module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1261(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1262(.a(gate11inter0), .b(s_102), .O(gate11inter1));
  and2  gate1263(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1264(.a(s_102), .O(gate11inter3));
  inv1  gate1265(.a(s_103), .O(gate11inter4));
  nand2 gate1266(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1267(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1268(.a(G5), .O(gate11inter7));
  inv1  gate1269(.a(G6), .O(gate11inter8));
  nand2 gate1270(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1271(.a(s_103), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1272(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1273(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1274(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1765(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1766(.a(gate16inter0), .b(s_174), .O(gate16inter1));
  and2  gate1767(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1768(.a(s_174), .O(gate16inter3));
  inv1  gate1769(.a(s_175), .O(gate16inter4));
  nand2 gate1770(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1771(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1772(.a(G15), .O(gate16inter7));
  inv1  gate1773(.a(G16), .O(gate16inter8));
  nand2 gate1774(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1775(.a(s_175), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1776(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1777(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1778(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1359(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1360(.a(gate17inter0), .b(s_116), .O(gate17inter1));
  and2  gate1361(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1362(.a(s_116), .O(gate17inter3));
  inv1  gate1363(.a(s_117), .O(gate17inter4));
  nand2 gate1364(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1365(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1366(.a(G17), .O(gate17inter7));
  inv1  gate1367(.a(G18), .O(gate17inter8));
  nand2 gate1368(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1369(.a(s_117), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1370(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1371(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1372(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1135(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1136(.a(gate27inter0), .b(s_84), .O(gate27inter1));
  and2  gate1137(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1138(.a(s_84), .O(gate27inter3));
  inv1  gate1139(.a(s_85), .O(gate27inter4));
  nand2 gate1140(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1141(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1142(.a(G2), .O(gate27inter7));
  inv1  gate1143(.a(G6), .O(gate27inter8));
  nand2 gate1144(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1145(.a(s_85), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1146(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1147(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1148(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1751(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1752(.a(gate29inter0), .b(s_172), .O(gate29inter1));
  and2  gate1753(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1754(.a(s_172), .O(gate29inter3));
  inv1  gate1755(.a(s_173), .O(gate29inter4));
  nand2 gate1756(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1757(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1758(.a(G3), .O(gate29inter7));
  inv1  gate1759(.a(G7), .O(gate29inter8));
  nand2 gate1760(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1761(.a(s_173), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1762(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1763(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1764(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate925(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate926(.a(gate31inter0), .b(s_54), .O(gate31inter1));
  and2  gate927(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate928(.a(s_54), .O(gate31inter3));
  inv1  gate929(.a(s_55), .O(gate31inter4));
  nand2 gate930(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate931(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate932(.a(G4), .O(gate31inter7));
  inv1  gate933(.a(G8), .O(gate31inter8));
  nand2 gate934(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate935(.a(s_55), .b(gate31inter3), .O(gate31inter10));
  nor2  gate936(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate937(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate938(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1667(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1668(.a(gate34inter0), .b(s_160), .O(gate34inter1));
  and2  gate1669(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1670(.a(s_160), .O(gate34inter3));
  inv1  gate1671(.a(s_161), .O(gate34inter4));
  nand2 gate1672(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1673(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1674(.a(G25), .O(gate34inter7));
  inv1  gate1675(.a(G29), .O(gate34inter8));
  nand2 gate1676(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1677(.a(s_161), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1678(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1679(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1680(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1457(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1458(.a(gate39inter0), .b(s_130), .O(gate39inter1));
  and2  gate1459(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1460(.a(s_130), .O(gate39inter3));
  inv1  gate1461(.a(s_131), .O(gate39inter4));
  nand2 gate1462(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1463(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1464(.a(G20), .O(gate39inter7));
  inv1  gate1465(.a(G24), .O(gate39inter8));
  nand2 gate1466(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1467(.a(s_131), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1468(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1469(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1470(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1499(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1500(.a(gate44inter0), .b(s_136), .O(gate44inter1));
  and2  gate1501(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1502(.a(s_136), .O(gate44inter3));
  inv1  gate1503(.a(s_137), .O(gate44inter4));
  nand2 gate1504(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1505(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1506(.a(G4), .O(gate44inter7));
  inv1  gate1507(.a(G269), .O(gate44inter8));
  nand2 gate1508(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1509(.a(s_137), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1510(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1511(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1512(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate869(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate870(.a(gate46inter0), .b(s_46), .O(gate46inter1));
  and2  gate871(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate872(.a(s_46), .O(gate46inter3));
  inv1  gate873(.a(s_47), .O(gate46inter4));
  nand2 gate874(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate875(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate876(.a(G6), .O(gate46inter7));
  inv1  gate877(.a(G272), .O(gate46inter8));
  nand2 gate878(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate879(.a(s_47), .b(gate46inter3), .O(gate46inter10));
  nor2  gate880(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate881(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate882(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1611(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1612(.a(gate52inter0), .b(s_152), .O(gate52inter1));
  and2  gate1613(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1614(.a(s_152), .O(gate52inter3));
  inv1  gate1615(.a(s_153), .O(gate52inter4));
  nand2 gate1616(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1617(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1618(.a(G12), .O(gate52inter7));
  inv1  gate1619(.a(G281), .O(gate52inter8));
  nand2 gate1620(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1621(.a(s_153), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1622(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1623(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1624(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate547(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate548(.a(gate59inter0), .b(s_0), .O(gate59inter1));
  and2  gate549(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate550(.a(s_0), .O(gate59inter3));
  inv1  gate551(.a(s_1), .O(gate59inter4));
  nand2 gate552(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate553(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate554(.a(G19), .O(gate59inter7));
  inv1  gate555(.a(G293), .O(gate59inter8));
  nand2 gate556(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate557(.a(s_1), .b(gate59inter3), .O(gate59inter10));
  nor2  gate558(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate559(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate560(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1289(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1290(.a(gate63inter0), .b(s_106), .O(gate63inter1));
  and2  gate1291(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1292(.a(s_106), .O(gate63inter3));
  inv1  gate1293(.a(s_107), .O(gate63inter4));
  nand2 gate1294(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1295(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1296(.a(G23), .O(gate63inter7));
  inv1  gate1297(.a(G299), .O(gate63inter8));
  nand2 gate1298(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1299(.a(s_107), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1300(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1301(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1302(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate743(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate744(.a(gate65inter0), .b(s_28), .O(gate65inter1));
  and2  gate745(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate746(.a(s_28), .O(gate65inter3));
  inv1  gate747(.a(s_29), .O(gate65inter4));
  nand2 gate748(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate749(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate750(.a(G25), .O(gate65inter7));
  inv1  gate751(.a(G302), .O(gate65inter8));
  nand2 gate752(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate753(.a(s_29), .b(gate65inter3), .O(gate65inter10));
  nor2  gate754(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate755(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate756(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate967(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate968(.a(gate70inter0), .b(s_60), .O(gate70inter1));
  and2  gate969(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate970(.a(s_60), .O(gate70inter3));
  inv1  gate971(.a(s_61), .O(gate70inter4));
  nand2 gate972(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate973(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate974(.a(G30), .O(gate70inter7));
  inv1  gate975(.a(G308), .O(gate70inter8));
  nand2 gate976(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate977(.a(s_61), .b(gate70inter3), .O(gate70inter10));
  nor2  gate978(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate979(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate980(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate785(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate786(.a(gate77inter0), .b(s_34), .O(gate77inter1));
  and2  gate787(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate788(.a(s_34), .O(gate77inter3));
  inv1  gate789(.a(s_35), .O(gate77inter4));
  nand2 gate790(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate791(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate792(.a(G2), .O(gate77inter7));
  inv1  gate793(.a(G320), .O(gate77inter8));
  nand2 gate794(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate795(.a(s_35), .b(gate77inter3), .O(gate77inter10));
  nor2  gate796(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate797(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate798(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1331(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1332(.a(gate83inter0), .b(s_112), .O(gate83inter1));
  and2  gate1333(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1334(.a(s_112), .O(gate83inter3));
  inv1  gate1335(.a(s_113), .O(gate83inter4));
  nand2 gate1336(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1337(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1338(.a(G11), .O(gate83inter7));
  inv1  gate1339(.a(G329), .O(gate83inter8));
  nand2 gate1340(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1341(.a(s_113), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1342(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1343(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1344(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate645(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate646(.a(gate88inter0), .b(s_14), .O(gate88inter1));
  and2  gate647(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate648(.a(s_14), .O(gate88inter3));
  inv1  gate649(.a(s_15), .O(gate88inter4));
  nand2 gate650(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate651(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate652(.a(G16), .O(gate88inter7));
  inv1  gate653(.a(G335), .O(gate88inter8));
  nand2 gate654(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate655(.a(s_15), .b(gate88inter3), .O(gate88inter10));
  nor2  gate656(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate657(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate658(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate673(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate674(.a(gate90inter0), .b(s_18), .O(gate90inter1));
  and2  gate675(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate676(.a(s_18), .O(gate90inter3));
  inv1  gate677(.a(s_19), .O(gate90inter4));
  nand2 gate678(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate679(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate680(.a(G21), .O(gate90inter7));
  inv1  gate681(.a(G338), .O(gate90inter8));
  nand2 gate682(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate683(.a(s_19), .b(gate90inter3), .O(gate90inter10));
  nor2  gate684(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate685(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate686(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate883(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate884(.a(gate91inter0), .b(s_48), .O(gate91inter1));
  and2  gate885(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate886(.a(s_48), .O(gate91inter3));
  inv1  gate887(.a(s_49), .O(gate91inter4));
  nand2 gate888(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate889(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate890(.a(G25), .O(gate91inter7));
  inv1  gate891(.a(G341), .O(gate91inter8));
  nand2 gate892(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate893(.a(s_49), .b(gate91inter3), .O(gate91inter10));
  nor2  gate894(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate895(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate896(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1471(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1472(.a(gate92inter0), .b(s_132), .O(gate92inter1));
  and2  gate1473(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1474(.a(s_132), .O(gate92inter3));
  inv1  gate1475(.a(s_133), .O(gate92inter4));
  nand2 gate1476(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1477(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1478(.a(G29), .O(gate92inter7));
  inv1  gate1479(.a(G341), .O(gate92inter8));
  nand2 gate1480(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1481(.a(s_133), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1482(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1483(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1484(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate995(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate996(.a(gate107inter0), .b(s_64), .O(gate107inter1));
  and2  gate997(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate998(.a(s_64), .O(gate107inter3));
  inv1  gate999(.a(s_65), .O(gate107inter4));
  nand2 gate1000(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1001(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1002(.a(G366), .O(gate107inter7));
  inv1  gate1003(.a(G367), .O(gate107inter8));
  nand2 gate1004(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1005(.a(s_65), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1006(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1007(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1008(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate981(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate982(.a(gate113inter0), .b(s_62), .O(gate113inter1));
  and2  gate983(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate984(.a(s_62), .O(gate113inter3));
  inv1  gate985(.a(s_63), .O(gate113inter4));
  nand2 gate986(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate987(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate988(.a(G378), .O(gate113inter7));
  inv1  gate989(.a(G379), .O(gate113inter8));
  nand2 gate990(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate991(.a(s_63), .b(gate113inter3), .O(gate113inter10));
  nor2  gate992(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate993(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate994(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate589(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate590(.a(gate119inter0), .b(s_6), .O(gate119inter1));
  and2  gate591(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate592(.a(s_6), .O(gate119inter3));
  inv1  gate593(.a(s_7), .O(gate119inter4));
  nand2 gate594(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate595(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate596(.a(G390), .O(gate119inter7));
  inv1  gate597(.a(G391), .O(gate119inter8));
  nand2 gate598(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate599(.a(s_7), .b(gate119inter3), .O(gate119inter10));
  nor2  gate600(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate601(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate602(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate799(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate800(.a(gate121inter0), .b(s_36), .O(gate121inter1));
  and2  gate801(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate802(.a(s_36), .O(gate121inter3));
  inv1  gate803(.a(s_37), .O(gate121inter4));
  nand2 gate804(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate805(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate806(.a(G394), .O(gate121inter7));
  inv1  gate807(.a(G395), .O(gate121inter8));
  nand2 gate808(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate809(.a(s_37), .b(gate121inter3), .O(gate121inter10));
  nor2  gate810(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate811(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate812(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1079(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1080(.a(gate123inter0), .b(s_76), .O(gate123inter1));
  and2  gate1081(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1082(.a(s_76), .O(gate123inter3));
  inv1  gate1083(.a(s_77), .O(gate123inter4));
  nand2 gate1084(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1085(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1086(.a(G398), .O(gate123inter7));
  inv1  gate1087(.a(G399), .O(gate123inter8));
  nand2 gate1088(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1089(.a(s_77), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1090(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1091(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1092(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate911(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate912(.a(gate128inter0), .b(s_52), .O(gate128inter1));
  and2  gate913(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate914(.a(s_52), .O(gate128inter3));
  inv1  gate915(.a(s_53), .O(gate128inter4));
  nand2 gate916(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate917(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate918(.a(G408), .O(gate128inter7));
  inv1  gate919(.a(G409), .O(gate128inter8));
  nand2 gate920(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate921(.a(s_53), .b(gate128inter3), .O(gate128inter10));
  nor2  gate922(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate923(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate924(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1583(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1584(.a(gate131inter0), .b(s_148), .O(gate131inter1));
  and2  gate1585(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1586(.a(s_148), .O(gate131inter3));
  inv1  gate1587(.a(s_149), .O(gate131inter4));
  nand2 gate1588(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1589(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1590(.a(G414), .O(gate131inter7));
  inv1  gate1591(.a(G415), .O(gate131inter8));
  nand2 gate1592(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1593(.a(s_149), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1594(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1595(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1596(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate897(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate898(.a(gate136inter0), .b(s_50), .O(gate136inter1));
  and2  gate899(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate900(.a(s_50), .O(gate136inter3));
  inv1  gate901(.a(s_51), .O(gate136inter4));
  nand2 gate902(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate903(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate904(.a(G424), .O(gate136inter7));
  inv1  gate905(.a(G425), .O(gate136inter8));
  nand2 gate906(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate907(.a(s_51), .b(gate136inter3), .O(gate136inter10));
  nor2  gate908(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate909(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate910(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1541(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1542(.a(gate139inter0), .b(s_142), .O(gate139inter1));
  and2  gate1543(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1544(.a(s_142), .O(gate139inter3));
  inv1  gate1545(.a(s_143), .O(gate139inter4));
  nand2 gate1546(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1547(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1548(.a(G438), .O(gate139inter7));
  inv1  gate1549(.a(G441), .O(gate139inter8));
  nand2 gate1550(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1551(.a(s_143), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1552(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1553(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1554(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1317(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1318(.a(gate142inter0), .b(s_110), .O(gate142inter1));
  and2  gate1319(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1320(.a(s_110), .O(gate142inter3));
  inv1  gate1321(.a(s_111), .O(gate142inter4));
  nand2 gate1322(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1323(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1324(.a(G456), .O(gate142inter7));
  inv1  gate1325(.a(G459), .O(gate142inter8));
  nand2 gate1326(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1327(.a(s_111), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1328(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1329(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1330(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1247(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1248(.a(gate144inter0), .b(s_100), .O(gate144inter1));
  and2  gate1249(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1250(.a(s_100), .O(gate144inter3));
  inv1  gate1251(.a(s_101), .O(gate144inter4));
  nand2 gate1252(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1253(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1254(.a(G468), .O(gate144inter7));
  inv1  gate1255(.a(G471), .O(gate144inter8));
  nand2 gate1256(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1257(.a(s_101), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1258(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1259(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1260(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1107(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1108(.a(gate149inter0), .b(s_80), .O(gate149inter1));
  and2  gate1109(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1110(.a(s_80), .O(gate149inter3));
  inv1  gate1111(.a(s_81), .O(gate149inter4));
  nand2 gate1112(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1113(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1114(.a(G498), .O(gate149inter7));
  inv1  gate1115(.a(G501), .O(gate149inter8));
  nand2 gate1116(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1117(.a(s_81), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1118(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1119(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1120(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1373(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1374(.a(gate154inter0), .b(s_118), .O(gate154inter1));
  and2  gate1375(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1376(.a(s_118), .O(gate154inter3));
  inv1  gate1377(.a(s_119), .O(gate154inter4));
  nand2 gate1378(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1379(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1380(.a(G429), .O(gate154inter7));
  inv1  gate1381(.a(G522), .O(gate154inter8));
  nand2 gate1382(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1383(.a(s_119), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1384(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1385(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1386(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate729(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate730(.a(gate157inter0), .b(s_26), .O(gate157inter1));
  and2  gate731(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate732(.a(s_26), .O(gate157inter3));
  inv1  gate733(.a(s_27), .O(gate157inter4));
  nand2 gate734(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate735(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate736(.a(G438), .O(gate157inter7));
  inv1  gate737(.a(G528), .O(gate157inter8));
  nand2 gate738(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate739(.a(s_27), .b(gate157inter3), .O(gate157inter10));
  nor2  gate740(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate741(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate742(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate813(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate814(.a(gate159inter0), .b(s_38), .O(gate159inter1));
  and2  gate815(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate816(.a(s_38), .O(gate159inter3));
  inv1  gate817(.a(s_39), .O(gate159inter4));
  nand2 gate818(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate819(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate820(.a(G444), .O(gate159inter7));
  inv1  gate821(.a(G531), .O(gate159inter8));
  nand2 gate822(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate823(.a(s_39), .b(gate159inter3), .O(gate159inter10));
  nor2  gate824(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate825(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate826(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1051(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1052(.a(gate160inter0), .b(s_72), .O(gate160inter1));
  and2  gate1053(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1054(.a(s_72), .O(gate160inter3));
  inv1  gate1055(.a(s_73), .O(gate160inter4));
  nand2 gate1056(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1057(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1058(.a(G447), .O(gate160inter7));
  inv1  gate1059(.a(G531), .O(gate160inter8));
  nand2 gate1060(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1061(.a(s_73), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1062(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1063(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1064(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1387(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1388(.a(gate162inter0), .b(s_120), .O(gate162inter1));
  and2  gate1389(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1390(.a(s_120), .O(gate162inter3));
  inv1  gate1391(.a(s_121), .O(gate162inter4));
  nand2 gate1392(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1393(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1394(.a(G453), .O(gate162inter7));
  inv1  gate1395(.a(G534), .O(gate162inter8));
  nand2 gate1396(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1397(.a(s_121), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1398(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1399(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1400(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1639(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1640(.a(gate165inter0), .b(s_156), .O(gate165inter1));
  and2  gate1641(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1642(.a(s_156), .O(gate165inter3));
  inv1  gate1643(.a(s_157), .O(gate165inter4));
  nand2 gate1644(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1645(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1646(.a(G462), .O(gate165inter7));
  inv1  gate1647(.a(G540), .O(gate165inter8));
  nand2 gate1648(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1649(.a(s_157), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1650(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1651(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1652(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1709(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1710(.a(gate171inter0), .b(s_166), .O(gate171inter1));
  and2  gate1711(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1712(.a(s_166), .O(gate171inter3));
  inv1  gate1713(.a(s_167), .O(gate171inter4));
  nand2 gate1714(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1715(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1716(.a(G480), .O(gate171inter7));
  inv1  gate1717(.a(G549), .O(gate171inter8));
  nand2 gate1718(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1719(.a(s_167), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1720(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1721(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1722(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1205(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1206(.a(gate172inter0), .b(s_94), .O(gate172inter1));
  and2  gate1207(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1208(.a(s_94), .O(gate172inter3));
  inv1  gate1209(.a(s_95), .O(gate172inter4));
  nand2 gate1210(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1211(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1212(.a(G483), .O(gate172inter7));
  inv1  gate1213(.a(G549), .O(gate172inter8));
  nand2 gate1214(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1215(.a(s_95), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1216(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1217(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1218(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1653(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1654(.a(gate175inter0), .b(s_158), .O(gate175inter1));
  and2  gate1655(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1656(.a(s_158), .O(gate175inter3));
  inv1  gate1657(.a(s_159), .O(gate175inter4));
  nand2 gate1658(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1659(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1660(.a(G492), .O(gate175inter7));
  inv1  gate1661(.a(G555), .O(gate175inter8));
  nand2 gate1662(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1663(.a(s_159), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1664(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1665(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1666(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1093(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1094(.a(gate176inter0), .b(s_78), .O(gate176inter1));
  and2  gate1095(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1096(.a(s_78), .O(gate176inter3));
  inv1  gate1097(.a(s_79), .O(gate176inter4));
  nand2 gate1098(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1099(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1100(.a(G495), .O(gate176inter7));
  inv1  gate1101(.a(G555), .O(gate176inter8));
  nand2 gate1102(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1103(.a(s_79), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1104(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1105(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1106(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate1037(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1038(.a(gate177inter0), .b(s_70), .O(gate177inter1));
  and2  gate1039(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1040(.a(s_70), .O(gate177inter3));
  inv1  gate1041(.a(s_71), .O(gate177inter4));
  nand2 gate1042(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1043(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1044(.a(G498), .O(gate177inter7));
  inv1  gate1045(.a(G558), .O(gate177inter8));
  nand2 gate1046(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1047(.a(s_71), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1048(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1049(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1050(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1821(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1822(.a(gate178inter0), .b(s_182), .O(gate178inter1));
  and2  gate1823(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1824(.a(s_182), .O(gate178inter3));
  inv1  gate1825(.a(s_183), .O(gate178inter4));
  nand2 gate1826(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1827(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1828(.a(G501), .O(gate178inter7));
  inv1  gate1829(.a(G558), .O(gate178inter8));
  nand2 gate1830(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1831(.a(s_183), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1832(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1833(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1834(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate953(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate954(.a(gate179inter0), .b(s_58), .O(gate179inter1));
  and2  gate955(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate956(.a(s_58), .O(gate179inter3));
  inv1  gate957(.a(s_59), .O(gate179inter4));
  nand2 gate958(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate959(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate960(.a(G504), .O(gate179inter7));
  inv1  gate961(.a(G561), .O(gate179inter8));
  nand2 gate962(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate963(.a(s_59), .b(gate179inter3), .O(gate179inter10));
  nor2  gate964(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate965(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate966(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate757(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate758(.a(gate187inter0), .b(s_30), .O(gate187inter1));
  and2  gate759(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate760(.a(s_30), .O(gate187inter3));
  inv1  gate761(.a(s_31), .O(gate187inter4));
  nand2 gate762(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate763(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate764(.a(G574), .O(gate187inter7));
  inv1  gate765(.a(G575), .O(gate187inter8));
  nand2 gate766(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate767(.a(s_31), .b(gate187inter3), .O(gate187inter10));
  nor2  gate768(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate769(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate770(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate575(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate576(.a(gate192inter0), .b(s_4), .O(gate192inter1));
  and2  gate577(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate578(.a(s_4), .O(gate192inter3));
  inv1  gate579(.a(s_5), .O(gate192inter4));
  nand2 gate580(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate581(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate582(.a(G584), .O(gate192inter7));
  inv1  gate583(.a(G585), .O(gate192inter8));
  nand2 gate584(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate585(.a(s_5), .b(gate192inter3), .O(gate192inter10));
  nor2  gate586(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate587(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate588(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1849(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1850(.a(gate196inter0), .b(s_186), .O(gate196inter1));
  and2  gate1851(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1852(.a(s_186), .O(gate196inter3));
  inv1  gate1853(.a(s_187), .O(gate196inter4));
  nand2 gate1854(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1855(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1856(.a(G592), .O(gate196inter7));
  inv1  gate1857(.a(G593), .O(gate196inter8));
  nand2 gate1858(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1859(.a(s_187), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1860(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1861(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1862(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1527(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1528(.a(gate198inter0), .b(s_140), .O(gate198inter1));
  and2  gate1529(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1530(.a(s_140), .O(gate198inter3));
  inv1  gate1531(.a(s_141), .O(gate198inter4));
  nand2 gate1532(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1533(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1534(.a(G596), .O(gate198inter7));
  inv1  gate1535(.a(G597), .O(gate198inter8));
  nand2 gate1536(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1537(.a(s_141), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1538(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1539(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1540(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1793(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1794(.a(gate202inter0), .b(s_178), .O(gate202inter1));
  and2  gate1795(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1796(.a(s_178), .O(gate202inter3));
  inv1  gate1797(.a(s_179), .O(gate202inter4));
  nand2 gate1798(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1799(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1800(.a(G612), .O(gate202inter7));
  inv1  gate1801(.a(G617), .O(gate202inter8));
  nand2 gate1802(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1803(.a(s_179), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1804(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1805(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1806(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1807(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1808(.a(gate215inter0), .b(s_180), .O(gate215inter1));
  and2  gate1809(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1810(.a(s_180), .O(gate215inter3));
  inv1  gate1811(.a(s_181), .O(gate215inter4));
  nand2 gate1812(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1813(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1814(.a(G607), .O(gate215inter7));
  inv1  gate1815(.a(G675), .O(gate215inter8));
  nand2 gate1816(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1817(.a(s_181), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1818(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1819(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1820(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1681(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1682(.a(gate217inter0), .b(s_162), .O(gate217inter1));
  and2  gate1683(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1684(.a(s_162), .O(gate217inter3));
  inv1  gate1685(.a(s_163), .O(gate217inter4));
  nand2 gate1686(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1687(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1688(.a(G622), .O(gate217inter7));
  inv1  gate1689(.a(G678), .O(gate217inter8));
  nand2 gate1690(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1691(.a(s_163), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1692(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1693(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1694(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1345(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1346(.a(gate218inter0), .b(s_114), .O(gate218inter1));
  and2  gate1347(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1348(.a(s_114), .O(gate218inter3));
  inv1  gate1349(.a(s_115), .O(gate218inter4));
  nand2 gate1350(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1351(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1352(.a(G627), .O(gate218inter7));
  inv1  gate1353(.a(G678), .O(gate218inter8));
  nand2 gate1354(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1355(.a(s_115), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1356(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1357(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1358(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1597(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1598(.a(gate223inter0), .b(s_150), .O(gate223inter1));
  and2  gate1599(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1600(.a(s_150), .O(gate223inter3));
  inv1  gate1601(.a(s_151), .O(gate223inter4));
  nand2 gate1602(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1603(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1604(.a(G627), .O(gate223inter7));
  inv1  gate1605(.a(G687), .O(gate223inter8));
  nand2 gate1606(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1607(.a(s_151), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1608(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1609(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1610(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1625(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1626(.a(gate227inter0), .b(s_154), .O(gate227inter1));
  and2  gate1627(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1628(.a(s_154), .O(gate227inter3));
  inv1  gate1629(.a(s_155), .O(gate227inter4));
  nand2 gate1630(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1631(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1632(.a(G694), .O(gate227inter7));
  inv1  gate1633(.a(G695), .O(gate227inter8));
  nand2 gate1634(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1635(.a(s_155), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1636(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1637(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1638(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1779(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1780(.a(gate228inter0), .b(s_176), .O(gate228inter1));
  and2  gate1781(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1782(.a(s_176), .O(gate228inter3));
  inv1  gate1783(.a(s_177), .O(gate228inter4));
  nand2 gate1784(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1785(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1786(.a(G696), .O(gate228inter7));
  inv1  gate1787(.a(G697), .O(gate228inter8));
  nand2 gate1788(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1789(.a(s_177), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1790(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1791(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1792(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate603(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate604(.a(gate237inter0), .b(s_8), .O(gate237inter1));
  and2  gate605(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate606(.a(s_8), .O(gate237inter3));
  inv1  gate607(.a(s_9), .O(gate237inter4));
  nand2 gate608(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate609(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate610(.a(G254), .O(gate237inter7));
  inv1  gate611(.a(G706), .O(gate237inter8));
  nand2 gate612(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate613(.a(s_9), .b(gate237inter3), .O(gate237inter10));
  nor2  gate614(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate615(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate616(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate841(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate842(.a(gate243inter0), .b(s_42), .O(gate243inter1));
  and2  gate843(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate844(.a(s_42), .O(gate243inter3));
  inv1  gate845(.a(s_43), .O(gate243inter4));
  nand2 gate846(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate847(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate848(.a(G245), .O(gate243inter7));
  inv1  gate849(.a(G733), .O(gate243inter8));
  nand2 gate850(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate851(.a(s_43), .b(gate243inter3), .O(gate243inter10));
  nor2  gate852(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate853(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate854(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1695(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1696(.a(gate247inter0), .b(s_164), .O(gate247inter1));
  and2  gate1697(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1698(.a(s_164), .O(gate247inter3));
  inv1  gate1699(.a(s_165), .O(gate247inter4));
  nand2 gate1700(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1701(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1702(.a(G251), .O(gate247inter7));
  inv1  gate1703(.a(G739), .O(gate247inter8));
  nand2 gate1704(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1705(.a(s_165), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1706(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1707(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1708(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1191(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1192(.a(gate248inter0), .b(s_92), .O(gate248inter1));
  and2  gate1193(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1194(.a(s_92), .O(gate248inter3));
  inv1  gate1195(.a(s_93), .O(gate248inter4));
  nand2 gate1196(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1197(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1198(.a(G727), .O(gate248inter7));
  inv1  gate1199(.a(G739), .O(gate248inter8));
  nand2 gate1200(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1201(.a(s_93), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1202(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1203(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1204(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1555(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1556(.a(gate249inter0), .b(s_144), .O(gate249inter1));
  and2  gate1557(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1558(.a(s_144), .O(gate249inter3));
  inv1  gate1559(.a(s_145), .O(gate249inter4));
  nand2 gate1560(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1561(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1562(.a(G254), .O(gate249inter7));
  inv1  gate1563(.a(G742), .O(gate249inter8));
  nand2 gate1564(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1565(.a(s_145), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1566(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1567(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1568(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1877(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1878(.a(gate251inter0), .b(s_190), .O(gate251inter1));
  and2  gate1879(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1880(.a(s_190), .O(gate251inter3));
  inv1  gate1881(.a(s_191), .O(gate251inter4));
  nand2 gate1882(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1883(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1884(.a(G257), .O(gate251inter7));
  inv1  gate1885(.a(G745), .O(gate251inter8));
  nand2 gate1886(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1887(.a(s_191), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1888(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1889(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1890(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1009(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1010(.a(gate253inter0), .b(s_66), .O(gate253inter1));
  and2  gate1011(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1012(.a(s_66), .O(gate253inter3));
  inv1  gate1013(.a(s_67), .O(gate253inter4));
  nand2 gate1014(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1015(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1016(.a(G260), .O(gate253inter7));
  inv1  gate1017(.a(G748), .O(gate253inter8));
  nand2 gate1018(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1019(.a(s_67), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1020(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1021(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1022(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1723(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1724(.a(gate258inter0), .b(s_168), .O(gate258inter1));
  and2  gate1725(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1726(.a(s_168), .O(gate258inter3));
  inv1  gate1727(.a(s_169), .O(gate258inter4));
  nand2 gate1728(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1729(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1730(.a(G756), .O(gate258inter7));
  inv1  gate1731(.a(G757), .O(gate258inter8));
  nand2 gate1732(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1733(.a(s_169), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1734(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1735(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1736(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1275(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1276(.a(gate260inter0), .b(s_104), .O(gate260inter1));
  and2  gate1277(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1278(.a(s_104), .O(gate260inter3));
  inv1  gate1279(.a(s_105), .O(gate260inter4));
  nand2 gate1280(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1281(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1282(.a(G760), .O(gate260inter7));
  inv1  gate1283(.a(G761), .O(gate260inter8));
  nand2 gate1284(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1285(.a(s_105), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1286(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1287(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1288(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1233(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1234(.a(gate264inter0), .b(s_98), .O(gate264inter1));
  and2  gate1235(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1236(.a(s_98), .O(gate264inter3));
  inv1  gate1237(.a(s_99), .O(gate264inter4));
  nand2 gate1238(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1239(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1240(.a(G768), .O(gate264inter7));
  inv1  gate1241(.a(G769), .O(gate264inter8));
  nand2 gate1242(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1243(.a(s_99), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1244(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1245(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1246(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1121(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1122(.a(gate267inter0), .b(s_82), .O(gate267inter1));
  and2  gate1123(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1124(.a(s_82), .O(gate267inter3));
  inv1  gate1125(.a(s_83), .O(gate267inter4));
  nand2 gate1126(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1127(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1128(.a(G648), .O(gate267inter7));
  inv1  gate1129(.a(G776), .O(gate267inter8));
  nand2 gate1130(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1131(.a(s_83), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1132(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1133(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1134(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate617(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate618(.a(gate268inter0), .b(s_10), .O(gate268inter1));
  and2  gate619(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate620(.a(s_10), .O(gate268inter3));
  inv1  gate621(.a(s_11), .O(gate268inter4));
  nand2 gate622(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate623(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate624(.a(G651), .O(gate268inter7));
  inv1  gate625(.a(G779), .O(gate268inter8));
  nand2 gate626(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate627(.a(s_11), .b(gate268inter3), .O(gate268inter10));
  nor2  gate628(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate629(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate630(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate659(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate660(.a(gate393inter0), .b(s_16), .O(gate393inter1));
  and2  gate661(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate662(.a(s_16), .O(gate393inter3));
  inv1  gate663(.a(s_17), .O(gate393inter4));
  nand2 gate664(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate665(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate666(.a(G7), .O(gate393inter7));
  inv1  gate667(.a(G1054), .O(gate393inter8));
  nand2 gate668(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate669(.a(s_17), .b(gate393inter3), .O(gate393inter10));
  nor2  gate670(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate671(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate672(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1863(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1864(.a(gate394inter0), .b(s_188), .O(gate394inter1));
  and2  gate1865(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1866(.a(s_188), .O(gate394inter3));
  inv1  gate1867(.a(s_189), .O(gate394inter4));
  nand2 gate1868(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1869(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1870(.a(G8), .O(gate394inter7));
  inv1  gate1871(.a(G1057), .O(gate394inter8));
  nand2 gate1872(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1873(.a(s_189), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1874(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1875(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1876(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1429(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1430(.a(gate397inter0), .b(s_126), .O(gate397inter1));
  and2  gate1431(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1432(.a(s_126), .O(gate397inter3));
  inv1  gate1433(.a(s_127), .O(gate397inter4));
  nand2 gate1434(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1435(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1436(.a(G11), .O(gate397inter7));
  inv1  gate1437(.a(G1066), .O(gate397inter8));
  nand2 gate1438(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1439(.a(s_127), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1440(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1441(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1442(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1149(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1150(.a(gate403inter0), .b(s_86), .O(gate403inter1));
  and2  gate1151(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1152(.a(s_86), .O(gate403inter3));
  inv1  gate1153(.a(s_87), .O(gate403inter4));
  nand2 gate1154(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1155(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1156(.a(G17), .O(gate403inter7));
  inv1  gate1157(.a(G1084), .O(gate403inter8));
  nand2 gate1158(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1159(.a(s_87), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1160(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1161(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1162(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1065(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1066(.a(gate414inter0), .b(s_74), .O(gate414inter1));
  and2  gate1067(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1068(.a(s_74), .O(gate414inter3));
  inv1  gate1069(.a(s_75), .O(gate414inter4));
  nand2 gate1070(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1071(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1072(.a(G28), .O(gate414inter7));
  inv1  gate1073(.a(G1117), .O(gate414inter8));
  nand2 gate1074(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1075(.a(s_75), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1076(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1077(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1078(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1401(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1402(.a(gate422inter0), .b(s_122), .O(gate422inter1));
  and2  gate1403(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1404(.a(s_122), .O(gate422inter3));
  inv1  gate1405(.a(s_123), .O(gate422inter4));
  nand2 gate1406(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1407(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1408(.a(G1039), .O(gate422inter7));
  inv1  gate1409(.a(G1135), .O(gate422inter8));
  nand2 gate1410(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1411(.a(s_123), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1412(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1413(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1414(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1219(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1220(.a(gate424inter0), .b(s_96), .O(gate424inter1));
  and2  gate1221(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1222(.a(s_96), .O(gate424inter3));
  inv1  gate1223(.a(s_97), .O(gate424inter4));
  nand2 gate1224(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1225(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1226(.a(G1042), .O(gate424inter7));
  inv1  gate1227(.a(G1138), .O(gate424inter8));
  nand2 gate1228(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1229(.a(s_97), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1230(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1231(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1232(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate855(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate856(.a(gate430inter0), .b(s_44), .O(gate430inter1));
  and2  gate857(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate858(.a(s_44), .O(gate430inter3));
  inv1  gate859(.a(s_45), .O(gate430inter4));
  nand2 gate860(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate861(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate862(.a(G1051), .O(gate430inter7));
  inv1  gate863(.a(G1147), .O(gate430inter8));
  nand2 gate864(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate865(.a(s_45), .b(gate430inter3), .O(gate430inter10));
  nor2  gate866(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate867(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate868(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1569(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1570(.a(gate432inter0), .b(s_146), .O(gate432inter1));
  and2  gate1571(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1572(.a(s_146), .O(gate432inter3));
  inv1  gate1573(.a(s_147), .O(gate432inter4));
  nand2 gate1574(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1575(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1576(.a(G1054), .O(gate432inter7));
  inv1  gate1577(.a(G1150), .O(gate432inter8));
  nand2 gate1578(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1579(.a(s_147), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1580(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1581(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1582(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1835(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1836(.a(gate437inter0), .b(s_184), .O(gate437inter1));
  and2  gate1837(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1838(.a(s_184), .O(gate437inter3));
  inv1  gate1839(.a(s_185), .O(gate437inter4));
  nand2 gate1840(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1841(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1842(.a(G10), .O(gate437inter7));
  inv1  gate1843(.a(G1159), .O(gate437inter8));
  nand2 gate1844(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1845(.a(s_185), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1846(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1847(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1848(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate561(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate562(.a(gate438inter0), .b(s_2), .O(gate438inter1));
  and2  gate563(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate564(.a(s_2), .O(gate438inter3));
  inv1  gate565(.a(s_3), .O(gate438inter4));
  nand2 gate566(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate567(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate568(.a(G1063), .O(gate438inter7));
  inv1  gate569(.a(G1159), .O(gate438inter8));
  nand2 gate570(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate571(.a(s_3), .b(gate438inter3), .O(gate438inter10));
  nor2  gate572(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate573(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate574(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate701(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate702(.a(gate447inter0), .b(s_22), .O(gate447inter1));
  and2  gate703(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate704(.a(s_22), .O(gate447inter3));
  inv1  gate705(.a(s_23), .O(gate447inter4));
  nand2 gate706(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate707(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate708(.a(G15), .O(gate447inter7));
  inv1  gate709(.a(G1174), .O(gate447inter8));
  nand2 gate710(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate711(.a(s_23), .b(gate447inter3), .O(gate447inter10));
  nor2  gate712(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate713(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate714(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate687(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate688(.a(gate452inter0), .b(s_20), .O(gate452inter1));
  and2  gate689(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate690(.a(s_20), .O(gate452inter3));
  inv1  gate691(.a(s_21), .O(gate452inter4));
  nand2 gate692(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate693(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate694(.a(G1084), .O(gate452inter7));
  inv1  gate695(.a(G1180), .O(gate452inter8));
  nand2 gate696(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate697(.a(s_21), .b(gate452inter3), .O(gate452inter10));
  nor2  gate698(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate699(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate700(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate771(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate772(.a(gate453inter0), .b(s_32), .O(gate453inter1));
  and2  gate773(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate774(.a(s_32), .O(gate453inter3));
  inv1  gate775(.a(s_33), .O(gate453inter4));
  nand2 gate776(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate777(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate778(.a(G18), .O(gate453inter7));
  inv1  gate779(.a(G1183), .O(gate453inter8));
  nand2 gate780(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate781(.a(s_33), .b(gate453inter3), .O(gate453inter10));
  nor2  gate782(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate783(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate784(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1485(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1486(.a(gate462inter0), .b(s_134), .O(gate462inter1));
  and2  gate1487(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1488(.a(s_134), .O(gate462inter3));
  inv1  gate1489(.a(s_135), .O(gate462inter4));
  nand2 gate1490(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1491(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1492(.a(G1099), .O(gate462inter7));
  inv1  gate1493(.a(G1195), .O(gate462inter8));
  nand2 gate1494(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1495(.a(s_135), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1496(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1497(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1498(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1513(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1514(.a(gate464inter0), .b(s_138), .O(gate464inter1));
  and2  gate1515(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1516(.a(s_138), .O(gate464inter3));
  inv1  gate1517(.a(s_139), .O(gate464inter4));
  nand2 gate1518(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1519(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1520(.a(G1102), .O(gate464inter7));
  inv1  gate1521(.a(G1198), .O(gate464inter8));
  nand2 gate1522(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1523(.a(s_139), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1524(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1525(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1526(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate715(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate716(.a(gate472inter0), .b(s_24), .O(gate472inter1));
  and2  gate717(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate718(.a(s_24), .O(gate472inter3));
  inv1  gate719(.a(s_25), .O(gate472inter4));
  nand2 gate720(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate721(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate722(.a(G1114), .O(gate472inter7));
  inv1  gate723(.a(G1210), .O(gate472inter8));
  nand2 gate724(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate725(.a(s_25), .b(gate472inter3), .O(gate472inter10));
  nor2  gate726(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate727(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate728(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1023(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1024(.a(gate477inter0), .b(s_68), .O(gate477inter1));
  and2  gate1025(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1026(.a(s_68), .O(gate477inter3));
  inv1  gate1027(.a(s_69), .O(gate477inter4));
  nand2 gate1028(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1029(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1030(.a(G30), .O(gate477inter7));
  inv1  gate1031(.a(G1219), .O(gate477inter8));
  nand2 gate1032(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1033(.a(s_69), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1034(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1035(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1036(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate939(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate940(.a(gate481inter0), .b(s_56), .O(gate481inter1));
  and2  gate941(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate942(.a(s_56), .O(gate481inter3));
  inv1  gate943(.a(s_57), .O(gate481inter4));
  nand2 gate944(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate945(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate946(.a(G32), .O(gate481inter7));
  inv1  gate947(.a(G1225), .O(gate481inter8));
  nand2 gate948(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate949(.a(s_57), .b(gate481inter3), .O(gate481inter10));
  nor2  gate950(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate951(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate952(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate827(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate828(.a(gate482inter0), .b(s_40), .O(gate482inter1));
  and2  gate829(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate830(.a(s_40), .O(gate482inter3));
  inv1  gate831(.a(s_41), .O(gate482inter4));
  nand2 gate832(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate833(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate834(.a(G1129), .O(gate482inter7));
  inv1  gate835(.a(G1225), .O(gate482inter8));
  nand2 gate836(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate837(.a(s_41), .b(gate482inter3), .O(gate482inter10));
  nor2  gate838(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate839(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate840(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1415(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1416(.a(gate488inter0), .b(s_124), .O(gate488inter1));
  and2  gate1417(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1418(.a(s_124), .O(gate488inter3));
  inv1  gate1419(.a(s_125), .O(gate488inter4));
  nand2 gate1420(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1421(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1422(.a(G1238), .O(gate488inter7));
  inv1  gate1423(.a(G1239), .O(gate488inter8));
  nand2 gate1424(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1425(.a(s_125), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1426(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1427(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1428(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1303(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1304(.a(gate490inter0), .b(s_108), .O(gate490inter1));
  and2  gate1305(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1306(.a(s_108), .O(gate490inter3));
  inv1  gate1307(.a(s_109), .O(gate490inter4));
  nand2 gate1308(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1309(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1310(.a(G1242), .O(gate490inter7));
  inv1  gate1311(.a(G1243), .O(gate490inter8));
  nand2 gate1312(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1313(.a(s_109), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1314(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1315(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1316(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate631(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate632(.a(gate491inter0), .b(s_12), .O(gate491inter1));
  and2  gate633(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate634(.a(s_12), .O(gate491inter3));
  inv1  gate635(.a(s_13), .O(gate491inter4));
  nand2 gate636(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate637(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate638(.a(G1244), .O(gate491inter7));
  inv1  gate639(.a(G1245), .O(gate491inter8));
  nand2 gate640(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate641(.a(s_13), .b(gate491inter3), .O(gate491inter10));
  nor2  gate642(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate643(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate644(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1443(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1444(.a(gate499inter0), .b(s_128), .O(gate499inter1));
  and2  gate1445(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1446(.a(s_128), .O(gate499inter3));
  inv1  gate1447(.a(s_129), .O(gate499inter4));
  nand2 gate1448(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1449(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1450(.a(G1260), .O(gate499inter7));
  inv1  gate1451(.a(G1261), .O(gate499inter8));
  nand2 gate1452(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1453(.a(s_129), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1454(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1455(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1456(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1163(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1164(.a(gate504inter0), .b(s_88), .O(gate504inter1));
  and2  gate1165(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1166(.a(s_88), .O(gate504inter3));
  inv1  gate1167(.a(s_89), .O(gate504inter4));
  nand2 gate1168(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1169(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1170(.a(G1270), .O(gate504inter7));
  inv1  gate1171(.a(G1271), .O(gate504inter8));
  nand2 gate1172(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1173(.a(s_89), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1174(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1175(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1176(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1177(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1178(.a(gate510inter0), .b(s_90), .O(gate510inter1));
  and2  gate1179(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1180(.a(s_90), .O(gate510inter3));
  inv1  gate1181(.a(s_91), .O(gate510inter4));
  nand2 gate1182(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1183(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1184(.a(G1282), .O(gate510inter7));
  inv1  gate1185(.a(G1283), .O(gate510inter8));
  nand2 gate1186(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1187(.a(s_91), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1188(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1189(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1190(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1737(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1738(.a(gate511inter0), .b(s_170), .O(gate511inter1));
  and2  gate1739(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1740(.a(s_170), .O(gate511inter3));
  inv1  gate1741(.a(s_171), .O(gate511inter4));
  nand2 gate1742(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1743(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1744(.a(G1284), .O(gate511inter7));
  inv1  gate1745(.a(G1285), .O(gate511inter8));
  nand2 gate1746(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1747(.a(s_171), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1748(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1749(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1750(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule