module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381, s_382, s_383, s_384, s_385, s_386, s_387, s_388, s_389, s_390, s_391, s_392, s_393, s_394, s_395, s_396, s_397, s_398, s_399, s_400, s_401;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2619(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2620(.a(gate10inter0), .b(s_296), .O(gate10inter1));
  and2  gate2621(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2622(.a(s_296), .O(gate10inter3));
  inv1  gate2623(.a(s_297), .O(gate10inter4));
  nand2 gate2624(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2625(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2626(.a(G3), .O(gate10inter7));
  inv1  gate2627(.a(G4), .O(gate10inter8));
  nand2 gate2628(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2629(.a(s_297), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2630(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2631(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2632(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate967(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate968(.a(gate13inter0), .b(s_60), .O(gate13inter1));
  and2  gate969(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate970(.a(s_60), .O(gate13inter3));
  inv1  gate971(.a(s_61), .O(gate13inter4));
  nand2 gate972(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate973(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate974(.a(G9), .O(gate13inter7));
  inv1  gate975(.a(G10), .O(gate13inter8));
  nand2 gate976(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate977(.a(s_61), .b(gate13inter3), .O(gate13inter10));
  nor2  gate978(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate979(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate980(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1233(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1234(.a(gate18inter0), .b(s_98), .O(gate18inter1));
  and2  gate1235(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1236(.a(s_98), .O(gate18inter3));
  inv1  gate1237(.a(s_99), .O(gate18inter4));
  nand2 gate1238(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1239(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1240(.a(G19), .O(gate18inter7));
  inv1  gate1241(.a(G20), .O(gate18inter8));
  nand2 gate1242(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1243(.a(s_99), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1244(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1245(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1246(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2871(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2872(.a(gate19inter0), .b(s_332), .O(gate19inter1));
  and2  gate2873(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2874(.a(s_332), .O(gate19inter3));
  inv1  gate2875(.a(s_333), .O(gate19inter4));
  nand2 gate2876(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2877(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2878(.a(G21), .O(gate19inter7));
  inv1  gate2879(.a(G22), .O(gate19inter8));
  nand2 gate2880(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2881(.a(s_333), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2882(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2883(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2884(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2969(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2970(.a(gate20inter0), .b(s_346), .O(gate20inter1));
  and2  gate2971(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2972(.a(s_346), .O(gate20inter3));
  inv1  gate2973(.a(s_347), .O(gate20inter4));
  nand2 gate2974(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2975(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2976(.a(G23), .O(gate20inter7));
  inv1  gate2977(.a(G24), .O(gate20inter8));
  nand2 gate2978(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2979(.a(s_347), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2980(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2981(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2982(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1275(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1276(.a(gate22inter0), .b(s_104), .O(gate22inter1));
  and2  gate1277(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1278(.a(s_104), .O(gate22inter3));
  inv1  gate1279(.a(s_105), .O(gate22inter4));
  nand2 gate1280(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1281(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1282(.a(G27), .O(gate22inter7));
  inv1  gate1283(.a(G28), .O(gate22inter8));
  nand2 gate1284(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1285(.a(s_105), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1286(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1287(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1288(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate799(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate800(.a(gate23inter0), .b(s_36), .O(gate23inter1));
  and2  gate801(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate802(.a(s_36), .O(gate23inter3));
  inv1  gate803(.a(s_37), .O(gate23inter4));
  nand2 gate804(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate805(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate806(.a(G29), .O(gate23inter7));
  inv1  gate807(.a(G30), .O(gate23inter8));
  nand2 gate808(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate809(.a(s_37), .b(gate23inter3), .O(gate23inter10));
  nor2  gate810(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate811(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate812(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1303(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1304(.a(gate25inter0), .b(s_108), .O(gate25inter1));
  and2  gate1305(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1306(.a(s_108), .O(gate25inter3));
  inv1  gate1307(.a(s_109), .O(gate25inter4));
  nand2 gate1308(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1309(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1310(.a(G1), .O(gate25inter7));
  inv1  gate1311(.a(G5), .O(gate25inter8));
  nand2 gate1312(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1313(.a(s_109), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1314(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1315(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1316(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate869(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate870(.a(gate26inter0), .b(s_46), .O(gate26inter1));
  and2  gate871(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate872(.a(s_46), .O(gate26inter3));
  inv1  gate873(.a(s_47), .O(gate26inter4));
  nand2 gate874(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate875(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate876(.a(G9), .O(gate26inter7));
  inv1  gate877(.a(G13), .O(gate26inter8));
  nand2 gate878(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate879(.a(s_47), .b(gate26inter3), .O(gate26inter10));
  nor2  gate880(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate881(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate882(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2381(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2382(.a(gate28inter0), .b(s_262), .O(gate28inter1));
  and2  gate2383(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2384(.a(s_262), .O(gate28inter3));
  inv1  gate2385(.a(s_263), .O(gate28inter4));
  nand2 gate2386(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2387(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2388(.a(G10), .O(gate28inter7));
  inv1  gate2389(.a(G14), .O(gate28inter8));
  nand2 gate2390(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2391(.a(s_263), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2392(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2393(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2394(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate3025(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate3026(.a(gate43inter0), .b(s_354), .O(gate43inter1));
  and2  gate3027(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate3028(.a(s_354), .O(gate43inter3));
  inv1  gate3029(.a(s_355), .O(gate43inter4));
  nand2 gate3030(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate3031(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate3032(.a(G3), .O(gate43inter7));
  inv1  gate3033(.a(G269), .O(gate43inter8));
  nand2 gate3034(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate3035(.a(s_355), .b(gate43inter3), .O(gate43inter10));
  nor2  gate3036(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate3037(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate3038(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2157(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2158(.a(gate44inter0), .b(s_230), .O(gate44inter1));
  and2  gate2159(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2160(.a(s_230), .O(gate44inter3));
  inv1  gate2161(.a(s_231), .O(gate44inter4));
  nand2 gate2162(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2163(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2164(.a(G4), .O(gate44inter7));
  inv1  gate2165(.a(G269), .O(gate44inter8));
  nand2 gate2166(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2167(.a(s_231), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2168(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2169(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2170(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate3249(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate3250(.a(gate46inter0), .b(s_386), .O(gate46inter1));
  and2  gate3251(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate3252(.a(s_386), .O(gate46inter3));
  inv1  gate3253(.a(s_387), .O(gate46inter4));
  nand2 gate3254(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate3255(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate3256(.a(G6), .O(gate46inter7));
  inv1  gate3257(.a(G272), .O(gate46inter8));
  nand2 gate3258(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate3259(.a(s_387), .b(gate46inter3), .O(gate46inter10));
  nor2  gate3260(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate3261(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate3262(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2437(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2438(.a(gate47inter0), .b(s_270), .O(gate47inter1));
  and2  gate2439(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2440(.a(s_270), .O(gate47inter3));
  inv1  gate2441(.a(s_271), .O(gate47inter4));
  nand2 gate2442(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2443(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2444(.a(G7), .O(gate47inter7));
  inv1  gate2445(.a(G275), .O(gate47inter8));
  nand2 gate2446(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2447(.a(s_271), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2448(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2449(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2450(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate3333(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate3334(.a(gate49inter0), .b(s_398), .O(gate49inter1));
  and2  gate3335(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate3336(.a(s_398), .O(gate49inter3));
  inv1  gate3337(.a(s_399), .O(gate49inter4));
  nand2 gate3338(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate3339(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate3340(.a(G9), .O(gate49inter7));
  inv1  gate3341(.a(G278), .O(gate49inter8));
  nand2 gate3342(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate3343(.a(s_399), .b(gate49inter3), .O(gate49inter10));
  nor2  gate3344(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate3345(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate3346(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate3263(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate3264(.a(gate54inter0), .b(s_388), .O(gate54inter1));
  and2  gate3265(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate3266(.a(s_388), .O(gate54inter3));
  inv1  gate3267(.a(s_389), .O(gate54inter4));
  nand2 gate3268(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate3269(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate3270(.a(G14), .O(gate54inter7));
  inv1  gate3271(.a(G284), .O(gate54inter8));
  nand2 gate3272(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate3273(.a(s_389), .b(gate54inter3), .O(gate54inter10));
  nor2  gate3274(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate3275(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate3276(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1093(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1094(.a(gate56inter0), .b(s_78), .O(gate56inter1));
  and2  gate1095(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1096(.a(s_78), .O(gate56inter3));
  inv1  gate1097(.a(s_79), .O(gate56inter4));
  nand2 gate1098(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1099(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1100(.a(G16), .O(gate56inter7));
  inv1  gate1101(.a(G287), .O(gate56inter8));
  nand2 gate1102(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1103(.a(s_79), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1104(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1105(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1106(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1065(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1066(.a(gate57inter0), .b(s_74), .O(gate57inter1));
  and2  gate1067(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1068(.a(s_74), .O(gate57inter3));
  inv1  gate1069(.a(s_75), .O(gate57inter4));
  nand2 gate1070(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1071(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1072(.a(G17), .O(gate57inter7));
  inv1  gate1073(.a(G290), .O(gate57inter8));
  nand2 gate1074(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1075(.a(s_75), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1076(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1077(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1078(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1261(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1262(.a(gate59inter0), .b(s_102), .O(gate59inter1));
  and2  gate1263(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1264(.a(s_102), .O(gate59inter3));
  inv1  gate1265(.a(s_103), .O(gate59inter4));
  nand2 gate1266(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1267(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1268(.a(G19), .O(gate59inter7));
  inv1  gate1269(.a(G293), .O(gate59inter8));
  nand2 gate1270(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1271(.a(s_103), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1272(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1273(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1274(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1947(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1948(.a(gate61inter0), .b(s_200), .O(gate61inter1));
  and2  gate1949(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1950(.a(s_200), .O(gate61inter3));
  inv1  gate1951(.a(s_201), .O(gate61inter4));
  nand2 gate1952(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1953(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1954(.a(G21), .O(gate61inter7));
  inv1  gate1955(.a(G296), .O(gate61inter8));
  nand2 gate1956(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1957(.a(s_201), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1958(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1959(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1960(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1653(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1654(.a(gate63inter0), .b(s_158), .O(gate63inter1));
  and2  gate1655(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1656(.a(s_158), .O(gate63inter3));
  inv1  gate1657(.a(s_159), .O(gate63inter4));
  nand2 gate1658(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1659(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1660(.a(G23), .O(gate63inter7));
  inv1  gate1661(.a(G299), .O(gate63inter8));
  nand2 gate1662(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1663(.a(s_159), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1664(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1665(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1666(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1569(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1570(.a(gate65inter0), .b(s_146), .O(gate65inter1));
  and2  gate1571(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1572(.a(s_146), .O(gate65inter3));
  inv1  gate1573(.a(s_147), .O(gate65inter4));
  nand2 gate1574(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1575(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1576(.a(G25), .O(gate65inter7));
  inv1  gate1577(.a(G302), .O(gate65inter8));
  nand2 gate1578(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1579(.a(s_147), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1580(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1581(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1582(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2829(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2830(.a(gate67inter0), .b(s_326), .O(gate67inter1));
  and2  gate2831(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2832(.a(s_326), .O(gate67inter3));
  inv1  gate2833(.a(s_327), .O(gate67inter4));
  nand2 gate2834(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2835(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2836(.a(G27), .O(gate67inter7));
  inv1  gate2837(.a(G305), .O(gate67inter8));
  nand2 gate2838(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2839(.a(s_327), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2840(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2841(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2842(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate3081(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate3082(.a(gate68inter0), .b(s_362), .O(gate68inter1));
  and2  gate3083(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate3084(.a(s_362), .O(gate68inter3));
  inv1  gate3085(.a(s_363), .O(gate68inter4));
  nand2 gate3086(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate3087(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate3088(.a(G28), .O(gate68inter7));
  inv1  gate3089(.a(G305), .O(gate68inter8));
  nand2 gate3090(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate3091(.a(s_363), .b(gate68inter3), .O(gate68inter10));
  nor2  gate3092(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate3093(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate3094(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate3235(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate3236(.a(gate69inter0), .b(s_384), .O(gate69inter1));
  and2  gate3237(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate3238(.a(s_384), .O(gate69inter3));
  inv1  gate3239(.a(s_385), .O(gate69inter4));
  nand2 gate3240(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate3241(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate3242(.a(G29), .O(gate69inter7));
  inv1  gate3243(.a(G308), .O(gate69inter8));
  nand2 gate3244(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate3245(.a(s_385), .b(gate69inter3), .O(gate69inter10));
  nor2  gate3246(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate3247(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate3248(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2045(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2046(.a(gate71inter0), .b(s_214), .O(gate71inter1));
  and2  gate2047(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2048(.a(s_214), .O(gate71inter3));
  inv1  gate2049(.a(s_215), .O(gate71inter4));
  nand2 gate2050(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2051(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2052(.a(G31), .O(gate71inter7));
  inv1  gate2053(.a(G311), .O(gate71inter8));
  nand2 gate2054(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2055(.a(s_215), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2056(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2057(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2058(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1289(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1290(.a(gate78inter0), .b(s_106), .O(gate78inter1));
  and2  gate1291(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1292(.a(s_106), .O(gate78inter3));
  inv1  gate1293(.a(s_107), .O(gate78inter4));
  nand2 gate1294(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1295(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1296(.a(G6), .O(gate78inter7));
  inv1  gate1297(.a(G320), .O(gate78inter8));
  nand2 gate1298(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1299(.a(s_107), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1300(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1301(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1302(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1107(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1108(.a(gate79inter0), .b(s_80), .O(gate79inter1));
  and2  gate1109(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1110(.a(s_80), .O(gate79inter3));
  inv1  gate1111(.a(s_81), .O(gate79inter4));
  nand2 gate1112(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1113(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1114(.a(G10), .O(gate79inter7));
  inv1  gate1115(.a(G323), .O(gate79inter8));
  nand2 gate1116(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1117(.a(s_81), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1118(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1119(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1120(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate3109(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate3110(.a(gate88inter0), .b(s_366), .O(gate88inter1));
  and2  gate3111(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate3112(.a(s_366), .O(gate88inter3));
  inv1  gate3113(.a(s_367), .O(gate88inter4));
  nand2 gate3114(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate3115(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate3116(.a(G16), .O(gate88inter7));
  inv1  gate3117(.a(G335), .O(gate88inter8));
  nand2 gate3118(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate3119(.a(s_367), .b(gate88inter3), .O(gate88inter10));
  nor2  gate3120(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate3121(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate3122(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2451(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2452(.a(gate89inter0), .b(s_272), .O(gate89inter1));
  and2  gate2453(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2454(.a(s_272), .O(gate89inter3));
  inv1  gate2455(.a(s_273), .O(gate89inter4));
  nand2 gate2456(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2457(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2458(.a(G17), .O(gate89inter7));
  inv1  gate2459(.a(G338), .O(gate89inter8));
  nand2 gate2460(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2461(.a(s_273), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2462(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2463(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2464(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate2773(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2774(.a(gate90inter0), .b(s_318), .O(gate90inter1));
  and2  gate2775(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2776(.a(s_318), .O(gate90inter3));
  inv1  gate2777(.a(s_319), .O(gate90inter4));
  nand2 gate2778(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2779(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2780(.a(G21), .O(gate90inter7));
  inv1  gate2781(.a(G338), .O(gate90inter8));
  nand2 gate2782(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2783(.a(s_319), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2784(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2785(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2786(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate3095(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate3096(.a(gate92inter0), .b(s_364), .O(gate92inter1));
  and2  gate3097(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate3098(.a(s_364), .O(gate92inter3));
  inv1  gate3099(.a(s_365), .O(gate92inter4));
  nand2 gate3100(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate3101(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate3102(.a(G29), .O(gate92inter7));
  inv1  gate3103(.a(G341), .O(gate92inter8));
  nand2 gate3104(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate3105(.a(s_365), .b(gate92inter3), .O(gate92inter10));
  nor2  gate3106(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate3107(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate3108(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2423(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2424(.a(gate94inter0), .b(s_268), .O(gate94inter1));
  and2  gate2425(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2426(.a(s_268), .O(gate94inter3));
  inv1  gate2427(.a(s_269), .O(gate94inter4));
  nand2 gate2428(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2429(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2430(.a(G22), .O(gate94inter7));
  inv1  gate2431(.a(G344), .O(gate94inter8));
  nand2 gate2432(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2433(.a(s_269), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2434(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2435(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2436(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1051(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1052(.a(gate96inter0), .b(s_72), .O(gate96inter1));
  and2  gate1053(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1054(.a(s_72), .O(gate96inter3));
  inv1  gate1055(.a(s_73), .O(gate96inter4));
  nand2 gate1056(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1057(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1058(.a(G30), .O(gate96inter7));
  inv1  gate1059(.a(G347), .O(gate96inter8));
  nand2 gate1060(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1061(.a(s_73), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1062(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1063(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1064(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2885(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2886(.a(gate97inter0), .b(s_334), .O(gate97inter1));
  and2  gate2887(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2888(.a(s_334), .O(gate97inter3));
  inv1  gate2889(.a(s_335), .O(gate97inter4));
  nand2 gate2890(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2891(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2892(.a(G19), .O(gate97inter7));
  inv1  gate2893(.a(G350), .O(gate97inter8));
  nand2 gate2894(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2895(.a(s_335), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2896(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2897(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2898(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate3165(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate3166(.a(gate98inter0), .b(s_374), .O(gate98inter1));
  and2  gate3167(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate3168(.a(s_374), .O(gate98inter3));
  inv1  gate3169(.a(s_375), .O(gate98inter4));
  nand2 gate3170(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate3171(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate3172(.a(G23), .O(gate98inter7));
  inv1  gate3173(.a(G350), .O(gate98inter8));
  nand2 gate3174(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate3175(.a(s_375), .b(gate98inter3), .O(gate98inter10));
  nor2  gate3176(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate3177(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate3178(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate3011(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate3012(.a(gate99inter0), .b(s_352), .O(gate99inter1));
  and2  gate3013(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate3014(.a(s_352), .O(gate99inter3));
  inv1  gate3015(.a(s_353), .O(gate99inter4));
  nand2 gate3016(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate3017(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate3018(.a(G27), .O(gate99inter7));
  inv1  gate3019(.a(G353), .O(gate99inter8));
  nand2 gate3020(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate3021(.a(s_353), .b(gate99inter3), .O(gate99inter10));
  nor2  gate3022(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate3023(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate3024(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate911(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate912(.a(gate102inter0), .b(s_52), .O(gate102inter1));
  and2  gate913(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate914(.a(s_52), .O(gate102inter3));
  inv1  gate915(.a(s_53), .O(gate102inter4));
  nand2 gate916(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate917(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate918(.a(G24), .O(gate102inter7));
  inv1  gate919(.a(G356), .O(gate102inter8));
  nand2 gate920(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate921(.a(s_53), .b(gate102inter3), .O(gate102inter10));
  nor2  gate922(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate923(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate924(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2535(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2536(.a(gate104inter0), .b(s_284), .O(gate104inter1));
  and2  gate2537(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2538(.a(s_284), .O(gate104inter3));
  inv1  gate2539(.a(s_285), .O(gate104inter4));
  nand2 gate2540(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2541(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2542(.a(G32), .O(gate104inter7));
  inv1  gate2543(.a(G359), .O(gate104inter8));
  nand2 gate2544(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2545(.a(s_285), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2546(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2547(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2548(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2479(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2480(.a(gate106inter0), .b(s_276), .O(gate106inter1));
  and2  gate2481(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2482(.a(s_276), .O(gate106inter3));
  inv1  gate2483(.a(s_277), .O(gate106inter4));
  nand2 gate2484(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2485(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2486(.a(G364), .O(gate106inter7));
  inv1  gate2487(.a(G365), .O(gate106inter8));
  nand2 gate2488(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2489(.a(s_277), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2490(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2491(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2492(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1471(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1472(.a(gate107inter0), .b(s_132), .O(gate107inter1));
  and2  gate1473(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1474(.a(s_132), .O(gate107inter3));
  inv1  gate1475(.a(s_133), .O(gate107inter4));
  nand2 gate1476(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1477(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1478(.a(G366), .O(gate107inter7));
  inv1  gate1479(.a(G367), .O(gate107inter8));
  nand2 gate1480(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1481(.a(s_133), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1482(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1483(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1484(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1555(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1556(.a(gate112inter0), .b(s_144), .O(gate112inter1));
  and2  gate1557(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1558(.a(s_144), .O(gate112inter3));
  inv1  gate1559(.a(s_145), .O(gate112inter4));
  nand2 gate1560(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1561(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1562(.a(G376), .O(gate112inter7));
  inv1  gate1563(.a(G377), .O(gate112inter8));
  nand2 gate1564(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1565(.a(s_145), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1566(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1567(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1568(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate603(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate604(.a(gate115inter0), .b(s_8), .O(gate115inter1));
  and2  gate605(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate606(.a(s_8), .O(gate115inter3));
  inv1  gate607(.a(s_9), .O(gate115inter4));
  nand2 gate608(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate609(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate610(.a(G382), .O(gate115inter7));
  inv1  gate611(.a(G383), .O(gate115inter8));
  nand2 gate612(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate613(.a(s_9), .b(gate115inter3), .O(gate115inter10));
  nor2  gate614(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate615(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate616(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate645(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate646(.a(gate116inter0), .b(s_14), .O(gate116inter1));
  and2  gate647(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate648(.a(s_14), .O(gate116inter3));
  inv1  gate649(.a(s_15), .O(gate116inter4));
  nand2 gate650(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate651(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate652(.a(G384), .O(gate116inter7));
  inv1  gate653(.a(G385), .O(gate116inter8));
  nand2 gate654(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate655(.a(s_15), .b(gate116inter3), .O(gate116inter10));
  nor2  gate656(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate657(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate658(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2591(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2592(.a(gate118inter0), .b(s_292), .O(gate118inter1));
  and2  gate2593(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2594(.a(s_292), .O(gate118inter3));
  inv1  gate2595(.a(s_293), .O(gate118inter4));
  nand2 gate2596(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2597(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2598(.a(G388), .O(gate118inter7));
  inv1  gate2599(.a(G389), .O(gate118inter8));
  nand2 gate2600(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2601(.a(s_293), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2602(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2603(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2604(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1121(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1122(.a(gate122inter0), .b(s_82), .O(gate122inter1));
  and2  gate1123(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1124(.a(s_82), .O(gate122inter3));
  inv1  gate1125(.a(s_83), .O(gate122inter4));
  nand2 gate1126(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1127(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1128(.a(G396), .O(gate122inter7));
  inv1  gate1129(.a(G397), .O(gate122inter8));
  nand2 gate1130(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1131(.a(s_83), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1132(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1133(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1134(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate855(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate856(.a(gate124inter0), .b(s_44), .O(gate124inter1));
  and2  gate857(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate858(.a(s_44), .O(gate124inter3));
  inv1  gate859(.a(s_45), .O(gate124inter4));
  nand2 gate860(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate861(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate862(.a(G400), .O(gate124inter7));
  inv1  gate863(.a(G401), .O(gate124inter8));
  nand2 gate864(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate865(.a(s_45), .b(gate124inter3), .O(gate124inter10));
  nor2  gate866(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate867(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate868(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1443(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1444(.a(gate125inter0), .b(s_128), .O(gate125inter1));
  and2  gate1445(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1446(.a(s_128), .O(gate125inter3));
  inv1  gate1447(.a(s_129), .O(gate125inter4));
  nand2 gate1448(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1449(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1450(.a(G402), .O(gate125inter7));
  inv1  gate1451(.a(G403), .O(gate125inter8));
  nand2 gate1452(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1453(.a(s_129), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1454(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1455(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1456(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate813(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate814(.a(gate127inter0), .b(s_38), .O(gate127inter1));
  and2  gate815(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate816(.a(s_38), .O(gate127inter3));
  inv1  gate817(.a(s_39), .O(gate127inter4));
  nand2 gate818(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate819(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate820(.a(G406), .O(gate127inter7));
  inv1  gate821(.a(G407), .O(gate127inter8));
  nand2 gate822(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate823(.a(s_39), .b(gate127inter3), .O(gate127inter10));
  nor2  gate824(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate825(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate826(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2717(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2718(.a(gate129inter0), .b(s_310), .O(gate129inter1));
  and2  gate2719(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2720(.a(s_310), .O(gate129inter3));
  inv1  gate2721(.a(s_311), .O(gate129inter4));
  nand2 gate2722(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2723(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2724(.a(G410), .O(gate129inter7));
  inv1  gate2725(.a(G411), .O(gate129inter8));
  nand2 gate2726(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2727(.a(s_311), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2728(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2729(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2730(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate2339(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2340(.a(gate133inter0), .b(s_256), .O(gate133inter1));
  and2  gate2341(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2342(.a(s_256), .O(gate133inter3));
  inv1  gate2343(.a(s_257), .O(gate133inter4));
  nand2 gate2344(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2345(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2346(.a(G418), .O(gate133inter7));
  inv1  gate2347(.a(G419), .O(gate133inter8));
  nand2 gate2348(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2349(.a(s_257), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2350(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2351(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2352(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate3067(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate3068(.a(gate136inter0), .b(s_360), .O(gate136inter1));
  and2  gate3069(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate3070(.a(s_360), .O(gate136inter3));
  inv1  gate3071(.a(s_361), .O(gate136inter4));
  nand2 gate3072(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate3073(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate3074(.a(G424), .O(gate136inter7));
  inv1  gate3075(.a(G425), .O(gate136inter8));
  nand2 gate3076(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate3077(.a(s_361), .b(gate136inter3), .O(gate136inter10));
  nor2  gate3078(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate3079(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate3080(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2759(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2760(.a(gate138inter0), .b(s_316), .O(gate138inter1));
  and2  gate2761(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2762(.a(s_316), .O(gate138inter3));
  inv1  gate2763(.a(s_317), .O(gate138inter4));
  nand2 gate2764(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2765(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2766(.a(G432), .O(gate138inter7));
  inv1  gate2767(.a(G435), .O(gate138inter8));
  nand2 gate2768(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2769(.a(s_317), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2770(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2771(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2772(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1779(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1780(.a(gate139inter0), .b(s_176), .O(gate139inter1));
  and2  gate1781(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1782(.a(s_176), .O(gate139inter3));
  inv1  gate1783(.a(s_177), .O(gate139inter4));
  nand2 gate1784(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1785(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1786(.a(G438), .O(gate139inter7));
  inv1  gate1787(.a(G441), .O(gate139inter8));
  nand2 gate1788(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1789(.a(s_177), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1790(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1791(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1792(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate953(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate954(.a(gate140inter0), .b(s_58), .O(gate140inter1));
  and2  gate955(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate956(.a(s_58), .O(gate140inter3));
  inv1  gate957(.a(s_59), .O(gate140inter4));
  nand2 gate958(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate959(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate960(.a(G444), .O(gate140inter7));
  inv1  gate961(.a(G447), .O(gate140inter8));
  nand2 gate962(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate963(.a(s_59), .b(gate140inter3), .O(gate140inter10));
  nor2  gate964(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate965(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate966(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1737(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1738(.a(gate142inter0), .b(s_170), .O(gate142inter1));
  and2  gate1739(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1740(.a(s_170), .O(gate142inter3));
  inv1  gate1741(.a(s_171), .O(gate142inter4));
  nand2 gate1742(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1743(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1744(.a(G456), .O(gate142inter7));
  inv1  gate1745(.a(G459), .O(gate142inter8));
  nand2 gate1746(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1747(.a(s_171), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1748(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1749(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1750(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2073(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2074(.a(gate144inter0), .b(s_218), .O(gate144inter1));
  and2  gate2075(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2076(.a(s_218), .O(gate144inter3));
  inv1  gate2077(.a(s_219), .O(gate144inter4));
  nand2 gate2078(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2079(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2080(.a(G468), .O(gate144inter7));
  inv1  gate2081(.a(G471), .O(gate144inter8));
  nand2 gate2082(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2083(.a(s_219), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2084(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2085(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2086(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1429(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1430(.a(gate145inter0), .b(s_126), .O(gate145inter1));
  and2  gate1431(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1432(.a(s_126), .O(gate145inter3));
  inv1  gate1433(.a(s_127), .O(gate145inter4));
  nand2 gate1434(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1435(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1436(.a(G474), .O(gate145inter7));
  inv1  gate1437(.a(G477), .O(gate145inter8));
  nand2 gate1438(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1439(.a(s_127), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1440(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1441(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1442(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate547(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate548(.a(gate146inter0), .b(s_0), .O(gate146inter1));
  and2  gate549(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate550(.a(s_0), .O(gate146inter3));
  inv1  gate551(.a(s_1), .O(gate146inter4));
  nand2 gate552(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate553(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate554(.a(G480), .O(gate146inter7));
  inv1  gate555(.a(G483), .O(gate146inter8));
  nand2 gate556(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate557(.a(s_1), .b(gate146inter3), .O(gate146inter10));
  nor2  gate558(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate559(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate560(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate743(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate744(.a(gate150inter0), .b(s_28), .O(gate150inter1));
  and2  gate745(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate746(.a(s_28), .O(gate150inter3));
  inv1  gate747(.a(s_29), .O(gate150inter4));
  nand2 gate748(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate749(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate750(.a(G504), .O(gate150inter7));
  inv1  gate751(.a(G507), .O(gate150inter8));
  nand2 gate752(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate753(.a(s_29), .b(gate150inter3), .O(gate150inter10));
  nor2  gate754(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate755(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate756(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1793(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1794(.a(gate154inter0), .b(s_178), .O(gate154inter1));
  and2  gate1795(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1796(.a(s_178), .O(gate154inter3));
  inv1  gate1797(.a(s_179), .O(gate154inter4));
  nand2 gate1798(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1799(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1800(.a(G429), .O(gate154inter7));
  inv1  gate1801(.a(G522), .O(gate154inter8));
  nand2 gate1802(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1803(.a(s_179), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1804(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1805(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1806(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1765(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1766(.a(gate155inter0), .b(s_174), .O(gate155inter1));
  and2  gate1767(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1768(.a(s_174), .O(gate155inter3));
  inv1  gate1769(.a(s_175), .O(gate155inter4));
  nand2 gate1770(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1771(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1772(.a(G432), .O(gate155inter7));
  inv1  gate1773(.a(G525), .O(gate155inter8));
  nand2 gate1774(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1775(.a(s_175), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1776(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1777(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1778(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2549(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2550(.a(gate156inter0), .b(s_286), .O(gate156inter1));
  and2  gate2551(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2552(.a(s_286), .O(gate156inter3));
  inv1  gate2553(.a(s_287), .O(gate156inter4));
  nand2 gate2554(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2555(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2556(.a(G435), .O(gate156inter7));
  inv1  gate2557(.a(G525), .O(gate156inter8));
  nand2 gate2558(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2559(.a(s_287), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2560(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2561(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2562(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1023(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1024(.a(gate158inter0), .b(s_68), .O(gate158inter1));
  and2  gate1025(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1026(.a(s_68), .O(gate158inter3));
  inv1  gate1027(.a(s_69), .O(gate158inter4));
  nand2 gate1028(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1029(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1030(.a(G441), .O(gate158inter7));
  inv1  gate1031(.a(G528), .O(gate158inter8));
  nand2 gate1032(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1033(.a(s_69), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1034(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1035(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1036(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2199(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2200(.a(gate160inter0), .b(s_236), .O(gate160inter1));
  and2  gate2201(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2202(.a(s_236), .O(gate160inter3));
  inv1  gate2203(.a(s_237), .O(gate160inter4));
  nand2 gate2204(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2205(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2206(.a(G447), .O(gate160inter7));
  inv1  gate2207(.a(G531), .O(gate160inter8));
  nand2 gate2208(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2209(.a(s_237), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2210(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2211(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2212(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate3305(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate3306(.a(gate161inter0), .b(s_394), .O(gate161inter1));
  and2  gate3307(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate3308(.a(s_394), .O(gate161inter3));
  inv1  gate3309(.a(s_395), .O(gate161inter4));
  nand2 gate3310(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate3311(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate3312(.a(G450), .O(gate161inter7));
  inv1  gate3313(.a(G534), .O(gate161inter8));
  nand2 gate3314(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate3315(.a(s_395), .b(gate161inter3), .O(gate161inter10));
  nor2  gate3316(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate3317(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate3318(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1177(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1178(.a(gate162inter0), .b(s_90), .O(gate162inter1));
  and2  gate1179(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1180(.a(s_90), .O(gate162inter3));
  inv1  gate1181(.a(s_91), .O(gate162inter4));
  nand2 gate1182(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1183(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1184(.a(G453), .O(gate162inter7));
  inv1  gate1185(.a(G534), .O(gate162inter8));
  nand2 gate1186(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1187(.a(s_91), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1188(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1189(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1190(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2815(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2816(.a(gate163inter0), .b(s_324), .O(gate163inter1));
  and2  gate2817(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2818(.a(s_324), .O(gate163inter3));
  inv1  gate2819(.a(s_325), .O(gate163inter4));
  nand2 gate2820(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2821(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2822(.a(G456), .O(gate163inter7));
  inv1  gate2823(.a(G537), .O(gate163inter8));
  nand2 gate2824(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2825(.a(s_325), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2826(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2827(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2828(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2367(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2368(.a(gate164inter0), .b(s_260), .O(gate164inter1));
  and2  gate2369(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2370(.a(s_260), .O(gate164inter3));
  inv1  gate2371(.a(s_261), .O(gate164inter4));
  nand2 gate2372(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2373(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2374(.a(G459), .O(gate164inter7));
  inv1  gate2375(.a(G537), .O(gate164inter8));
  nand2 gate2376(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2377(.a(s_261), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2378(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2379(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2380(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1863(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1864(.a(gate167inter0), .b(s_188), .O(gate167inter1));
  and2  gate1865(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1866(.a(s_188), .O(gate167inter3));
  inv1  gate1867(.a(s_189), .O(gate167inter4));
  nand2 gate1868(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1869(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1870(.a(G468), .O(gate167inter7));
  inv1  gate1871(.a(G543), .O(gate167inter8));
  nand2 gate1872(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1873(.a(s_189), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1874(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1875(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1876(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1961(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1962(.a(gate168inter0), .b(s_202), .O(gate168inter1));
  and2  gate1963(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1964(.a(s_202), .O(gate168inter3));
  inv1  gate1965(.a(s_203), .O(gate168inter4));
  nand2 gate1966(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1967(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1968(.a(G471), .O(gate168inter7));
  inv1  gate1969(.a(G543), .O(gate168inter8));
  nand2 gate1970(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1971(.a(s_203), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1972(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1973(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1974(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2465(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2466(.a(gate170inter0), .b(s_274), .O(gate170inter1));
  and2  gate2467(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2468(.a(s_274), .O(gate170inter3));
  inv1  gate2469(.a(s_275), .O(gate170inter4));
  nand2 gate2470(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2471(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2472(.a(G477), .O(gate170inter7));
  inv1  gate2473(.a(G546), .O(gate170inter8));
  nand2 gate2474(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2475(.a(s_275), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2476(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2477(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2478(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1415(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1416(.a(gate171inter0), .b(s_124), .O(gate171inter1));
  and2  gate1417(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1418(.a(s_124), .O(gate171inter3));
  inv1  gate1419(.a(s_125), .O(gate171inter4));
  nand2 gate1420(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1421(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1422(.a(G480), .O(gate171inter7));
  inv1  gate1423(.a(G549), .O(gate171inter8));
  nand2 gate1424(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1425(.a(s_125), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1426(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1427(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1428(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2129(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2130(.a(gate172inter0), .b(s_226), .O(gate172inter1));
  and2  gate2131(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2132(.a(s_226), .O(gate172inter3));
  inv1  gate2133(.a(s_227), .O(gate172inter4));
  nand2 gate2134(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2135(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2136(.a(G483), .O(gate172inter7));
  inv1  gate2137(.a(G549), .O(gate172inter8));
  nand2 gate2138(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2139(.a(s_227), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2140(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2141(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2142(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2395(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2396(.a(gate175inter0), .b(s_264), .O(gate175inter1));
  and2  gate2397(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2398(.a(s_264), .O(gate175inter3));
  inv1  gate2399(.a(s_265), .O(gate175inter4));
  nand2 gate2400(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2401(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2402(.a(G492), .O(gate175inter7));
  inv1  gate2403(.a(G555), .O(gate175inter8));
  nand2 gate2404(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2405(.a(s_265), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2406(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2407(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2408(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1695(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1696(.a(gate176inter0), .b(s_164), .O(gate176inter1));
  and2  gate1697(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1698(.a(s_164), .O(gate176inter3));
  inv1  gate1699(.a(s_165), .O(gate176inter4));
  nand2 gate1700(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1701(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1702(.a(G495), .O(gate176inter7));
  inv1  gate1703(.a(G555), .O(gate176inter8));
  nand2 gate1704(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1705(.a(s_165), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1706(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1707(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1708(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate3319(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate3320(.a(gate177inter0), .b(s_396), .O(gate177inter1));
  and2  gate3321(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate3322(.a(s_396), .O(gate177inter3));
  inv1  gate3323(.a(s_397), .O(gate177inter4));
  nand2 gate3324(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate3325(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate3326(.a(G498), .O(gate177inter7));
  inv1  gate3327(.a(G558), .O(gate177inter8));
  nand2 gate3328(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate3329(.a(s_397), .b(gate177inter3), .O(gate177inter10));
  nor2  gate3330(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate3331(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate3332(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate2521(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2522(.a(gate178inter0), .b(s_282), .O(gate178inter1));
  and2  gate2523(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2524(.a(s_282), .O(gate178inter3));
  inv1  gate2525(.a(s_283), .O(gate178inter4));
  nand2 gate2526(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2527(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2528(.a(G501), .O(gate178inter7));
  inv1  gate2529(.a(G558), .O(gate178inter8));
  nand2 gate2530(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2531(.a(s_283), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2532(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2533(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2534(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate3053(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate3054(.a(gate179inter0), .b(s_358), .O(gate179inter1));
  and2  gate3055(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate3056(.a(s_358), .O(gate179inter3));
  inv1  gate3057(.a(s_359), .O(gate179inter4));
  nand2 gate3058(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate3059(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate3060(.a(G504), .O(gate179inter7));
  inv1  gate3061(.a(G561), .O(gate179inter8));
  nand2 gate3062(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate3063(.a(s_359), .b(gate179inter3), .O(gate179inter10));
  nor2  gate3064(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate3065(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate3066(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate3347(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate3348(.a(gate180inter0), .b(s_400), .O(gate180inter1));
  and2  gate3349(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate3350(.a(s_400), .O(gate180inter3));
  inv1  gate3351(.a(s_401), .O(gate180inter4));
  nand2 gate3352(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate3353(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate3354(.a(G507), .O(gate180inter7));
  inv1  gate3355(.a(G561), .O(gate180inter8));
  nand2 gate3356(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate3357(.a(s_401), .b(gate180inter3), .O(gate180inter10));
  nor2  gate3358(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate3359(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate3360(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2955(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2956(.a(gate182inter0), .b(s_344), .O(gate182inter1));
  and2  gate2957(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2958(.a(s_344), .O(gate182inter3));
  inv1  gate2959(.a(s_345), .O(gate182inter4));
  nand2 gate2960(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2961(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2962(.a(G513), .O(gate182inter7));
  inv1  gate2963(.a(G564), .O(gate182inter8));
  nand2 gate2964(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2965(.a(s_345), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2966(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2967(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2968(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1359(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1360(.a(gate183inter0), .b(s_116), .O(gate183inter1));
  and2  gate1361(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1362(.a(s_116), .O(gate183inter3));
  inv1  gate1363(.a(s_117), .O(gate183inter4));
  nand2 gate1364(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1365(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1366(.a(G516), .O(gate183inter7));
  inv1  gate1367(.a(G567), .O(gate183inter8));
  nand2 gate1368(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1369(.a(s_117), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1370(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1371(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1372(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2297(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2298(.a(gate190inter0), .b(s_250), .O(gate190inter1));
  and2  gate2299(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2300(.a(s_250), .O(gate190inter3));
  inv1  gate2301(.a(s_251), .O(gate190inter4));
  nand2 gate2302(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2303(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2304(.a(G580), .O(gate190inter7));
  inv1  gate2305(.a(G581), .O(gate190inter8));
  nand2 gate2306(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2307(.a(s_251), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2308(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2309(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2310(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1597(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1598(.a(gate191inter0), .b(s_150), .O(gate191inter1));
  and2  gate1599(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1600(.a(s_150), .O(gate191inter3));
  inv1  gate1601(.a(s_151), .O(gate191inter4));
  nand2 gate1602(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1603(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1604(.a(G582), .O(gate191inter7));
  inv1  gate1605(.a(G583), .O(gate191inter8));
  nand2 gate1606(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1607(.a(s_151), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1608(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1609(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1610(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2927(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2928(.a(gate194inter0), .b(s_340), .O(gate194inter1));
  and2  gate2929(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2930(.a(s_340), .O(gate194inter3));
  inv1  gate2931(.a(s_341), .O(gate194inter4));
  nand2 gate2932(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2933(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2934(.a(G588), .O(gate194inter7));
  inv1  gate2935(.a(G589), .O(gate194inter8));
  nand2 gate2936(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2937(.a(s_341), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2938(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2939(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2940(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2563(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2564(.a(gate198inter0), .b(s_288), .O(gate198inter1));
  and2  gate2565(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2566(.a(s_288), .O(gate198inter3));
  inv1  gate2567(.a(s_289), .O(gate198inter4));
  nand2 gate2568(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2569(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2570(.a(G596), .O(gate198inter7));
  inv1  gate2571(.a(G597), .O(gate198inter8));
  nand2 gate2572(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2573(.a(s_289), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2574(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2575(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2576(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2171(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2172(.a(gate200inter0), .b(s_232), .O(gate200inter1));
  and2  gate2173(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2174(.a(s_232), .O(gate200inter3));
  inv1  gate2175(.a(s_233), .O(gate200inter4));
  nand2 gate2176(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2177(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2178(.a(G600), .O(gate200inter7));
  inv1  gate2179(.a(G601), .O(gate200inter8));
  nand2 gate2180(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2181(.a(s_233), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2182(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2183(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2184(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1667(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1668(.a(gate201inter0), .b(s_160), .O(gate201inter1));
  and2  gate1669(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1670(.a(s_160), .O(gate201inter3));
  inv1  gate1671(.a(s_161), .O(gate201inter4));
  nand2 gate1672(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1673(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1674(.a(G602), .O(gate201inter7));
  inv1  gate1675(.a(G607), .O(gate201inter8));
  nand2 gate1676(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1677(.a(s_161), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1678(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1679(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1680(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate3123(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate3124(.a(gate203inter0), .b(s_368), .O(gate203inter1));
  and2  gate3125(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate3126(.a(s_368), .O(gate203inter3));
  inv1  gate3127(.a(s_369), .O(gate203inter4));
  nand2 gate3128(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate3129(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate3130(.a(G602), .O(gate203inter7));
  inv1  gate3131(.a(G612), .O(gate203inter8));
  nand2 gate3132(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate3133(.a(s_369), .b(gate203inter3), .O(gate203inter10));
  nor2  gate3134(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate3135(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate3136(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1513(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1514(.a(gate205inter0), .b(s_138), .O(gate205inter1));
  and2  gate1515(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1516(.a(s_138), .O(gate205inter3));
  inv1  gate1517(.a(s_139), .O(gate205inter4));
  nand2 gate1518(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1519(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1520(.a(G622), .O(gate205inter7));
  inv1  gate1521(.a(G627), .O(gate205inter8));
  nand2 gate1522(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1523(.a(s_139), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1524(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1525(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1526(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2801(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2802(.a(gate206inter0), .b(s_322), .O(gate206inter1));
  and2  gate2803(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2804(.a(s_322), .O(gate206inter3));
  inv1  gate2805(.a(s_323), .O(gate206inter4));
  nand2 gate2806(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2807(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2808(.a(G632), .O(gate206inter7));
  inv1  gate2809(.a(G637), .O(gate206inter8));
  nand2 gate2810(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2811(.a(s_323), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2812(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2813(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2814(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate3179(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate3180(.a(gate207inter0), .b(s_376), .O(gate207inter1));
  and2  gate3181(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate3182(.a(s_376), .O(gate207inter3));
  inv1  gate3183(.a(s_377), .O(gate207inter4));
  nand2 gate3184(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate3185(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate3186(.a(G622), .O(gate207inter7));
  inv1  gate3187(.a(G632), .O(gate207inter8));
  nand2 gate3188(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate3189(.a(s_377), .b(gate207inter3), .O(gate207inter10));
  nor2  gate3190(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate3191(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate3192(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate3277(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate3278(.a(gate208inter0), .b(s_390), .O(gate208inter1));
  and2  gate3279(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate3280(.a(s_390), .O(gate208inter3));
  inv1  gate3281(.a(s_391), .O(gate208inter4));
  nand2 gate3282(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate3283(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate3284(.a(G627), .O(gate208inter7));
  inv1  gate3285(.a(G637), .O(gate208inter8));
  nand2 gate3286(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate3287(.a(s_391), .b(gate208inter3), .O(gate208inter10));
  nor2  gate3288(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate3289(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate3290(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1373(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1374(.a(gate209inter0), .b(s_118), .O(gate209inter1));
  and2  gate1375(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1376(.a(s_118), .O(gate209inter3));
  inv1  gate1377(.a(s_119), .O(gate209inter4));
  nand2 gate1378(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1379(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1380(.a(G602), .O(gate209inter7));
  inv1  gate1381(.a(G666), .O(gate209inter8));
  nand2 gate1382(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1383(.a(s_119), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1384(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1385(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1386(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate757(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate758(.a(gate210inter0), .b(s_30), .O(gate210inter1));
  and2  gate759(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate760(.a(s_30), .O(gate210inter3));
  inv1  gate761(.a(s_31), .O(gate210inter4));
  nand2 gate762(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate763(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate764(.a(G607), .O(gate210inter7));
  inv1  gate765(.a(G666), .O(gate210inter8));
  nand2 gate766(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate767(.a(s_31), .b(gate210inter3), .O(gate210inter10));
  nor2  gate768(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate769(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate770(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1905(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1906(.a(gate214inter0), .b(s_194), .O(gate214inter1));
  and2  gate1907(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1908(.a(s_194), .O(gate214inter3));
  inv1  gate1909(.a(s_195), .O(gate214inter4));
  nand2 gate1910(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1911(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1912(.a(G612), .O(gate214inter7));
  inv1  gate1913(.a(G672), .O(gate214inter8));
  nand2 gate1914(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1915(.a(s_195), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1916(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1917(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1918(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1975(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1976(.a(gate220inter0), .b(s_204), .O(gate220inter1));
  and2  gate1977(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1978(.a(s_204), .O(gate220inter3));
  inv1  gate1979(.a(s_205), .O(gate220inter4));
  nand2 gate1980(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1981(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1982(.a(G637), .O(gate220inter7));
  inv1  gate1983(.a(G681), .O(gate220inter8));
  nand2 gate1984(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1985(.a(s_205), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1986(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1987(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1988(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2913(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2914(.a(gate223inter0), .b(s_338), .O(gate223inter1));
  and2  gate2915(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2916(.a(s_338), .O(gate223inter3));
  inv1  gate2917(.a(s_339), .O(gate223inter4));
  nand2 gate2918(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2919(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2920(.a(G627), .O(gate223inter7));
  inv1  gate2921(.a(G687), .O(gate223inter8));
  nand2 gate2922(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2923(.a(s_339), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2924(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2925(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2926(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1877(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1878(.a(gate225inter0), .b(s_190), .O(gate225inter1));
  and2  gate1879(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1880(.a(s_190), .O(gate225inter3));
  inv1  gate1881(.a(s_191), .O(gate225inter4));
  nand2 gate1882(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1883(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1884(.a(G690), .O(gate225inter7));
  inv1  gate1885(.a(G691), .O(gate225inter8));
  nand2 gate1886(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1887(.a(s_191), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1888(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1889(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1890(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1387(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1388(.a(gate226inter0), .b(s_120), .O(gate226inter1));
  and2  gate1389(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1390(.a(s_120), .O(gate226inter3));
  inv1  gate1391(.a(s_121), .O(gate226inter4));
  nand2 gate1392(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1393(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1394(.a(G692), .O(gate226inter7));
  inv1  gate1395(.a(G693), .O(gate226inter8));
  nand2 gate1396(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1397(.a(s_121), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1398(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1399(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1400(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate827(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate828(.a(gate227inter0), .b(s_40), .O(gate227inter1));
  and2  gate829(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate830(.a(s_40), .O(gate227inter3));
  inv1  gate831(.a(s_41), .O(gate227inter4));
  nand2 gate832(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate833(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate834(.a(G694), .O(gate227inter7));
  inv1  gate835(.a(G695), .O(gate227inter8));
  nand2 gate836(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate837(.a(s_41), .b(gate227inter3), .O(gate227inter10));
  nor2  gate838(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate839(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate840(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2115(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2116(.a(gate229inter0), .b(s_224), .O(gate229inter1));
  and2  gate2117(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2118(.a(s_224), .O(gate229inter3));
  inv1  gate2119(.a(s_225), .O(gate229inter4));
  nand2 gate2120(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2121(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2122(.a(G698), .O(gate229inter7));
  inv1  gate2123(.a(G699), .O(gate229inter8));
  nand2 gate2124(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2125(.a(s_225), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2126(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2127(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2128(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1709(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1710(.a(gate231inter0), .b(s_166), .O(gate231inter1));
  and2  gate1711(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1712(.a(s_166), .O(gate231inter3));
  inv1  gate1713(.a(s_167), .O(gate231inter4));
  nand2 gate1714(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1715(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1716(.a(G702), .O(gate231inter7));
  inv1  gate1717(.a(G703), .O(gate231inter8));
  nand2 gate1718(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1719(.a(s_167), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1720(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1721(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1722(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1499(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1500(.a(gate233inter0), .b(s_136), .O(gate233inter1));
  and2  gate1501(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1502(.a(s_136), .O(gate233inter3));
  inv1  gate1503(.a(s_137), .O(gate233inter4));
  nand2 gate1504(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1505(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1506(.a(G242), .O(gate233inter7));
  inv1  gate1507(.a(G718), .O(gate233inter8));
  nand2 gate1508(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1509(.a(s_137), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1510(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1511(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1512(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2731(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2732(.a(gate234inter0), .b(s_312), .O(gate234inter1));
  and2  gate2733(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2734(.a(s_312), .O(gate234inter3));
  inv1  gate2735(.a(s_313), .O(gate234inter4));
  nand2 gate2736(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2737(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2738(.a(G245), .O(gate234inter7));
  inv1  gate2739(.a(G721), .O(gate234inter8));
  nand2 gate2740(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2741(.a(s_313), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2742(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2743(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2744(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1541(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1542(.a(gate236inter0), .b(s_142), .O(gate236inter1));
  and2  gate1543(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1544(.a(s_142), .O(gate236inter3));
  inv1  gate1545(.a(s_143), .O(gate236inter4));
  nand2 gate1546(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1547(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1548(.a(G251), .O(gate236inter7));
  inv1  gate1549(.a(G727), .O(gate236inter8));
  nand2 gate1550(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1551(.a(s_143), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1552(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1553(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1554(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate617(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate618(.a(gate238inter0), .b(s_10), .O(gate238inter1));
  and2  gate619(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate620(.a(s_10), .O(gate238inter3));
  inv1  gate621(.a(s_11), .O(gate238inter4));
  nand2 gate622(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate623(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate624(.a(G257), .O(gate238inter7));
  inv1  gate625(.a(G709), .O(gate238inter8));
  nand2 gate626(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate627(.a(s_11), .b(gate238inter3), .O(gate238inter10));
  nor2  gate628(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate629(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate630(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate3221(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate3222(.a(gate239inter0), .b(s_382), .O(gate239inter1));
  and2  gate3223(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate3224(.a(s_382), .O(gate239inter3));
  inv1  gate3225(.a(s_383), .O(gate239inter4));
  nand2 gate3226(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate3227(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate3228(.a(G260), .O(gate239inter7));
  inv1  gate3229(.a(G712), .O(gate239inter8));
  nand2 gate3230(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate3231(.a(s_383), .b(gate239inter3), .O(gate239inter10));
  nor2  gate3232(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate3233(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate3234(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate883(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate884(.a(gate240inter0), .b(s_48), .O(gate240inter1));
  and2  gate885(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate886(.a(s_48), .O(gate240inter3));
  inv1  gate887(.a(s_49), .O(gate240inter4));
  nand2 gate888(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate889(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate890(.a(G263), .O(gate240inter7));
  inv1  gate891(.a(G715), .O(gate240inter8));
  nand2 gate892(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate893(.a(s_49), .b(gate240inter3), .O(gate240inter10));
  nor2  gate894(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate895(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate896(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate673(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate674(.a(gate241inter0), .b(s_18), .O(gate241inter1));
  and2  gate675(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate676(.a(s_18), .O(gate241inter3));
  inv1  gate677(.a(s_19), .O(gate241inter4));
  nand2 gate678(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate679(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate680(.a(G242), .O(gate241inter7));
  inv1  gate681(.a(G730), .O(gate241inter8));
  nand2 gate682(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate683(.a(s_19), .b(gate241inter3), .O(gate241inter10));
  nor2  gate684(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate685(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate686(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2143(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2144(.a(gate243inter0), .b(s_228), .O(gate243inter1));
  and2  gate2145(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2146(.a(s_228), .O(gate243inter3));
  inv1  gate2147(.a(s_229), .O(gate243inter4));
  nand2 gate2148(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2149(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2150(.a(G245), .O(gate243inter7));
  inv1  gate2151(.a(G733), .O(gate243inter8));
  nand2 gate2152(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2153(.a(s_229), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2154(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2155(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2156(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate3151(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate3152(.a(gate245inter0), .b(s_372), .O(gate245inter1));
  and2  gate3153(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate3154(.a(s_372), .O(gate245inter3));
  inv1  gate3155(.a(s_373), .O(gate245inter4));
  nand2 gate3156(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate3157(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate3158(.a(G248), .O(gate245inter7));
  inv1  gate3159(.a(G736), .O(gate245inter8));
  nand2 gate3160(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate3161(.a(s_373), .b(gate245inter3), .O(gate245inter10));
  nor2  gate3162(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate3163(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate3164(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1485(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1486(.a(gate247inter0), .b(s_134), .O(gate247inter1));
  and2  gate1487(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1488(.a(s_134), .O(gate247inter3));
  inv1  gate1489(.a(s_135), .O(gate247inter4));
  nand2 gate1490(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1491(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1492(.a(G251), .O(gate247inter7));
  inv1  gate1493(.a(G739), .O(gate247inter8));
  nand2 gate1494(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1495(.a(s_135), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1496(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1497(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1498(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1149(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1150(.a(gate250inter0), .b(s_86), .O(gate250inter1));
  and2  gate1151(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1152(.a(s_86), .O(gate250inter3));
  inv1  gate1153(.a(s_87), .O(gate250inter4));
  nand2 gate1154(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1155(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1156(.a(G706), .O(gate250inter7));
  inv1  gate1157(.a(G742), .O(gate250inter8));
  nand2 gate1158(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1159(.a(s_87), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1160(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1161(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1162(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2787(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2788(.a(gate251inter0), .b(s_320), .O(gate251inter1));
  and2  gate2789(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2790(.a(s_320), .O(gate251inter3));
  inv1  gate2791(.a(s_321), .O(gate251inter4));
  nand2 gate2792(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2793(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2794(.a(G257), .O(gate251inter7));
  inv1  gate2795(.a(G745), .O(gate251inter8));
  nand2 gate2796(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2797(.a(s_321), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2798(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2799(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2800(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate2843(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2844(.a(gate252inter0), .b(s_328), .O(gate252inter1));
  and2  gate2845(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2846(.a(s_328), .O(gate252inter3));
  inv1  gate2847(.a(s_329), .O(gate252inter4));
  nand2 gate2848(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2849(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2850(.a(G709), .O(gate252inter7));
  inv1  gate2851(.a(G745), .O(gate252inter8));
  nand2 gate2852(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2853(.a(s_329), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2854(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2855(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2856(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate939(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate940(.a(gate254inter0), .b(s_56), .O(gate254inter1));
  and2  gate941(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate942(.a(s_56), .O(gate254inter3));
  inv1  gate943(.a(s_57), .O(gate254inter4));
  nand2 gate944(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate945(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate946(.a(G712), .O(gate254inter7));
  inv1  gate947(.a(G748), .O(gate254inter8));
  nand2 gate948(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate949(.a(s_57), .b(gate254inter3), .O(gate254inter10));
  nor2  gate950(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate951(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate952(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2577(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2578(.a(gate257inter0), .b(s_290), .O(gate257inter1));
  and2  gate2579(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2580(.a(s_290), .O(gate257inter3));
  inv1  gate2581(.a(s_291), .O(gate257inter4));
  nand2 gate2582(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2583(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2584(.a(G754), .O(gate257inter7));
  inv1  gate2585(.a(G755), .O(gate257inter8));
  nand2 gate2586(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2587(.a(s_291), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2588(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2589(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2590(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1317(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1318(.a(gate258inter0), .b(s_110), .O(gate258inter1));
  and2  gate1319(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1320(.a(s_110), .O(gate258inter3));
  inv1  gate1321(.a(s_111), .O(gate258inter4));
  nand2 gate1322(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1323(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1324(.a(G756), .O(gate258inter7));
  inv1  gate1325(.a(G757), .O(gate258inter8));
  nand2 gate1326(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1327(.a(s_111), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1328(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1329(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1330(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate3039(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate3040(.a(gate259inter0), .b(s_356), .O(gate259inter1));
  and2  gate3041(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate3042(.a(s_356), .O(gate259inter3));
  inv1  gate3043(.a(s_357), .O(gate259inter4));
  nand2 gate3044(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate3045(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate3046(.a(G758), .O(gate259inter7));
  inv1  gate3047(.a(G759), .O(gate259inter8));
  nand2 gate3048(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate3049(.a(s_357), .b(gate259inter3), .O(gate259inter10));
  nor2  gate3050(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate3051(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate3052(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1583(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1584(.a(gate260inter0), .b(s_148), .O(gate260inter1));
  and2  gate1585(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1586(.a(s_148), .O(gate260inter3));
  inv1  gate1587(.a(s_149), .O(gate260inter4));
  nand2 gate1588(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1589(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1590(.a(G760), .O(gate260inter7));
  inv1  gate1591(.a(G761), .O(gate260inter8));
  nand2 gate1592(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1593(.a(s_149), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1594(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1595(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1596(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1849(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1850(.a(gate261inter0), .b(s_186), .O(gate261inter1));
  and2  gate1851(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1852(.a(s_186), .O(gate261inter3));
  inv1  gate1853(.a(s_187), .O(gate261inter4));
  nand2 gate1854(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1855(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1856(.a(G762), .O(gate261inter7));
  inv1  gate1857(.a(G763), .O(gate261inter8));
  nand2 gate1858(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1859(.a(s_187), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1860(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1861(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1862(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate729(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate730(.a(gate262inter0), .b(s_26), .O(gate262inter1));
  and2  gate731(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate732(.a(s_26), .O(gate262inter3));
  inv1  gate733(.a(s_27), .O(gate262inter4));
  nand2 gate734(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate735(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate736(.a(G764), .O(gate262inter7));
  inv1  gate737(.a(G765), .O(gate262inter8));
  nand2 gate738(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate739(.a(s_27), .b(gate262inter3), .O(gate262inter10));
  nor2  gate740(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate741(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate742(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate981(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate982(.a(gate263inter0), .b(s_62), .O(gate263inter1));
  and2  gate983(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate984(.a(s_62), .O(gate263inter3));
  inv1  gate985(.a(s_63), .O(gate263inter4));
  nand2 gate986(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate987(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate988(.a(G766), .O(gate263inter7));
  inv1  gate989(.a(G767), .O(gate263inter8));
  nand2 gate990(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate991(.a(s_63), .b(gate263inter3), .O(gate263inter10));
  nor2  gate992(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate993(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate994(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate659(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate660(.a(gate265inter0), .b(s_16), .O(gate265inter1));
  and2  gate661(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate662(.a(s_16), .O(gate265inter3));
  inv1  gate663(.a(s_17), .O(gate265inter4));
  nand2 gate664(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate665(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate666(.a(G642), .O(gate265inter7));
  inv1  gate667(.a(G770), .O(gate265inter8));
  nand2 gate668(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate669(.a(s_17), .b(gate265inter3), .O(gate265inter10));
  nor2  gate670(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate671(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate672(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate2311(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2312(.a(gate266inter0), .b(s_252), .O(gate266inter1));
  and2  gate2313(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2314(.a(s_252), .O(gate266inter3));
  inv1  gate2315(.a(s_253), .O(gate266inter4));
  nand2 gate2316(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2317(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2318(.a(G645), .O(gate266inter7));
  inv1  gate2319(.a(G773), .O(gate266inter8));
  nand2 gate2320(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2321(.a(s_253), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2322(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2323(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2324(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate925(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate926(.a(gate268inter0), .b(s_54), .O(gate268inter1));
  and2  gate927(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate928(.a(s_54), .O(gate268inter3));
  inv1  gate929(.a(s_55), .O(gate268inter4));
  nand2 gate930(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate931(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate932(.a(G651), .O(gate268inter7));
  inv1  gate933(.a(G779), .O(gate268inter8));
  nand2 gate934(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate935(.a(s_55), .b(gate268inter3), .O(gate268inter10));
  nor2  gate936(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate937(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate938(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2941(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2942(.a(gate269inter0), .b(s_342), .O(gate269inter1));
  and2  gate2943(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2944(.a(s_342), .O(gate269inter3));
  inv1  gate2945(.a(s_343), .O(gate269inter4));
  nand2 gate2946(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2947(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2948(.a(G654), .O(gate269inter7));
  inv1  gate2949(.a(G782), .O(gate269inter8));
  nand2 gate2950(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2951(.a(s_343), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2952(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2953(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2954(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate1247(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1248(.a(gate270inter0), .b(s_100), .O(gate270inter1));
  and2  gate1249(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1250(.a(s_100), .O(gate270inter3));
  inv1  gate1251(.a(s_101), .O(gate270inter4));
  nand2 gate1252(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1253(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1254(.a(G657), .O(gate270inter7));
  inv1  gate1255(.a(G785), .O(gate270inter8));
  nand2 gate1256(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1257(.a(s_101), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1258(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1259(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1260(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2255(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2256(.a(gate272inter0), .b(s_244), .O(gate272inter1));
  and2  gate2257(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2258(.a(s_244), .O(gate272inter3));
  inv1  gate2259(.a(s_245), .O(gate272inter4));
  nand2 gate2260(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2261(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2262(.a(G663), .O(gate272inter7));
  inv1  gate2263(.a(G791), .O(gate272inter8));
  nand2 gate2264(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2265(.a(s_245), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2266(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2267(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2268(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1191(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1192(.a(gate273inter0), .b(s_92), .O(gate273inter1));
  and2  gate1193(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1194(.a(s_92), .O(gate273inter3));
  inv1  gate1195(.a(s_93), .O(gate273inter4));
  nand2 gate1196(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1197(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1198(.a(G642), .O(gate273inter7));
  inv1  gate1199(.a(G794), .O(gate273inter8));
  nand2 gate1200(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1201(.a(s_93), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1202(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1203(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1204(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate701(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate702(.a(gate275inter0), .b(s_22), .O(gate275inter1));
  and2  gate703(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate704(.a(s_22), .O(gate275inter3));
  inv1  gate705(.a(s_23), .O(gate275inter4));
  nand2 gate706(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate707(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate708(.a(G645), .O(gate275inter7));
  inv1  gate709(.a(G797), .O(gate275inter8));
  nand2 gate710(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate711(.a(s_23), .b(gate275inter3), .O(gate275inter10));
  nor2  gate712(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate713(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate714(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2241(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2242(.a(gate279inter0), .b(s_242), .O(gate279inter1));
  and2  gate2243(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2244(.a(s_242), .O(gate279inter3));
  inv1  gate2245(.a(s_243), .O(gate279inter4));
  nand2 gate2246(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2247(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2248(.a(G651), .O(gate279inter7));
  inv1  gate2249(.a(G803), .O(gate279inter8));
  nand2 gate2250(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2251(.a(s_243), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2252(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2253(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2254(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2227(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2228(.a(gate283inter0), .b(s_240), .O(gate283inter1));
  and2  gate2229(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2230(.a(s_240), .O(gate283inter3));
  inv1  gate2231(.a(s_241), .O(gate283inter4));
  nand2 gate2232(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2233(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2234(.a(G657), .O(gate283inter7));
  inv1  gate2235(.a(G809), .O(gate283inter8));
  nand2 gate2236(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2237(.a(s_241), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2238(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2239(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2240(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2059(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2060(.a(gate285inter0), .b(s_216), .O(gate285inter1));
  and2  gate2061(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2062(.a(s_216), .O(gate285inter3));
  inv1  gate2063(.a(s_217), .O(gate285inter4));
  nand2 gate2064(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2065(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2066(.a(G660), .O(gate285inter7));
  inv1  gate2067(.a(G812), .O(gate285inter8));
  nand2 gate2068(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2069(.a(s_217), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2070(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2071(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2072(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1205(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1206(.a(gate286inter0), .b(s_94), .O(gate286inter1));
  and2  gate1207(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1208(.a(s_94), .O(gate286inter3));
  inv1  gate1209(.a(s_95), .O(gate286inter4));
  nand2 gate1210(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1211(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1212(.a(G788), .O(gate286inter7));
  inv1  gate1213(.a(G812), .O(gate286inter8));
  nand2 gate1214(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1215(.a(s_95), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1216(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1217(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1218(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate631(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate632(.a(gate287inter0), .b(s_12), .O(gate287inter1));
  and2  gate633(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate634(.a(s_12), .O(gate287inter3));
  inv1  gate635(.a(s_13), .O(gate287inter4));
  nand2 gate636(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate637(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate638(.a(G663), .O(gate287inter7));
  inv1  gate639(.a(G815), .O(gate287inter8));
  nand2 gate640(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate641(.a(s_13), .b(gate287inter3), .O(gate287inter10));
  nor2  gate642(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate643(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate644(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate687(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate688(.a(gate292inter0), .b(s_20), .O(gate292inter1));
  and2  gate689(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate690(.a(s_20), .O(gate292inter3));
  inv1  gate691(.a(s_21), .O(gate292inter4));
  nand2 gate692(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate693(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate694(.a(G824), .O(gate292inter7));
  inv1  gate695(.a(G825), .O(gate292inter8));
  nand2 gate696(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate697(.a(s_21), .b(gate292inter3), .O(gate292inter10));
  nor2  gate698(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate699(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate700(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2213(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2214(.a(gate294inter0), .b(s_238), .O(gate294inter1));
  and2  gate2215(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2216(.a(s_238), .O(gate294inter3));
  inv1  gate2217(.a(s_239), .O(gate294inter4));
  nand2 gate2218(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2219(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2220(.a(G832), .O(gate294inter7));
  inv1  gate2221(.a(G833), .O(gate294inter8));
  nand2 gate2222(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2223(.a(s_239), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2224(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2225(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2226(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate575(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate576(.a(gate295inter0), .b(s_4), .O(gate295inter1));
  and2  gate577(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate578(.a(s_4), .O(gate295inter3));
  inv1  gate579(.a(s_5), .O(gate295inter4));
  nand2 gate580(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate581(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate582(.a(G830), .O(gate295inter7));
  inv1  gate583(.a(G831), .O(gate295inter8));
  nand2 gate584(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate585(.a(s_5), .b(gate295inter3), .O(gate295inter10));
  nor2  gate586(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate587(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate588(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate3137(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate3138(.a(gate296inter0), .b(s_370), .O(gate296inter1));
  and2  gate3139(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate3140(.a(s_370), .O(gate296inter3));
  inv1  gate3141(.a(s_371), .O(gate296inter4));
  nand2 gate3142(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate3143(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate3144(.a(G826), .O(gate296inter7));
  inv1  gate3145(.a(G827), .O(gate296inter8));
  nand2 gate3146(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate3147(.a(s_371), .b(gate296inter3), .O(gate296inter10));
  nor2  gate3148(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate3149(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate3150(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1611(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1612(.a(gate387inter0), .b(s_152), .O(gate387inter1));
  and2  gate1613(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1614(.a(s_152), .O(gate387inter3));
  inv1  gate1615(.a(s_153), .O(gate387inter4));
  nand2 gate1616(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1617(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1618(.a(G1), .O(gate387inter7));
  inv1  gate1619(.a(G1036), .O(gate387inter8));
  nand2 gate1620(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1621(.a(s_153), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1622(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1623(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1624(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1037(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1038(.a(gate389inter0), .b(s_70), .O(gate389inter1));
  and2  gate1039(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1040(.a(s_70), .O(gate389inter3));
  inv1  gate1041(.a(s_71), .O(gate389inter4));
  nand2 gate1042(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1043(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1044(.a(G3), .O(gate389inter7));
  inv1  gate1045(.a(G1042), .O(gate389inter8));
  nand2 gate1046(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1047(.a(s_71), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1048(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1049(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1050(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate715(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate716(.a(gate390inter0), .b(s_24), .O(gate390inter1));
  and2  gate717(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate718(.a(s_24), .O(gate390inter3));
  inv1  gate719(.a(s_25), .O(gate390inter4));
  nand2 gate720(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate721(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate722(.a(G4), .O(gate390inter7));
  inv1  gate723(.a(G1045), .O(gate390inter8));
  nand2 gate724(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate725(.a(s_25), .b(gate390inter3), .O(gate390inter10));
  nor2  gate726(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate727(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate728(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate2605(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2606(.a(gate391inter0), .b(s_294), .O(gate391inter1));
  and2  gate2607(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2608(.a(s_294), .O(gate391inter3));
  inv1  gate2609(.a(s_295), .O(gate391inter4));
  nand2 gate2610(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2611(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2612(.a(G5), .O(gate391inter7));
  inv1  gate2613(.a(G1048), .O(gate391inter8));
  nand2 gate2614(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2615(.a(s_295), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2616(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2617(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2618(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1457(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1458(.a(gate393inter0), .b(s_130), .O(gate393inter1));
  and2  gate1459(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1460(.a(s_130), .O(gate393inter3));
  inv1  gate1461(.a(s_131), .O(gate393inter4));
  nand2 gate1462(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1463(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1464(.a(G7), .O(gate393inter7));
  inv1  gate1465(.a(G1054), .O(gate393inter8));
  nand2 gate1466(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1467(.a(s_131), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1468(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1469(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1470(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2633(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2634(.a(gate394inter0), .b(s_298), .O(gate394inter1));
  and2  gate2635(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2636(.a(s_298), .O(gate394inter3));
  inv1  gate2637(.a(s_299), .O(gate394inter4));
  nand2 gate2638(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2639(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2640(.a(G8), .O(gate394inter7));
  inv1  gate2641(.a(G1057), .O(gate394inter8));
  nand2 gate2642(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2643(.a(s_299), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2644(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2645(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2646(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1625(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1626(.a(gate396inter0), .b(s_154), .O(gate396inter1));
  and2  gate1627(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1628(.a(s_154), .O(gate396inter3));
  inv1  gate1629(.a(s_155), .O(gate396inter4));
  nand2 gate1630(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1631(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1632(.a(G10), .O(gate396inter7));
  inv1  gate1633(.a(G1063), .O(gate396inter8));
  nand2 gate1634(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1635(.a(s_155), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1636(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1637(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1638(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1751(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1752(.a(gate400inter0), .b(s_172), .O(gate400inter1));
  and2  gate1753(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1754(.a(s_172), .O(gate400inter3));
  inv1  gate1755(.a(s_173), .O(gate400inter4));
  nand2 gate1756(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1757(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1758(.a(G14), .O(gate400inter7));
  inv1  gate1759(.a(G1075), .O(gate400inter8));
  nand2 gate1760(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1761(.a(s_173), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1762(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1763(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1764(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2409(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2410(.a(gate402inter0), .b(s_266), .O(gate402inter1));
  and2  gate2411(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2412(.a(s_266), .O(gate402inter3));
  inv1  gate2413(.a(s_267), .O(gate402inter4));
  nand2 gate2414(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2415(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2416(.a(G16), .O(gate402inter7));
  inv1  gate2417(.a(G1081), .O(gate402inter8));
  nand2 gate2418(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2419(.a(s_267), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2420(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2421(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2422(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate2087(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2088(.a(gate403inter0), .b(s_220), .O(gate403inter1));
  and2  gate2089(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2090(.a(s_220), .O(gate403inter3));
  inv1  gate2091(.a(s_221), .O(gate403inter4));
  nand2 gate2092(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2093(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2094(.a(G17), .O(gate403inter7));
  inv1  gate2095(.a(G1084), .O(gate403inter8));
  nand2 gate2096(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2097(.a(s_221), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2098(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2099(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2100(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1989(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1990(.a(gate404inter0), .b(s_206), .O(gate404inter1));
  and2  gate1991(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1992(.a(s_206), .O(gate404inter3));
  inv1  gate1993(.a(s_207), .O(gate404inter4));
  nand2 gate1994(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1995(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1996(.a(G18), .O(gate404inter7));
  inv1  gate1997(.a(G1087), .O(gate404inter8));
  nand2 gate1998(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1999(.a(s_207), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2000(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2001(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2002(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2353(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2354(.a(gate409inter0), .b(s_258), .O(gate409inter1));
  and2  gate2355(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2356(.a(s_258), .O(gate409inter3));
  inv1  gate2357(.a(s_259), .O(gate409inter4));
  nand2 gate2358(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2359(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2360(.a(G23), .O(gate409inter7));
  inv1  gate2361(.a(G1102), .O(gate409inter8));
  nand2 gate2362(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2363(.a(s_259), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2364(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2365(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2366(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1345(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1346(.a(gate410inter0), .b(s_114), .O(gate410inter1));
  and2  gate1347(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1348(.a(s_114), .O(gate410inter3));
  inv1  gate1349(.a(s_115), .O(gate410inter4));
  nand2 gate1350(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1351(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1352(.a(G24), .O(gate410inter7));
  inv1  gate1353(.a(G1105), .O(gate410inter8));
  nand2 gate1354(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1355(.a(s_115), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1356(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1357(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1358(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate2745(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2746(.a(gate411inter0), .b(s_314), .O(gate411inter1));
  and2  gate2747(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2748(.a(s_314), .O(gate411inter3));
  inv1  gate2749(.a(s_315), .O(gate411inter4));
  nand2 gate2750(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2751(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2752(.a(G25), .O(gate411inter7));
  inv1  gate2753(.a(G1108), .O(gate411inter8));
  nand2 gate2754(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2755(.a(s_315), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2756(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2757(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2758(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1331(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1332(.a(gate412inter0), .b(s_112), .O(gate412inter1));
  and2  gate1333(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1334(.a(s_112), .O(gate412inter3));
  inv1  gate1335(.a(s_113), .O(gate412inter4));
  nand2 gate1336(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1337(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1338(.a(G26), .O(gate412inter7));
  inv1  gate1339(.a(G1111), .O(gate412inter8));
  nand2 gate1340(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1341(.a(s_113), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1342(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1343(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1344(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2857(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2858(.a(gate414inter0), .b(s_330), .O(gate414inter1));
  and2  gate2859(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2860(.a(s_330), .O(gate414inter3));
  inv1  gate2861(.a(s_331), .O(gate414inter4));
  nand2 gate2862(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2863(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2864(.a(G28), .O(gate414inter7));
  inv1  gate2865(.a(G1117), .O(gate414inter8));
  nand2 gate2866(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2867(.a(s_331), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2868(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2869(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2870(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2031(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2032(.a(gate416inter0), .b(s_212), .O(gate416inter1));
  and2  gate2033(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2034(.a(s_212), .O(gate416inter3));
  inv1  gate2035(.a(s_213), .O(gate416inter4));
  nand2 gate2036(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2037(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2038(.a(G30), .O(gate416inter7));
  inv1  gate2039(.a(G1123), .O(gate416inter8));
  nand2 gate2040(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2041(.a(s_213), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2042(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2043(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2044(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1933(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1934(.a(gate417inter0), .b(s_198), .O(gate417inter1));
  and2  gate1935(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1936(.a(s_198), .O(gate417inter3));
  inv1  gate1937(.a(s_199), .O(gate417inter4));
  nand2 gate1938(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1939(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1940(.a(G31), .O(gate417inter7));
  inv1  gate1941(.a(G1126), .O(gate417inter8));
  nand2 gate1942(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1943(.a(s_199), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1944(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1945(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1946(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate589(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate590(.a(gate418inter0), .b(s_6), .O(gate418inter1));
  and2  gate591(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate592(.a(s_6), .O(gate418inter3));
  inv1  gate593(.a(s_7), .O(gate418inter4));
  nand2 gate594(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate595(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate596(.a(G32), .O(gate418inter7));
  inv1  gate597(.a(G1129), .O(gate418inter8));
  nand2 gate598(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate599(.a(s_7), .b(gate418inter3), .O(gate418inter10));
  nor2  gate600(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate601(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate602(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2703(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2704(.a(gate420inter0), .b(s_308), .O(gate420inter1));
  and2  gate2705(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2706(.a(s_308), .O(gate420inter3));
  inv1  gate2707(.a(s_309), .O(gate420inter4));
  nand2 gate2708(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2709(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2710(.a(G1036), .O(gate420inter7));
  inv1  gate2711(.a(G1132), .O(gate420inter8));
  nand2 gate2712(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2713(.a(s_309), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2714(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2715(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2716(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2325(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2326(.a(gate421inter0), .b(s_254), .O(gate421inter1));
  and2  gate2327(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2328(.a(s_254), .O(gate421inter3));
  inv1  gate2329(.a(s_255), .O(gate421inter4));
  nand2 gate2330(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2331(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2332(.a(G2), .O(gate421inter7));
  inv1  gate2333(.a(G1135), .O(gate421inter8));
  nand2 gate2334(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2335(.a(s_255), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2336(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2337(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2338(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2661(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2662(.a(gate422inter0), .b(s_302), .O(gate422inter1));
  and2  gate2663(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2664(.a(s_302), .O(gate422inter3));
  inv1  gate2665(.a(s_303), .O(gate422inter4));
  nand2 gate2666(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2667(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2668(.a(G1039), .O(gate422inter7));
  inv1  gate2669(.a(G1135), .O(gate422inter8));
  nand2 gate2670(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2671(.a(s_303), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2672(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2673(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2674(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2003(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2004(.a(gate425inter0), .b(s_208), .O(gate425inter1));
  and2  gate2005(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2006(.a(s_208), .O(gate425inter3));
  inv1  gate2007(.a(s_209), .O(gate425inter4));
  nand2 gate2008(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2009(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2010(.a(G4), .O(gate425inter7));
  inv1  gate2011(.a(G1141), .O(gate425inter8));
  nand2 gate2012(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2013(.a(s_209), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2014(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2015(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2016(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate3207(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate3208(.a(gate426inter0), .b(s_380), .O(gate426inter1));
  and2  gate3209(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate3210(.a(s_380), .O(gate426inter3));
  inv1  gate3211(.a(s_381), .O(gate426inter4));
  nand2 gate3212(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate3213(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate3214(.a(G1045), .O(gate426inter7));
  inv1  gate3215(.a(G1141), .O(gate426inter8));
  nand2 gate3216(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate3217(.a(s_381), .b(gate426inter3), .O(gate426inter10));
  nor2  gate3218(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate3219(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate3220(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate561(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate562(.a(gate428inter0), .b(s_2), .O(gate428inter1));
  and2  gate563(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate564(.a(s_2), .O(gate428inter3));
  inv1  gate565(.a(s_3), .O(gate428inter4));
  nand2 gate566(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate567(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate568(.a(G1048), .O(gate428inter7));
  inv1  gate569(.a(G1144), .O(gate428inter8));
  nand2 gate570(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate571(.a(s_3), .b(gate428inter3), .O(gate428inter10));
  nor2  gate572(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate573(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate574(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate771(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate772(.a(gate430inter0), .b(s_32), .O(gate430inter1));
  and2  gate773(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate774(.a(s_32), .O(gate430inter3));
  inv1  gate775(.a(s_33), .O(gate430inter4));
  nand2 gate776(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate777(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate778(.a(G1051), .O(gate430inter7));
  inv1  gate779(.a(G1147), .O(gate430inter8));
  nand2 gate780(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate781(.a(s_33), .b(gate430inter3), .O(gate430inter10));
  nor2  gate782(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate783(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate784(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1401(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1402(.a(gate436inter0), .b(s_122), .O(gate436inter1));
  and2  gate1403(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1404(.a(s_122), .O(gate436inter3));
  inv1  gate1405(.a(s_123), .O(gate436inter4));
  nand2 gate1406(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1407(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1408(.a(G1060), .O(gate436inter7));
  inv1  gate1409(.a(G1156), .O(gate436inter8));
  nand2 gate1410(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1411(.a(s_123), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1412(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1413(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1414(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2507(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2508(.a(gate441inter0), .b(s_280), .O(gate441inter1));
  and2  gate2509(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2510(.a(s_280), .O(gate441inter3));
  inv1  gate2511(.a(s_281), .O(gate441inter4));
  nand2 gate2512(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2513(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2514(.a(G12), .O(gate441inter7));
  inv1  gate2515(.a(G1165), .O(gate441inter8));
  nand2 gate2516(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2517(.a(s_281), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2518(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2519(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2520(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1919(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1920(.a(gate443inter0), .b(s_196), .O(gate443inter1));
  and2  gate1921(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1922(.a(s_196), .O(gate443inter3));
  inv1  gate1923(.a(s_197), .O(gate443inter4));
  nand2 gate1924(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1925(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1926(.a(G13), .O(gate443inter7));
  inv1  gate1927(.a(G1168), .O(gate443inter8));
  nand2 gate1928(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1929(.a(s_197), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1930(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1931(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1932(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1079(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1080(.a(gate446inter0), .b(s_76), .O(gate446inter1));
  and2  gate1081(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1082(.a(s_76), .O(gate446inter3));
  inv1  gate1083(.a(s_77), .O(gate446inter4));
  nand2 gate1084(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1085(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1086(.a(G1075), .O(gate446inter7));
  inv1  gate1087(.a(G1171), .O(gate446inter8));
  nand2 gate1088(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1089(.a(s_77), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1090(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1091(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1092(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2899(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2900(.a(gate448inter0), .b(s_336), .O(gate448inter1));
  and2  gate2901(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2902(.a(s_336), .O(gate448inter3));
  inv1  gate2903(.a(s_337), .O(gate448inter4));
  nand2 gate2904(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2905(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2906(.a(G1078), .O(gate448inter7));
  inv1  gate2907(.a(G1174), .O(gate448inter8));
  nand2 gate2908(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2909(.a(s_337), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2910(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2911(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2912(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1219(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1220(.a(gate449inter0), .b(s_96), .O(gate449inter1));
  and2  gate1221(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1222(.a(s_96), .O(gate449inter3));
  inv1  gate1223(.a(s_97), .O(gate449inter4));
  nand2 gate1224(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1225(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1226(.a(G16), .O(gate449inter7));
  inv1  gate1227(.a(G1177), .O(gate449inter8));
  nand2 gate1228(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1229(.a(s_97), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1230(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1231(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1232(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1135(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1136(.a(gate454inter0), .b(s_84), .O(gate454inter1));
  and2  gate1137(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1138(.a(s_84), .O(gate454inter3));
  inv1  gate1139(.a(s_85), .O(gate454inter4));
  nand2 gate1140(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1141(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1142(.a(G1087), .O(gate454inter7));
  inv1  gate1143(.a(G1183), .O(gate454inter8));
  nand2 gate1144(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1145(.a(s_85), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1146(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1147(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1148(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2983(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2984(.a(gate457inter0), .b(s_348), .O(gate457inter1));
  and2  gate2985(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2986(.a(s_348), .O(gate457inter3));
  inv1  gate2987(.a(s_349), .O(gate457inter4));
  nand2 gate2988(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2989(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2990(.a(G20), .O(gate457inter7));
  inv1  gate2991(.a(G1189), .O(gate457inter8));
  nand2 gate2992(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2993(.a(s_349), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2994(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2995(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2996(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1163(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1164(.a(gate458inter0), .b(s_88), .O(gate458inter1));
  and2  gate1165(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1166(.a(s_88), .O(gate458inter3));
  inv1  gate1167(.a(s_89), .O(gate458inter4));
  nand2 gate1168(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1169(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1170(.a(G1093), .O(gate458inter7));
  inv1  gate1171(.a(G1189), .O(gate458inter8));
  nand2 gate1172(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1173(.a(s_89), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1174(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1175(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1176(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1639(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1640(.a(gate469inter0), .b(s_156), .O(gate469inter1));
  and2  gate1641(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1642(.a(s_156), .O(gate469inter3));
  inv1  gate1643(.a(s_157), .O(gate469inter4));
  nand2 gate1644(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1645(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1646(.a(G26), .O(gate469inter7));
  inv1  gate1647(.a(G1207), .O(gate469inter8));
  nand2 gate1648(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1649(.a(s_157), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1650(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1651(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1652(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2017(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2018(.a(gate470inter0), .b(s_210), .O(gate470inter1));
  and2  gate2019(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2020(.a(s_210), .O(gate470inter3));
  inv1  gate2021(.a(s_211), .O(gate470inter4));
  nand2 gate2022(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2023(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2024(.a(G1111), .O(gate470inter7));
  inv1  gate2025(.a(G1207), .O(gate470inter8));
  nand2 gate2026(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2027(.a(s_211), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2028(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2029(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2030(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2283(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2284(.a(gate471inter0), .b(s_248), .O(gate471inter1));
  and2  gate2285(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2286(.a(s_248), .O(gate471inter3));
  inv1  gate2287(.a(s_249), .O(gate471inter4));
  nand2 gate2288(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2289(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2290(.a(G27), .O(gate471inter7));
  inv1  gate2291(.a(G1210), .O(gate471inter8));
  nand2 gate2292(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2293(.a(s_249), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2294(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2295(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2296(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2493(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2494(.a(gate472inter0), .b(s_278), .O(gate472inter1));
  and2  gate2495(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2496(.a(s_278), .O(gate472inter3));
  inv1  gate2497(.a(s_279), .O(gate472inter4));
  nand2 gate2498(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2499(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2500(.a(G1114), .O(gate472inter7));
  inv1  gate2501(.a(G1210), .O(gate472inter8));
  nand2 gate2502(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2503(.a(s_279), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2504(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2505(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2506(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate995(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate996(.a(gate473inter0), .b(s_64), .O(gate473inter1));
  and2  gate997(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate998(.a(s_64), .O(gate473inter3));
  inv1  gate999(.a(s_65), .O(gate473inter4));
  nand2 gate1000(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1001(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1002(.a(G28), .O(gate473inter7));
  inv1  gate1003(.a(G1213), .O(gate473inter8));
  nand2 gate1004(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1005(.a(s_65), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1006(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1007(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1008(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate3193(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate3194(.a(gate474inter0), .b(s_378), .O(gate474inter1));
  and2  gate3195(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate3196(.a(s_378), .O(gate474inter3));
  inv1  gate3197(.a(s_379), .O(gate474inter4));
  nand2 gate3198(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate3199(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate3200(.a(G1117), .O(gate474inter7));
  inv1  gate3201(.a(G1213), .O(gate474inter8));
  nand2 gate3202(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate3203(.a(s_379), .b(gate474inter3), .O(gate474inter10));
  nor2  gate3204(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate3205(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate3206(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate785(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate786(.a(gate475inter0), .b(s_34), .O(gate475inter1));
  and2  gate787(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate788(.a(s_34), .O(gate475inter3));
  inv1  gate789(.a(s_35), .O(gate475inter4));
  nand2 gate790(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate791(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate792(.a(G29), .O(gate475inter7));
  inv1  gate793(.a(G1216), .O(gate475inter8));
  nand2 gate794(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate795(.a(s_35), .b(gate475inter3), .O(gate475inter10));
  nor2  gate796(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate797(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate798(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2997(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2998(.a(gate476inter0), .b(s_350), .O(gate476inter1));
  and2  gate2999(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate3000(.a(s_350), .O(gate476inter3));
  inv1  gate3001(.a(s_351), .O(gate476inter4));
  nand2 gate3002(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate3003(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate3004(.a(G1120), .O(gate476inter7));
  inv1  gate3005(.a(G1216), .O(gate476inter8));
  nand2 gate3006(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate3007(.a(s_351), .b(gate476inter3), .O(gate476inter10));
  nor2  gate3008(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate3009(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate3010(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1891(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1892(.a(gate477inter0), .b(s_192), .O(gate477inter1));
  and2  gate1893(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1894(.a(s_192), .O(gate477inter3));
  inv1  gate1895(.a(s_193), .O(gate477inter4));
  nand2 gate1896(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1897(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1898(.a(G30), .O(gate477inter7));
  inv1  gate1899(.a(G1219), .O(gate477inter8));
  nand2 gate1900(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1901(.a(s_193), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1902(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1903(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1904(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1009(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1010(.a(gate481inter0), .b(s_66), .O(gate481inter1));
  and2  gate1011(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1012(.a(s_66), .O(gate481inter3));
  inv1  gate1013(.a(s_67), .O(gate481inter4));
  nand2 gate1014(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1015(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1016(.a(G32), .O(gate481inter7));
  inv1  gate1017(.a(G1225), .O(gate481inter8));
  nand2 gate1018(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1019(.a(s_67), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1020(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1021(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1022(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2101(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2102(.a(gate483inter0), .b(s_222), .O(gate483inter1));
  and2  gate2103(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2104(.a(s_222), .O(gate483inter3));
  inv1  gate2105(.a(s_223), .O(gate483inter4));
  nand2 gate2106(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2107(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2108(.a(G1228), .O(gate483inter7));
  inv1  gate2109(.a(G1229), .O(gate483inter8));
  nand2 gate2110(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2111(.a(s_223), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2112(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2113(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2114(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate3291(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate3292(.a(gate487inter0), .b(s_392), .O(gate487inter1));
  and2  gate3293(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate3294(.a(s_392), .O(gate487inter3));
  inv1  gate3295(.a(s_393), .O(gate487inter4));
  nand2 gate3296(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate3297(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate3298(.a(G1236), .O(gate487inter7));
  inv1  gate3299(.a(G1237), .O(gate487inter8));
  nand2 gate3300(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate3301(.a(s_393), .b(gate487inter3), .O(gate487inter10));
  nor2  gate3302(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate3303(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate3304(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1723(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1724(.a(gate489inter0), .b(s_168), .O(gate489inter1));
  and2  gate1725(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1726(.a(s_168), .O(gate489inter3));
  inv1  gate1727(.a(s_169), .O(gate489inter4));
  nand2 gate1728(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1729(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1730(.a(G1240), .O(gate489inter7));
  inv1  gate1731(.a(G1241), .O(gate489inter8));
  nand2 gate1732(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1733(.a(s_169), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1734(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1735(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1736(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1807(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1808(.a(gate490inter0), .b(s_180), .O(gate490inter1));
  and2  gate1809(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1810(.a(s_180), .O(gate490inter3));
  inv1  gate1811(.a(s_181), .O(gate490inter4));
  nand2 gate1812(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1813(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1814(.a(G1242), .O(gate490inter7));
  inv1  gate1815(.a(G1243), .O(gate490inter8));
  nand2 gate1816(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1817(.a(s_181), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1818(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1819(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1820(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1821(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1822(.a(gate492inter0), .b(s_182), .O(gate492inter1));
  and2  gate1823(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1824(.a(s_182), .O(gate492inter3));
  inv1  gate1825(.a(s_183), .O(gate492inter4));
  nand2 gate1826(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1827(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1828(.a(G1246), .O(gate492inter7));
  inv1  gate1829(.a(G1247), .O(gate492inter8));
  nand2 gate1830(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1831(.a(s_183), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1832(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1833(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1834(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1527(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1528(.a(gate495inter0), .b(s_140), .O(gate495inter1));
  and2  gate1529(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1530(.a(s_140), .O(gate495inter3));
  inv1  gate1531(.a(s_141), .O(gate495inter4));
  nand2 gate1532(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1533(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1534(.a(G1252), .O(gate495inter7));
  inv1  gate1535(.a(G1253), .O(gate495inter8));
  nand2 gate1536(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1537(.a(s_141), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1538(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1539(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1540(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate841(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate842(.a(gate500inter0), .b(s_42), .O(gate500inter1));
  and2  gate843(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate844(.a(s_42), .O(gate500inter3));
  inv1  gate845(.a(s_43), .O(gate500inter4));
  nand2 gate846(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate847(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate848(.a(G1262), .O(gate500inter7));
  inv1  gate849(.a(G1263), .O(gate500inter8));
  nand2 gate850(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate851(.a(s_43), .b(gate500inter3), .O(gate500inter10));
  nor2  gate852(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate853(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate854(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2647(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2648(.a(gate501inter0), .b(s_300), .O(gate501inter1));
  and2  gate2649(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2650(.a(s_300), .O(gate501inter3));
  inv1  gate2651(.a(s_301), .O(gate501inter4));
  nand2 gate2652(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2653(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2654(.a(G1264), .O(gate501inter7));
  inv1  gate2655(.a(G1265), .O(gate501inter8));
  nand2 gate2656(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2657(.a(s_301), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2658(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2659(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2660(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1835(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1836(.a(gate502inter0), .b(s_184), .O(gate502inter1));
  and2  gate1837(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1838(.a(s_184), .O(gate502inter3));
  inv1  gate1839(.a(s_185), .O(gate502inter4));
  nand2 gate1840(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1841(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1842(.a(G1266), .O(gate502inter7));
  inv1  gate1843(.a(G1267), .O(gate502inter8));
  nand2 gate1844(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1845(.a(s_185), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1846(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1847(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1848(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate2185(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2186(.a(gate504inter0), .b(s_234), .O(gate504inter1));
  and2  gate2187(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2188(.a(s_234), .O(gate504inter3));
  inv1  gate2189(.a(s_235), .O(gate504inter4));
  nand2 gate2190(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2191(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2192(.a(G1270), .O(gate504inter7));
  inv1  gate2193(.a(G1271), .O(gate504inter8));
  nand2 gate2194(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2195(.a(s_235), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2196(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2197(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2198(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2269(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2270(.a(gate507inter0), .b(s_246), .O(gate507inter1));
  and2  gate2271(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2272(.a(s_246), .O(gate507inter3));
  inv1  gate2273(.a(s_247), .O(gate507inter4));
  nand2 gate2274(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2275(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2276(.a(G1276), .O(gate507inter7));
  inv1  gate2277(.a(G1277), .O(gate507inter8));
  nand2 gate2278(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2279(.a(s_247), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2280(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2281(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2282(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2689(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2690(.a(gate508inter0), .b(s_306), .O(gate508inter1));
  and2  gate2691(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2692(.a(s_306), .O(gate508inter3));
  inv1  gate2693(.a(s_307), .O(gate508inter4));
  nand2 gate2694(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2695(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2696(.a(G1278), .O(gate508inter7));
  inv1  gate2697(.a(G1279), .O(gate508inter8));
  nand2 gate2698(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2699(.a(s_307), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2700(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2701(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2702(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2675(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2676(.a(gate510inter0), .b(s_304), .O(gate510inter1));
  and2  gate2677(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2678(.a(s_304), .O(gate510inter3));
  inv1  gate2679(.a(s_305), .O(gate510inter4));
  nand2 gate2680(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2681(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2682(.a(G1282), .O(gate510inter7));
  inv1  gate2683(.a(G1283), .O(gate510inter8));
  nand2 gate2684(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2685(.a(s_305), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2686(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2687(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2688(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate897(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate898(.a(gate513inter0), .b(s_50), .O(gate513inter1));
  and2  gate899(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate900(.a(s_50), .O(gate513inter3));
  inv1  gate901(.a(s_51), .O(gate513inter4));
  nand2 gate902(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate903(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate904(.a(G1288), .O(gate513inter7));
  inv1  gate905(.a(G1289), .O(gate513inter8));
  nand2 gate906(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate907(.a(s_51), .b(gate513inter3), .O(gate513inter10));
  nor2  gate908(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate909(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate910(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1681(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1682(.a(gate514inter0), .b(s_162), .O(gate514inter1));
  and2  gate1683(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1684(.a(s_162), .O(gate514inter3));
  inv1  gate1685(.a(s_163), .O(gate514inter4));
  nand2 gate1686(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1687(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1688(.a(G1290), .O(gate514inter7));
  inv1  gate1689(.a(G1291), .O(gate514inter8));
  nand2 gate1690(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1691(.a(s_163), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1692(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1693(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1694(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule