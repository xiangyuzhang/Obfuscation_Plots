module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2297(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2298(.a(gate10inter0), .b(s_250), .O(gate10inter1));
  and2  gate2299(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2300(.a(s_250), .O(gate10inter3));
  inv1  gate2301(.a(s_251), .O(gate10inter4));
  nand2 gate2302(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2303(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2304(.a(G3), .O(gate10inter7));
  inv1  gate2305(.a(G4), .O(gate10inter8));
  nand2 gate2306(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2307(.a(s_251), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2308(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2309(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2310(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate1443(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1444(.a(gate11inter0), .b(s_128), .O(gate11inter1));
  and2  gate1445(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1446(.a(s_128), .O(gate11inter3));
  inv1  gate1447(.a(s_129), .O(gate11inter4));
  nand2 gate1448(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1449(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1450(.a(G5), .O(gate11inter7));
  inv1  gate1451(.a(G6), .O(gate11inter8));
  nand2 gate1452(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1453(.a(s_129), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1454(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1455(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1456(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1051(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1052(.a(gate14inter0), .b(s_72), .O(gate14inter1));
  and2  gate1053(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1054(.a(s_72), .O(gate14inter3));
  inv1  gate1055(.a(s_73), .O(gate14inter4));
  nand2 gate1056(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1057(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1058(.a(G11), .O(gate14inter7));
  inv1  gate1059(.a(G12), .O(gate14inter8));
  nand2 gate1060(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1061(.a(s_73), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1062(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1063(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1064(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1023(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1024(.a(gate15inter0), .b(s_68), .O(gate15inter1));
  and2  gate1025(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1026(.a(s_68), .O(gate15inter3));
  inv1  gate1027(.a(s_69), .O(gate15inter4));
  nand2 gate1028(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1029(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1030(.a(G13), .O(gate15inter7));
  inv1  gate1031(.a(G14), .O(gate15inter8));
  nand2 gate1032(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1033(.a(s_69), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1034(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1035(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1036(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate939(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate940(.a(gate16inter0), .b(s_56), .O(gate16inter1));
  and2  gate941(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate942(.a(s_56), .O(gate16inter3));
  inv1  gate943(.a(s_57), .O(gate16inter4));
  nand2 gate944(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate945(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate946(.a(G15), .O(gate16inter7));
  inv1  gate947(.a(G16), .O(gate16inter8));
  nand2 gate948(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate949(.a(s_57), .b(gate16inter3), .O(gate16inter10));
  nor2  gate950(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate951(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate952(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2493(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2494(.a(gate18inter0), .b(s_278), .O(gate18inter1));
  and2  gate2495(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2496(.a(s_278), .O(gate18inter3));
  inv1  gate2497(.a(s_279), .O(gate18inter4));
  nand2 gate2498(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2499(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2500(.a(G19), .O(gate18inter7));
  inv1  gate2501(.a(G20), .O(gate18inter8));
  nand2 gate2502(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2503(.a(s_279), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2504(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2505(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2506(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2213(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2214(.a(gate20inter0), .b(s_238), .O(gate20inter1));
  and2  gate2215(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2216(.a(s_238), .O(gate20inter3));
  inv1  gate2217(.a(s_239), .O(gate20inter4));
  nand2 gate2218(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2219(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2220(.a(G23), .O(gate20inter7));
  inv1  gate2221(.a(G24), .O(gate20inter8));
  nand2 gate2222(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2223(.a(s_239), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2224(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2225(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2226(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1723(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1724(.a(gate22inter0), .b(s_168), .O(gate22inter1));
  and2  gate1725(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1726(.a(s_168), .O(gate22inter3));
  inv1  gate1727(.a(s_169), .O(gate22inter4));
  nand2 gate1728(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1729(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1730(.a(G27), .O(gate22inter7));
  inv1  gate1731(.a(G28), .O(gate22inter8));
  nand2 gate1732(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1733(.a(s_169), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1734(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1735(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1736(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1639(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1640(.a(gate23inter0), .b(s_156), .O(gate23inter1));
  and2  gate1641(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1642(.a(s_156), .O(gate23inter3));
  inv1  gate1643(.a(s_157), .O(gate23inter4));
  nand2 gate1644(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1645(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1646(.a(G29), .O(gate23inter7));
  inv1  gate1647(.a(G30), .O(gate23inter8));
  nand2 gate1648(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1649(.a(s_157), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1650(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1651(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1652(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1891(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1892(.a(gate26inter0), .b(s_192), .O(gate26inter1));
  and2  gate1893(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1894(.a(s_192), .O(gate26inter3));
  inv1  gate1895(.a(s_193), .O(gate26inter4));
  nand2 gate1896(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1897(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1898(.a(G9), .O(gate26inter7));
  inv1  gate1899(.a(G13), .O(gate26inter8));
  nand2 gate1900(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1901(.a(s_193), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1902(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1903(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1904(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1807(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1808(.a(gate29inter0), .b(s_180), .O(gate29inter1));
  and2  gate1809(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1810(.a(s_180), .O(gate29inter3));
  inv1  gate1811(.a(s_181), .O(gate29inter4));
  nand2 gate1812(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1813(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1814(.a(G3), .O(gate29inter7));
  inv1  gate1815(.a(G7), .O(gate29inter8));
  nand2 gate1816(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1817(.a(s_181), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1818(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1819(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1820(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1989(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1990(.a(gate34inter0), .b(s_206), .O(gate34inter1));
  and2  gate1991(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1992(.a(s_206), .O(gate34inter3));
  inv1  gate1993(.a(s_207), .O(gate34inter4));
  nand2 gate1994(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1995(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1996(.a(G25), .O(gate34inter7));
  inv1  gate1997(.a(G29), .O(gate34inter8));
  nand2 gate1998(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1999(.a(s_207), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2000(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2001(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2002(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate2157(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2158(.a(gate35inter0), .b(s_230), .O(gate35inter1));
  and2  gate2159(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2160(.a(s_230), .O(gate35inter3));
  inv1  gate2161(.a(s_231), .O(gate35inter4));
  nand2 gate2162(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2163(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2164(.a(G18), .O(gate35inter7));
  inv1  gate2165(.a(G22), .O(gate35inter8));
  nand2 gate2166(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2167(.a(s_231), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2168(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2169(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2170(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2241(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2242(.a(gate36inter0), .b(s_242), .O(gate36inter1));
  and2  gate2243(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2244(.a(s_242), .O(gate36inter3));
  inv1  gate2245(.a(s_243), .O(gate36inter4));
  nand2 gate2246(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2247(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2248(.a(G26), .O(gate36inter7));
  inv1  gate2249(.a(G30), .O(gate36inter8));
  nand2 gate2250(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2251(.a(s_243), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2252(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2253(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2254(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate855(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate856(.a(gate37inter0), .b(s_44), .O(gate37inter1));
  and2  gate857(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate858(.a(s_44), .O(gate37inter3));
  inv1  gate859(.a(s_45), .O(gate37inter4));
  nand2 gate860(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate861(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate862(.a(G19), .O(gate37inter7));
  inv1  gate863(.a(G23), .O(gate37inter8));
  nand2 gate864(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate865(.a(s_45), .b(gate37inter3), .O(gate37inter10));
  nor2  gate866(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate867(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate868(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1947(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1948(.a(gate38inter0), .b(s_200), .O(gate38inter1));
  and2  gate1949(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1950(.a(s_200), .O(gate38inter3));
  inv1  gate1951(.a(s_201), .O(gate38inter4));
  nand2 gate1952(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1953(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1954(.a(G27), .O(gate38inter7));
  inv1  gate1955(.a(G31), .O(gate38inter8));
  nand2 gate1956(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1957(.a(s_201), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1958(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1959(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1960(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2255(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2256(.a(gate40inter0), .b(s_244), .O(gate40inter1));
  and2  gate2257(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2258(.a(s_244), .O(gate40inter3));
  inv1  gate2259(.a(s_245), .O(gate40inter4));
  nand2 gate2260(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2261(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2262(.a(G28), .O(gate40inter7));
  inv1  gate2263(.a(G32), .O(gate40inter8));
  nand2 gate2264(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2265(.a(s_245), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2266(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2267(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2268(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate659(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate660(.a(gate45inter0), .b(s_16), .O(gate45inter1));
  and2  gate661(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate662(.a(s_16), .O(gate45inter3));
  inv1  gate663(.a(s_17), .O(gate45inter4));
  nand2 gate664(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate665(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate666(.a(G5), .O(gate45inter7));
  inv1  gate667(.a(G272), .O(gate45inter8));
  nand2 gate668(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate669(.a(s_17), .b(gate45inter3), .O(gate45inter10));
  nor2  gate670(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate671(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate672(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate701(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate702(.a(gate46inter0), .b(s_22), .O(gate46inter1));
  and2  gate703(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate704(.a(s_22), .O(gate46inter3));
  inv1  gate705(.a(s_23), .O(gate46inter4));
  nand2 gate706(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate707(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate708(.a(G6), .O(gate46inter7));
  inv1  gate709(.a(G272), .O(gate46inter8));
  nand2 gate710(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate711(.a(s_23), .b(gate46inter3), .O(gate46inter10));
  nor2  gate712(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate713(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate714(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1709(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1710(.a(gate47inter0), .b(s_166), .O(gate47inter1));
  and2  gate1711(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1712(.a(s_166), .O(gate47inter3));
  inv1  gate1713(.a(s_167), .O(gate47inter4));
  nand2 gate1714(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1715(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1716(.a(G7), .O(gate47inter7));
  inv1  gate1717(.a(G275), .O(gate47inter8));
  nand2 gate1718(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1719(.a(s_167), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1720(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1721(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1722(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2101(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2102(.a(gate51inter0), .b(s_222), .O(gate51inter1));
  and2  gate2103(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2104(.a(s_222), .O(gate51inter3));
  inv1  gate2105(.a(s_223), .O(gate51inter4));
  nand2 gate2106(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2107(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2108(.a(G11), .O(gate51inter7));
  inv1  gate2109(.a(G281), .O(gate51inter8));
  nand2 gate2110(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2111(.a(s_223), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2112(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2113(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2114(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate2381(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2382(.a(gate52inter0), .b(s_262), .O(gate52inter1));
  and2  gate2383(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2384(.a(s_262), .O(gate52inter3));
  inv1  gate2385(.a(s_263), .O(gate52inter4));
  nand2 gate2386(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2387(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2388(.a(G12), .O(gate52inter7));
  inv1  gate2389(.a(G281), .O(gate52inter8));
  nand2 gate2390(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2391(.a(s_263), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2392(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2393(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2394(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1779(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1780(.a(gate57inter0), .b(s_176), .O(gate57inter1));
  and2  gate1781(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1782(.a(s_176), .O(gate57inter3));
  inv1  gate1783(.a(s_177), .O(gate57inter4));
  nand2 gate1784(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1785(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1786(.a(G17), .O(gate57inter7));
  inv1  gate1787(.a(G290), .O(gate57inter8));
  nand2 gate1788(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1789(.a(s_177), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1790(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1791(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1792(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate715(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate716(.a(gate64inter0), .b(s_24), .O(gate64inter1));
  and2  gate717(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate718(.a(s_24), .O(gate64inter3));
  inv1  gate719(.a(s_25), .O(gate64inter4));
  nand2 gate720(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate721(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate722(.a(G24), .O(gate64inter7));
  inv1  gate723(.a(G299), .O(gate64inter8));
  nand2 gate724(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate725(.a(s_25), .b(gate64inter3), .O(gate64inter10));
  nor2  gate726(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate727(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate728(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate561(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate562(.a(gate65inter0), .b(s_2), .O(gate65inter1));
  and2  gate563(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate564(.a(s_2), .O(gate65inter3));
  inv1  gate565(.a(s_3), .O(gate65inter4));
  nand2 gate566(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate567(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate568(.a(G25), .O(gate65inter7));
  inv1  gate569(.a(G302), .O(gate65inter8));
  nand2 gate570(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate571(.a(s_3), .b(gate65inter3), .O(gate65inter10));
  nor2  gate572(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate573(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate574(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1205(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1206(.a(gate66inter0), .b(s_94), .O(gate66inter1));
  and2  gate1207(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1208(.a(s_94), .O(gate66inter3));
  inv1  gate1209(.a(s_95), .O(gate66inter4));
  nand2 gate1210(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1211(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1212(.a(G26), .O(gate66inter7));
  inv1  gate1213(.a(G302), .O(gate66inter8));
  nand2 gate1214(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1215(.a(s_95), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1216(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1217(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1218(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate603(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate604(.a(gate69inter0), .b(s_8), .O(gate69inter1));
  and2  gate605(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate606(.a(s_8), .O(gate69inter3));
  inv1  gate607(.a(s_9), .O(gate69inter4));
  nand2 gate608(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate609(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate610(.a(G29), .O(gate69inter7));
  inv1  gate611(.a(G308), .O(gate69inter8));
  nand2 gate612(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate613(.a(s_9), .b(gate69inter3), .O(gate69inter10));
  nor2  gate614(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate615(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate616(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2017(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2018(.a(gate71inter0), .b(s_210), .O(gate71inter1));
  and2  gate2019(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2020(.a(s_210), .O(gate71inter3));
  inv1  gate2021(.a(s_211), .O(gate71inter4));
  nand2 gate2022(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2023(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2024(.a(G31), .O(gate71inter7));
  inv1  gate2025(.a(G311), .O(gate71inter8));
  nand2 gate2026(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2027(.a(s_211), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2028(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2029(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2030(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate841(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate842(.a(gate73inter0), .b(s_42), .O(gate73inter1));
  and2  gate843(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate844(.a(s_42), .O(gate73inter3));
  inv1  gate845(.a(s_43), .O(gate73inter4));
  nand2 gate846(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate847(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate848(.a(G1), .O(gate73inter7));
  inv1  gate849(.a(G314), .O(gate73inter8));
  nand2 gate850(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate851(.a(s_43), .b(gate73inter3), .O(gate73inter10));
  nor2  gate852(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate853(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate854(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2199(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2200(.a(gate74inter0), .b(s_236), .O(gate74inter1));
  and2  gate2201(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2202(.a(s_236), .O(gate74inter3));
  inv1  gate2203(.a(s_237), .O(gate74inter4));
  nand2 gate2204(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2205(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2206(.a(G5), .O(gate74inter7));
  inv1  gate2207(.a(G314), .O(gate74inter8));
  nand2 gate2208(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2209(.a(s_237), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2210(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2211(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2212(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1135(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1136(.a(gate76inter0), .b(s_84), .O(gate76inter1));
  and2  gate1137(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1138(.a(s_84), .O(gate76inter3));
  inv1  gate1139(.a(s_85), .O(gate76inter4));
  nand2 gate1140(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1141(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1142(.a(G13), .O(gate76inter7));
  inv1  gate1143(.a(G317), .O(gate76inter8));
  nand2 gate1144(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1145(.a(s_85), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1146(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1147(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1148(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate2227(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2228(.a(gate77inter0), .b(s_240), .O(gate77inter1));
  and2  gate2229(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2230(.a(s_240), .O(gate77inter3));
  inv1  gate2231(.a(s_241), .O(gate77inter4));
  nand2 gate2232(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2233(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2234(.a(G2), .O(gate77inter7));
  inv1  gate2235(.a(G320), .O(gate77inter8));
  nand2 gate2236(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2237(.a(s_241), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2238(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2239(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2240(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1247(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1248(.a(gate78inter0), .b(s_100), .O(gate78inter1));
  and2  gate1249(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1250(.a(s_100), .O(gate78inter3));
  inv1  gate1251(.a(s_101), .O(gate78inter4));
  nand2 gate1252(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1253(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1254(.a(G6), .O(gate78inter7));
  inv1  gate1255(.a(G320), .O(gate78inter8));
  nand2 gate1256(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1257(.a(s_101), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1258(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1259(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1260(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1961(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1962(.a(gate80inter0), .b(s_202), .O(gate80inter1));
  and2  gate1963(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1964(.a(s_202), .O(gate80inter3));
  inv1  gate1965(.a(s_203), .O(gate80inter4));
  nand2 gate1966(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1967(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1968(.a(G14), .O(gate80inter7));
  inv1  gate1969(.a(G323), .O(gate80inter8));
  nand2 gate1970(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1971(.a(s_203), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1972(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1973(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1974(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate869(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate870(.a(gate81inter0), .b(s_46), .O(gate81inter1));
  and2  gate871(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate872(.a(s_46), .O(gate81inter3));
  inv1  gate873(.a(s_47), .O(gate81inter4));
  nand2 gate874(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate875(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate876(.a(G3), .O(gate81inter7));
  inv1  gate877(.a(G326), .O(gate81inter8));
  nand2 gate878(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate879(.a(s_47), .b(gate81inter3), .O(gate81inter10));
  nor2  gate880(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate881(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate882(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate883(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate884(.a(gate82inter0), .b(s_48), .O(gate82inter1));
  and2  gate885(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate886(.a(s_48), .O(gate82inter3));
  inv1  gate887(.a(s_49), .O(gate82inter4));
  nand2 gate888(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate889(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate890(.a(G7), .O(gate82inter7));
  inv1  gate891(.a(G326), .O(gate82inter8));
  nand2 gate892(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate893(.a(s_49), .b(gate82inter3), .O(gate82inter10));
  nor2  gate894(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate895(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate896(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2465(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2466(.a(gate84inter0), .b(s_274), .O(gate84inter1));
  and2  gate2467(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2468(.a(s_274), .O(gate84inter3));
  inv1  gate2469(.a(s_275), .O(gate84inter4));
  nand2 gate2470(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2471(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2472(.a(G15), .O(gate84inter7));
  inv1  gate2473(.a(G329), .O(gate84inter8));
  nand2 gate2474(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2475(.a(s_275), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2476(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2477(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2478(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1415(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1416(.a(gate85inter0), .b(s_124), .O(gate85inter1));
  and2  gate1417(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1418(.a(s_124), .O(gate85inter3));
  inv1  gate1419(.a(s_125), .O(gate85inter4));
  nand2 gate1420(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1421(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1422(.a(G4), .O(gate85inter7));
  inv1  gate1423(.a(G332), .O(gate85inter8));
  nand2 gate1424(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1425(.a(s_125), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1426(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1427(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1428(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate617(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate618(.a(gate90inter0), .b(s_10), .O(gate90inter1));
  and2  gate619(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate620(.a(s_10), .O(gate90inter3));
  inv1  gate621(.a(s_11), .O(gate90inter4));
  nand2 gate622(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate623(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate624(.a(G21), .O(gate90inter7));
  inv1  gate625(.a(G338), .O(gate90inter8));
  nand2 gate626(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate627(.a(s_11), .b(gate90inter3), .O(gate90inter10));
  nor2  gate628(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate629(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate630(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1695(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1696(.a(gate93inter0), .b(s_164), .O(gate93inter1));
  and2  gate1697(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1698(.a(s_164), .O(gate93inter3));
  inv1  gate1699(.a(s_165), .O(gate93inter4));
  nand2 gate1700(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1701(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1702(.a(G18), .O(gate93inter7));
  inv1  gate1703(.a(G344), .O(gate93inter8));
  nand2 gate1704(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1705(.a(s_165), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1706(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1707(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1708(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1429(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1430(.a(gate96inter0), .b(s_126), .O(gate96inter1));
  and2  gate1431(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1432(.a(s_126), .O(gate96inter3));
  inv1  gate1433(.a(s_127), .O(gate96inter4));
  nand2 gate1434(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1435(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1436(.a(G30), .O(gate96inter7));
  inv1  gate1437(.a(G347), .O(gate96inter8));
  nand2 gate1438(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1439(.a(s_127), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1440(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1441(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1442(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1499(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1500(.a(gate101inter0), .b(s_136), .O(gate101inter1));
  and2  gate1501(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1502(.a(s_136), .O(gate101inter3));
  inv1  gate1503(.a(s_137), .O(gate101inter4));
  nand2 gate1504(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1505(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1506(.a(G20), .O(gate101inter7));
  inv1  gate1507(.a(G356), .O(gate101inter8));
  nand2 gate1508(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1509(.a(s_137), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1510(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1511(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1512(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2031(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2032(.a(gate110inter0), .b(s_212), .O(gate110inter1));
  and2  gate2033(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2034(.a(s_212), .O(gate110inter3));
  inv1  gate2035(.a(s_213), .O(gate110inter4));
  nand2 gate2036(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2037(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2038(.a(G372), .O(gate110inter7));
  inv1  gate2039(.a(G373), .O(gate110inter8));
  nand2 gate2040(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2041(.a(s_213), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2042(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2043(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2044(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1583(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1584(.a(gate113inter0), .b(s_148), .O(gate113inter1));
  and2  gate1585(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1586(.a(s_148), .O(gate113inter3));
  inv1  gate1587(.a(s_149), .O(gate113inter4));
  nand2 gate1588(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1589(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1590(.a(G378), .O(gate113inter7));
  inv1  gate1591(.a(G379), .O(gate113inter8));
  nand2 gate1592(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1593(.a(s_149), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1594(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1595(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1596(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate1037(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1038(.a(gate114inter0), .b(s_70), .O(gate114inter1));
  and2  gate1039(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1040(.a(s_70), .O(gate114inter3));
  inv1  gate1041(.a(s_71), .O(gate114inter4));
  nand2 gate1042(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1043(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1044(.a(G380), .O(gate114inter7));
  inv1  gate1045(.a(G381), .O(gate114inter8));
  nand2 gate1046(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1047(.a(s_71), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1048(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1049(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1050(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2521(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2522(.a(gate120inter0), .b(s_282), .O(gate120inter1));
  and2  gate2523(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2524(.a(s_282), .O(gate120inter3));
  inv1  gate2525(.a(s_283), .O(gate120inter4));
  nand2 gate2526(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2527(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2528(.a(G392), .O(gate120inter7));
  inv1  gate2529(.a(G393), .O(gate120inter8));
  nand2 gate2530(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2531(.a(s_283), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2532(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2533(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2534(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1485(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1486(.a(gate121inter0), .b(s_134), .O(gate121inter1));
  and2  gate1487(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1488(.a(s_134), .O(gate121inter3));
  inv1  gate1489(.a(s_135), .O(gate121inter4));
  nand2 gate1490(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1491(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1492(.a(G394), .O(gate121inter7));
  inv1  gate1493(.a(G395), .O(gate121inter8));
  nand2 gate1494(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1495(.a(s_135), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1496(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1497(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1498(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2269(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2270(.a(gate127inter0), .b(s_246), .O(gate127inter1));
  and2  gate2271(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2272(.a(s_246), .O(gate127inter3));
  inv1  gate2273(.a(s_247), .O(gate127inter4));
  nand2 gate2274(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2275(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2276(.a(G406), .O(gate127inter7));
  inv1  gate2277(.a(G407), .O(gate127inter8));
  nand2 gate2278(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2279(.a(s_247), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2280(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2281(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2282(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1079(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1080(.a(gate129inter0), .b(s_76), .O(gate129inter1));
  and2  gate1081(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1082(.a(s_76), .O(gate129inter3));
  inv1  gate1083(.a(s_77), .O(gate129inter4));
  nand2 gate1084(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1085(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1086(.a(G410), .O(gate129inter7));
  inv1  gate1087(.a(G411), .O(gate129inter8));
  nand2 gate1088(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1089(.a(s_77), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1090(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1091(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1092(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate995(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate996(.a(gate130inter0), .b(s_64), .O(gate130inter1));
  and2  gate997(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate998(.a(s_64), .O(gate130inter3));
  inv1  gate999(.a(s_65), .O(gate130inter4));
  nand2 gate1000(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1001(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1002(.a(G412), .O(gate130inter7));
  inv1  gate1003(.a(G413), .O(gate130inter8));
  nand2 gate1004(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1005(.a(s_65), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1006(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1007(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1008(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2577(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2578(.a(gate134inter0), .b(s_290), .O(gate134inter1));
  and2  gate2579(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2580(.a(s_290), .O(gate134inter3));
  inv1  gate2581(.a(s_291), .O(gate134inter4));
  nand2 gate2582(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2583(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2584(.a(G420), .O(gate134inter7));
  inv1  gate2585(.a(G421), .O(gate134inter8));
  nand2 gate2586(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2587(.a(s_291), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2588(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2589(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2590(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate799(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate800(.a(gate137inter0), .b(s_36), .O(gate137inter1));
  and2  gate801(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate802(.a(s_36), .O(gate137inter3));
  inv1  gate803(.a(s_37), .O(gate137inter4));
  nand2 gate804(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate805(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate806(.a(G426), .O(gate137inter7));
  inv1  gate807(.a(G429), .O(gate137inter8));
  nand2 gate808(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate809(.a(s_37), .b(gate137inter3), .O(gate137inter10));
  nor2  gate810(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate811(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate812(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2073(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2074(.a(gate139inter0), .b(s_218), .O(gate139inter1));
  and2  gate2075(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2076(.a(s_218), .O(gate139inter3));
  inv1  gate2077(.a(s_219), .O(gate139inter4));
  nand2 gate2078(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2079(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2080(.a(G438), .O(gate139inter7));
  inv1  gate2081(.a(G441), .O(gate139inter8));
  nand2 gate2082(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2083(.a(s_219), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2084(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2085(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2086(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2507(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2508(.a(gate146inter0), .b(s_280), .O(gate146inter1));
  and2  gate2509(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2510(.a(s_280), .O(gate146inter3));
  inv1  gate2511(.a(s_281), .O(gate146inter4));
  nand2 gate2512(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2513(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2514(.a(G480), .O(gate146inter7));
  inv1  gate2515(.a(G483), .O(gate146inter8));
  nand2 gate2516(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2517(.a(s_281), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2518(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2519(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2520(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1149(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1150(.a(gate151inter0), .b(s_86), .O(gate151inter1));
  and2  gate1151(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1152(.a(s_86), .O(gate151inter3));
  inv1  gate1153(.a(s_87), .O(gate151inter4));
  nand2 gate1154(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1155(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1156(.a(G510), .O(gate151inter7));
  inv1  gate1157(.a(G513), .O(gate151inter8));
  nand2 gate1158(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1159(.a(s_87), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1160(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1161(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1162(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1009(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1010(.a(gate155inter0), .b(s_66), .O(gate155inter1));
  and2  gate1011(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1012(.a(s_66), .O(gate155inter3));
  inv1  gate1013(.a(s_67), .O(gate155inter4));
  nand2 gate1014(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1015(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1016(.a(G432), .O(gate155inter7));
  inv1  gate1017(.a(G525), .O(gate155inter8));
  nand2 gate1018(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1019(.a(s_67), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1020(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1021(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1022(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1611(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1612(.a(gate157inter0), .b(s_152), .O(gate157inter1));
  and2  gate1613(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1614(.a(s_152), .O(gate157inter3));
  inv1  gate1615(.a(s_153), .O(gate157inter4));
  nand2 gate1616(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1617(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1618(.a(G438), .O(gate157inter7));
  inv1  gate1619(.a(G528), .O(gate157inter8));
  nand2 gate1620(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1621(.a(s_153), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1622(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1623(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1624(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2171(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2172(.a(gate158inter0), .b(s_232), .O(gate158inter1));
  and2  gate2173(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2174(.a(s_232), .O(gate158inter3));
  inv1  gate2175(.a(s_233), .O(gate158inter4));
  nand2 gate2176(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2177(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2178(.a(G441), .O(gate158inter7));
  inv1  gate2179(.a(G528), .O(gate158inter8));
  nand2 gate2180(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2181(.a(s_233), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2182(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2183(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2184(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate673(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate674(.a(gate159inter0), .b(s_18), .O(gate159inter1));
  and2  gate675(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate676(.a(s_18), .O(gate159inter3));
  inv1  gate677(.a(s_19), .O(gate159inter4));
  nand2 gate678(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate679(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate680(.a(G444), .O(gate159inter7));
  inv1  gate681(.a(G531), .O(gate159inter8));
  nand2 gate682(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate683(.a(s_19), .b(gate159inter3), .O(gate159inter10));
  nor2  gate684(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate685(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate686(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate743(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate744(.a(gate164inter0), .b(s_28), .O(gate164inter1));
  and2  gate745(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate746(.a(s_28), .O(gate164inter3));
  inv1  gate747(.a(s_29), .O(gate164inter4));
  nand2 gate748(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate749(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate750(.a(G459), .O(gate164inter7));
  inv1  gate751(.a(G537), .O(gate164inter8));
  nand2 gate752(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate753(.a(s_29), .b(gate164inter3), .O(gate164inter10));
  nor2  gate754(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate755(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate756(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate771(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate772(.a(gate165inter0), .b(s_32), .O(gate165inter1));
  and2  gate773(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate774(.a(s_32), .O(gate165inter3));
  inv1  gate775(.a(s_33), .O(gate165inter4));
  nand2 gate776(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate777(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate778(.a(G462), .O(gate165inter7));
  inv1  gate779(.a(G540), .O(gate165inter8));
  nand2 gate780(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate781(.a(s_33), .b(gate165inter3), .O(gate165inter10));
  nor2  gate782(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate783(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate784(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1359(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1360(.a(gate169inter0), .b(s_116), .O(gate169inter1));
  and2  gate1361(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1362(.a(s_116), .O(gate169inter3));
  inv1  gate1363(.a(s_117), .O(gate169inter4));
  nand2 gate1364(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1365(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1366(.a(G474), .O(gate169inter7));
  inv1  gate1367(.a(G546), .O(gate169inter8));
  nand2 gate1368(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1369(.a(s_117), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1370(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1371(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1372(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2563(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2564(.a(gate170inter0), .b(s_288), .O(gate170inter1));
  and2  gate2565(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2566(.a(s_288), .O(gate170inter3));
  inv1  gate2567(.a(s_289), .O(gate170inter4));
  nand2 gate2568(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2569(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2570(.a(G477), .O(gate170inter7));
  inv1  gate2571(.a(G546), .O(gate170inter8));
  nand2 gate2572(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2573(.a(s_289), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2574(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2575(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2576(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate757(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate758(.a(gate172inter0), .b(s_30), .O(gate172inter1));
  and2  gate759(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate760(.a(s_30), .O(gate172inter3));
  inv1  gate761(.a(s_31), .O(gate172inter4));
  nand2 gate762(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate763(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate764(.a(G483), .O(gate172inter7));
  inv1  gate765(.a(G549), .O(gate172inter8));
  nand2 gate766(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate767(.a(s_31), .b(gate172inter3), .O(gate172inter10));
  nor2  gate768(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate769(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate770(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1541(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1542(.a(gate174inter0), .b(s_142), .O(gate174inter1));
  and2  gate1543(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1544(.a(s_142), .O(gate174inter3));
  inv1  gate1545(.a(s_143), .O(gate174inter4));
  nand2 gate1546(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1547(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1548(.a(G489), .O(gate174inter7));
  inv1  gate1549(.a(G552), .O(gate174inter8));
  nand2 gate1550(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1551(.a(s_143), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1552(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1553(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1554(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1527(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1528(.a(gate179inter0), .b(s_140), .O(gate179inter1));
  and2  gate1529(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1530(.a(s_140), .O(gate179inter3));
  inv1  gate1531(.a(s_141), .O(gate179inter4));
  nand2 gate1532(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1533(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1534(.a(G504), .O(gate179inter7));
  inv1  gate1535(.a(G561), .O(gate179inter8));
  nand2 gate1536(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1537(.a(s_141), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1538(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1539(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1540(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2087(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2088(.a(gate182inter0), .b(s_220), .O(gate182inter1));
  and2  gate2089(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2090(.a(s_220), .O(gate182inter3));
  inv1  gate2091(.a(s_221), .O(gate182inter4));
  nand2 gate2092(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2093(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2094(.a(G513), .O(gate182inter7));
  inv1  gate2095(.a(G564), .O(gate182inter8));
  nand2 gate2096(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2097(.a(s_221), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2098(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2099(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2100(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate575(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate576(.a(gate183inter0), .b(s_4), .O(gate183inter1));
  and2  gate577(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate578(.a(s_4), .O(gate183inter3));
  inv1  gate579(.a(s_5), .O(gate183inter4));
  nand2 gate580(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate581(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate582(.a(G516), .O(gate183inter7));
  inv1  gate583(.a(G567), .O(gate183inter8));
  nand2 gate584(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate585(.a(s_5), .b(gate183inter3), .O(gate183inter10));
  nor2  gate586(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate587(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate588(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1513(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1514(.a(gate191inter0), .b(s_138), .O(gate191inter1));
  and2  gate1515(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1516(.a(s_138), .O(gate191inter3));
  inv1  gate1517(.a(s_139), .O(gate191inter4));
  nand2 gate1518(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1519(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1520(.a(G582), .O(gate191inter7));
  inv1  gate1521(.a(G583), .O(gate191inter8));
  nand2 gate1522(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1523(.a(s_139), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1524(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1525(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1526(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1345(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1346(.a(gate196inter0), .b(s_114), .O(gate196inter1));
  and2  gate1347(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1348(.a(s_114), .O(gate196inter3));
  inv1  gate1349(.a(s_115), .O(gate196inter4));
  nand2 gate1350(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1351(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1352(.a(G592), .O(gate196inter7));
  inv1  gate1353(.a(G593), .O(gate196inter8));
  nand2 gate1354(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1355(.a(s_115), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1356(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1357(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1358(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate645(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate646(.a(gate203inter0), .b(s_14), .O(gate203inter1));
  and2  gate647(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate648(.a(s_14), .O(gate203inter3));
  inv1  gate649(.a(s_15), .O(gate203inter4));
  nand2 gate650(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate651(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate652(.a(G602), .O(gate203inter7));
  inv1  gate653(.a(G612), .O(gate203inter8));
  nand2 gate654(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate655(.a(s_15), .b(gate203inter3), .O(gate203inter10));
  nor2  gate656(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate657(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate658(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1569(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1570(.a(gate207inter0), .b(s_146), .O(gate207inter1));
  and2  gate1571(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1572(.a(s_146), .O(gate207inter3));
  inv1  gate1573(.a(s_147), .O(gate207inter4));
  nand2 gate1574(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1575(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1576(.a(G622), .O(gate207inter7));
  inv1  gate1577(.a(G632), .O(gate207inter8));
  nand2 gate1578(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1579(.a(s_147), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1580(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1581(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1582(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2045(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2046(.a(gate209inter0), .b(s_214), .O(gate209inter1));
  and2  gate2047(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2048(.a(s_214), .O(gate209inter3));
  inv1  gate2049(.a(s_215), .O(gate209inter4));
  nand2 gate2050(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2051(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2052(.a(G602), .O(gate209inter7));
  inv1  gate2053(.a(G666), .O(gate209inter8));
  nand2 gate2054(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2055(.a(s_215), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2056(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2057(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2058(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2535(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2536(.a(gate211inter0), .b(s_284), .O(gate211inter1));
  and2  gate2537(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2538(.a(s_284), .O(gate211inter3));
  inv1  gate2539(.a(s_285), .O(gate211inter4));
  nand2 gate2540(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2541(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2542(.a(G612), .O(gate211inter7));
  inv1  gate2543(.a(G669), .O(gate211inter8));
  nand2 gate2544(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2545(.a(s_285), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2546(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2547(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2548(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1975(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1976(.a(gate215inter0), .b(s_204), .O(gate215inter1));
  and2  gate1977(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1978(.a(s_204), .O(gate215inter3));
  inv1  gate1979(.a(s_205), .O(gate215inter4));
  nand2 gate1980(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1981(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1982(.a(G607), .O(gate215inter7));
  inv1  gate1983(.a(G675), .O(gate215inter8));
  nand2 gate1984(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1985(.a(s_205), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1986(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1987(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1988(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2409(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2410(.a(gate217inter0), .b(s_266), .O(gate217inter1));
  and2  gate2411(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2412(.a(s_266), .O(gate217inter3));
  inv1  gate2413(.a(s_267), .O(gate217inter4));
  nand2 gate2414(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2415(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2416(.a(G622), .O(gate217inter7));
  inv1  gate2417(.a(G678), .O(gate217inter8));
  nand2 gate2418(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2419(.a(s_267), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2420(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2421(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2422(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1289(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1290(.a(gate218inter0), .b(s_106), .O(gate218inter1));
  and2  gate1291(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1292(.a(s_106), .O(gate218inter3));
  inv1  gate1293(.a(s_107), .O(gate218inter4));
  nand2 gate1294(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1295(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1296(.a(G627), .O(gate218inter7));
  inv1  gate1297(.a(G678), .O(gate218inter8));
  nand2 gate1298(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1299(.a(s_107), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1300(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1301(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1302(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2003(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2004(.a(gate219inter0), .b(s_208), .O(gate219inter1));
  and2  gate2005(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2006(.a(s_208), .O(gate219inter3));
  inv1  gate2007(.a(s_209), .O(gate219inter4));
  nand2 gate2008(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2009(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2010(.a(G632), .O(gate219inter7));
  inv1  gate2011(.a(G681), .O(gate219inter8));
  nand2 gate2012(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2013(.a(s_209), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2014(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2015(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2016(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1905(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1906(.a(gate220inter0), .b(s_194), .O(gate220inter1));
  and2  gate1907(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1908(.a(s_194), .O(gate220inter3));
  inv1  gate1909(.a(s_195), .O(gate220inter4));
  nand2 gate1910(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1911(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1912(.a(G637), .O(gate220inter7));
  inv1  gate1913(.a(G681), .O(gate220inter8));
  nand2 gate1914(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1915(.a(s_195), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1916(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1917(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1918(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2283(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2284(.a(gate222inter0), .b(s_248), .O(gate222inter1));
  and2  gate2285(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2286(.a(s_248), .O(gate222inter3));
  inv1  gate2287(.a(s_249), .O(gate222inter4));
  nand2 gate2288(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2289(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2290(.a(G632), .O(gate222inter7));
  inv1  gate2291(.a(G684), .O(gate222inter8));
  nand2 gate2292(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2293(.a(s_249), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2294(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2295(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2296(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1093(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1094(.a(gate228inter0), .b(s_78), .O(gate228inter1));
  and2  gate1095(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1096(.a(s_78), .O(gate228inter3));
  inv1  gate1097(.a(s_79), .O(gate228inter4));
  nand2 gate1098(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1099(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1100(.a(G696), .O(gate228inter7));
  inv1  gate1101(.a(G697), .O(gate228inter8));
  nand2 gate1102(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1103(.a(s_79), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1104(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1105(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1106(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1177(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1178(.a(gate231inter0), .b(s_90), .O(gate231inter1));
  and2  gate1179(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1180(.a(s_90), .O(gate231inter3));
  inv1  gate1181(.a(s_91), .O(gate231inter4));
  nand2 gate1182(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1183(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1184(.a(G702), .O(gate231inter7));
  inv1  gate1185(.a(G703), .O(gate231inter8));
  nand2 gate1186(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1187(.a(s_91), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1188(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1189(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1190(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1471(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1472(.a(gate234inter0), .b(s_132), .O(gate234inter1));
  and2  gate1473(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1474(.a(s_132), .O(gate234inter3));
  inv1  gate1475(.a(s_133), .O(gate234inter4));
  nand2 gate1476(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1477(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1478(.a(G245), .O(gate234inter7));
  inv1  gate1479(.a(G721), .O(gate234inter8));
  nand2 gate1480(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1481(.a(s_133), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1482(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1483(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1484(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate981(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate982(.a(gate237inter0), .b(s_62), .O(gate237inter1));
  and2  gate983(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate984(.a(s_62), .O(gate237inter3));
  inv1  gate985(.a(s_63), .O(gate237inter4));
  nand2 gate986(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate987(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate988(.a(G254), .O(gate237inter7));
  inv1  gate989(.a(G706), .O(gate237inter8));
  nand2 gate990(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate991(.a(s_63), .b(gate237inter3), .O(gate237inter10));
  nor2  gate992(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate993(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate994(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1065(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1066(.a(gate242inter0), .b(s_74), .O(gate242inter1));
  and2  gate1067(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1068(.a(s_74), .O(gate242inter3));
  inv1  gate1069(.a(s_75), .O(gate242inter4));
  nand2 gate1070(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1071(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1072(.a(G718), .O(gate242inter7));
  inv1  gate1073(.a(G730), .O(gate242inter8));
  nand2 gate1074(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1075(.a(s_75), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1076(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1077(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1078(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1107(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1108(.a(gate247inter0), .b(s_80), .O(gate247inter1));
  and2  gate1109(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1110(.a(s_80), .O(gate247inter3));
  inv1  gate1111(.a(s_81), .O(gate247inter4));
  nand2 gate1112(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1113(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1114(.a(G251), .O(gate247inter7));
  inv1  gate1115(.a(G739), .O(gate247inter8));
  nand2 gate1116(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1117(.a(s_81), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1118(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1119(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1120(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate911(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate912(.a(gate260inter0), .b(s_52), .O(gate260inter1));
  and2  gate913(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate914(.a(s_52), .O(gate260inter3));
  inv1  gate915(.a(s_53), .O(gate260inter4));
  nand2 gate916(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate917(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate918(.a(G760), .O(gate260inter7));
  inv1  gate919(.a(G761), .O(gate260inter8));
  nand2 gate920(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate921(.a(s_53), .b(gate260inter3), .O(gate260inter10));
  nor2  gate922(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate923(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate924(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2353(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2354(.a(gate265inter0), .b(s_258), .O(gate265inter1));
  and2  gate2355(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2356(.a(s_258), .O(gate265inter3));
  inv1  gate2357(.a(s_259), .O(gate265inter4));
  nand2 gate2358(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2359(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2360(.a(G642), .O(gate265inter7));
  inv1  gate2361(.a(G770), .O(gate265inter8));
  nand2 gate2362(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2363(.a(s_259), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2364(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2365(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2366(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate953(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate954(.a(gate270inter0), .b(s_58), .O(gate270inter1));
  and2  gate955(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate956(.a(s_58), .O(gate270inter3));
  inv1  gate957(.a(s_59), .O(gate270inter4));
  nand2 gate958(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate959(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate960(.a(G657), .O(gate270inter7));
  inv1  gate961(.a(G785), .O(gate270inter8));
  nand2 gate962(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate963(.a(s_59), .b(gate270inter3), .O(gate270inter10));
  nor2  gate964(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate965(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate966(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2143(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2144(.a(gate273inter0), .b(s_228), .O(gate273inter1));
  and2  gate2145(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2146(.a(s_228), .O(gate273inter3));
  inv1  gate2147(.a(s_229), .O(gate273inter4));
  nand2 gate2148(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2149(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2150(.a(G642), .O(gate273inter7));
  inv1  gate2151(.a(G794), .O(gate273inter8));
  nand2 gate2152(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2153(.a(s_229), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2154(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2155(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2156(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1275(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1276(.a(gate275inter0), .b(s_104), .O(gate275inter1));
  and2  gate1277(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1278(.a(s_104), .O(gate275inter3));
  inv1  gate1279(.a(s_105), .O(gate275inter4));
  nand2 gate1280(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1281(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1282(.a(G645), .O(gate275inter7));
  inv1  gate1283(.a(G797), .O(gate275inter8));
  nand2 gate1284(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1285(.a(s_105), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1286(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1287(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1288(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate2423(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2424(.a(gate276inter0), .b(s_268), .O(gate276inter1));
  and2  gate2425(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2426(.a(s_268), .O(gate276inter3));
  inv1  gate2427(.a(s_269), .O(gate276inter4));
  nand2 gate2428(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2429(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2430(.a(G773), .O(gate276inter7));
  inv1  gate2431(.a(G797), .O(gate276inter8));
  nand2 gate2432(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2433(.a(s_269), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2434(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2435(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2436(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1191(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1192(.a(gate278inter0), .b(s_92), .O(gate278inter1));
  and2  gate1193(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1194(.a(s_92), .O(gate278inter3));
  inv1  gate1195(.a(s_93), .O(gate278inter4));
  nand2 gate1196(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1197(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1198(.a(G776), .O(gate278inter7));
  inv1  gate1199(.a(G800), .O(gate278inter8));
  nand2 gate1200(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1201(.a(s_93), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1202(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1203(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1204(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1555(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1556(.a(gate280inter0), .b(s_144), .O(gate280inter1));
  and2  gate1557(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1558(.a(s_144), .O(gate280inter3));
  inv1  gate1559(.a(s_145), .O(gate280inter4));
  nand2 gate1560(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1561(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1562(.a(G779), .O(gate280inter7));
  inv1  gate1563(.a(G803), .O(gate280inter8));
  nand2 gate1564(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1565(.a(s_145), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1566(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1567(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1568(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate897(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate898(.a(gate283inter0), .b(s_50), .O(gate283inter1));
  and2  gate899(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate900(.a(s_50), .O(gate283inter3));
  inv1  gate901(.a(s_51), .O(gate283inter4));
  nand2 gate902(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate903(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate904(.a(G657), .O(gate283inter7));
  inv1  gate905(.a(G809), .O(gate283inter8));
  nand2 gate906(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate907(.a(s_51), .b(gate283inter3), .O(gate283inter10));
  nor2  gate908(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate909(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate910(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1331(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1332(.a(gate287inter0), .b(s_112), .O(gate287inter1));
  and2  gate1333(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1334(.a(s_112), .O(gate287inter3));
  inv1  gate1335(.a(s_113), .O(gate287inter4));
  nand2 gate1336(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1337(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1338(.a(G663), .O(gate287inter7));
  inv1  gate1339(.a(G815), .O(gate287inter8));
  nand2 gate1340(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1341(.a(s_113), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1342(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1343(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1344(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2367(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2368(.a(gate290inter0), .b(s_260), .O(gate290inter1));
  and2  gate2369(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2370(.a(s_260), .O(gate290inter3));
  inv1  gate2371(.a(s_261), .O(gate290inter4));
  nand2 gate2372(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2373(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2374(.a(G820), .O(gate290inter7));
  inv1  gate2375(.a(G821), .O(gate290inter8));
  nand2 gate2376(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2377(.a(s_261), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2378(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2379(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2380(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1933(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1934(.a(gate293inter0), .b(s_198), .O(gate293inter1));
  and2  gate1935(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1936(.a(s_198), .O(gate293inter3));
  inv1  gate1937(.a(s_199), .O(gate293inter4));
  nand2 gate1938(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1939(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1940(.a(G828), .O(gate293inter7));
  inv1  gate1941(.a(G829), .O(gate293inter8));
  nand2 gate1942(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1943(.a(s_199), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1944(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1945(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1946(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1317(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1318(.a(gate294inter0), .b(s_110), .O(gate294inter1));
  and2  gate1319(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1320(.a(s_110), .O(gate294inter3));
  inv1  gate1321(.a(s_111), .O(gate294inter4));
  nand2 gate1322(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1323(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1324(.a(G832), .O(gate294inter7));
  inv1  gate1325(.a(G833), .O(gate294inter8));
  nand2 gate1326(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1327(.a(s_111), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1328(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1329(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1330(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1681(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1682(.a(gate388inter0), .b(s_162), .O(gate388inter1));
  and2  gate1683(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1684(.a(s_162), .O(gate388inter3));
  inv1  gate1685(.a(s_163), .O(gate388inter4));
  nand2 gate1686(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1687(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1688(.a(G2), .O(gate388inter7));
  inv1  gate1689(.a(G1039), .O(gate388inter8));
  nand2 gate1690(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1691(.a(s_163), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1692(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1693(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1694(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1751(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1752(.a(gate390inter0), .b(s_172), .O(gate390inter1));
  and2  gate1753(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1754(.a(s_172), .O(gate390inter3));
  inv1  gate1755(.a(s_173), .O(gate390inter4));
  nand2 gate1756(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1757(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1758(.a(G4), .O(gate390inter7));
  inv1  gate1759(.a(G1045), .O(gate390inter8));
  nand2 gate1760(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1761(.a(s_173), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1762(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1763(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1764(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate547(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate548(.a(gate391inter0), .b(s_0), .O(gate391inter1));
  and2  gate549(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate550(.a(s_0), .O(gate391inter3));
  inv1  gate551(.a(s_1), .O(gate391inter4));
  nand2 gate552(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate553(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate554(.a(G5), .O(gate391inter7));
  inv1  gate555(.a(G1048), .O(gate391inter8));
  nand2 gate556(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate557(.a(s_1), .b(gate391inter3), .O(gate391inter10));
  nor2  gate558(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate559(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate560(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1835(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1836(.a(gate397inter0), .b(s_184), .O(gate397inter1));
  and2  gate1837(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1838(.a(s_184), .O(gate397inter3));
  inv1  gate1839(.a(s_185), .O(gate397inter4));
  nand2 gate1840(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1841(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1842(.a(G11), .O(gate397inter7));
  inv1  gate1843(.a(G1066), .O(gate397inter8));
  nand2 gate1844(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1845(.a(s_185), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1846(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1847(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1848(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1163(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1164(.a(gate399inter0), .b(s_88), .O(gate399inter1));
  and2  gate1165(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1166(.a(s_88), .O(gate399inter3));
  inv1  gate1167(.a(s_89), .O(gate399inter4));
  nand2 gate1168(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1169(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1170(.a(G13), .O(gate399inter7));
  inv1  gate1171(.a(G1072), .O(gate399inter8));
  nand2 gate1172(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1173(.a(s_89), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1174(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1175(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1176(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate813(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate814(.a(gate400inter0), .b(s_38), .O(gate400inter1));
  and2  gate815(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate816(.a(s_38), .O(gate400inter3));
  inv1  gate817(.a(s_39), .O(gate400inter4));
  nand2 gate818(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate819(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate820(.a(G14), .O(gate400inter7));
  inv1  gate821(.a(G1075), .O(gate400inter8));
  nand2 gate822(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate823(.a(s_39), .b(gate400inter3), .O(gate400inter10));
  nor2  gate824(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate825(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate826(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1387(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1388(.a(gate402inter0), .b(s_120), .O(gate402inter1));
  and2  gate1389(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1390(.a(s_120), .O(gate402inter3));
  inv1  gate1391(.a(s_121), .O(gate402inter4));
  nand2 gate1392(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1393(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1394(.a(G16), .O(gate402inter7));
  inv1  gate1395(.a(G1081), .O(gate402inter8));
  nand2 gate1396(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1397(.a(s_121), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1398(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1399(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1400(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1737(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1738(.a(gate405inter0), .b(s_170), .O(gate405inter1));
  and2  gate1739(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1740(.a(s_170), .O(gate405inter3));
  inv1  gate1741(.a(s_171), .O(gate405inter4));
  nand2 gate1742(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1743(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1744(.a(G19), .O(gate405inter7));
  inv1  gate1745(.a(G1090), .O(gate405inter8));
  nand2 gate1746(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1747(.a(s_171), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1748(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1749(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1750(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1597(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1598(.a(gate408inter0), .b(s_150), .O(gate408inter1));
  and2  gate1599(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1600(.a(s_150), .O(gate408inter3));
  inv1  gate1601(.a(s_151), .O(gate408inter4));
  nand2 gate1602(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1603(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1604(.a(G22), .O(gate408inter7));
  inv1  gate1605(.a(G1099), .O(gate408inter8));
  nand2 gate1606(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1607(.a(s_151), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1608(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1609(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1610(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1667(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1668(.a(gate411inter0), .b(s_160), .O(gate411inter1));
  and2  gate1669(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1670(.a(s_160), .O(gate411inter3));
  inv1  gate1671(.a(s_161), .O(gate411inter4));
  nand2 gate1672(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1673(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1674(.a(G25), .O(gate411inter7));
  inv1  gate1675(.a(G1108), .O(gate411inter8));
  nand2 gate1676(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1677(.a(s_161), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1678(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1679(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1680(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1261(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1262(.a(gate413inter0), .b(s_102), .O(gate413inter1));
  and2  gate1263(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1264(.a(s_102), .O(gate413inter3));
  inv1  gate1265(.a(s_103), .O(gate413inter4));
  nand2 gate1266(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1267(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1268(.a(G27), .O(gate413inter7));
  inv1  gate1269(.a(G1114), .O(gate413inter8));
  nand2 gate1270(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1271(.a(s_103), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1272(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1273(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1274(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1653(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1654(.a(gate418inter0), .b(s_158), .O(gate418inter1));
  and2  gate1655(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1656(.a(s_158), .O(gate418inter3));
  inv1  gate1657(.a(s_159), .O(gate418inter4));
  nand2 gate1658(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1659(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1660(.a(G32), .O(gate418inter7));
  inv1  gate1661(.a(G1129), .O(gate418inter8));
  nand2 gate1662(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1663(.a(s_159), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1664(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1665(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1666(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate729(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate730(.a(gate422inter0), .b(s_26), .O(gate422inter1));
  and2  gate731(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate732(.a(s_26), .O(gate422inter3));
  inv1  gate733(.a(s_27), .O(gate422inter4));
  nand2 gate734(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate735(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate736(.a(G1039), .O(gate422inter7));
  inv1  gate737(.a(G1135), .O(gate422inter8));
  nand2 gate738(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate739(.a(s_27), .b(gate422inter3), .O(gate422inter10));
  nor2  gate740(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate741(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate742(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate631(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate632(.a(gate424inter0), .b(s_12), .O(gate424inter1));
  and2  gate633(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate634(.a(s_12), .O(gate424inter3));
  inv1  gate635(.a(s_13), .O(gate424inter4));
  nand2 gate636(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate637(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate638(.a(G1042), .O(gate424inter7));
  inv1  gate639(.a(G1138), .O(gate424inter8));
  nand2 gate640(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate641(.a(s_13), .b(gate424inter3), .O(gate424inter10));
  nor2  gate642(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate643(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate644(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1373(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1374(.a(gate425inter0), .b(s_118), .O(gate425inter1));
  and2  gate1375(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1376(.a(s_118), .O(gate425inter3));
  inv1  gate1377(.a(s_119), .O(gate425inter4));
  nand2 gate1378(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1379(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1380(.a(G4), .O(gate425inter7));
  inv1  gate1381(.a(G1141), .O(gate425inter8));
  nand2 gate1382(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1383(.a(s_119), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1384(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1385(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1386(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2115(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2116(.a(gate427inter0), .b(s_224), .O(gate427inter1));
  and2  gate2117(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2118(.a(s_224), .O(gate427inter3));
  inv1  gate2119(.a(s_225), .O(gate427inter4));
  nand2 gate2120(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2121(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2122(.a(G5), .O(gate427inter7));
  inv1  gate2123(.a(G1144), .O(gate427inter8));
  nand2 gate2124(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2125(.a(s_225), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2126(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2127(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2128(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1863(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1864(.a(gate429inter0), .b(s_188), .O(gate429inter1));
  and2  gate1865(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1866(.a(s_188), .O(gate429inter3));
  inv1  gate1867(.a(s_189), .O(gate429inter4));
  nand2 gate1868(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1869(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1870(.a(G6), .O(gate429inter7));
  inv1  gate1871(.a(G1147), .O(gate429inter8));
  nand2 gate1872(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1873(.a(s_189), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1874(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1875(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1876(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1849(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1850(.a(gate430inter0), .b(s_186), .O(gate430inter1));
  and2  gate1851(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1852(.a(s_186), .O(gate430inter3));
  inv1  gate1853(.a(s_187), .O(gate430inter4));
  nand2 gate1854(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1855(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1856(.a(G1051), .O(gate430inter7));
  inv1  gate1857(.a(G1147), .O(gate430inter8));
  nand2 gate1858(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1859(.a(s_187), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1860(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1861(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1862(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1303(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1304(.a(gate431inter0), .b(s_108), .O(gate431inter1));
  and2  gate1305(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1306(.a(s_108), .O(gate431inter3));
  inv1  gate1307(.a(s_109), .O(gate431inter4));
  nand2 gate1308(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1309(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1310(.a(G7), .O(gate431inter7));
  inv1  gate1311(.a(G1150), .O(gate431inter8));
  nand2 gate1312(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1313(.a(s_109), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1314(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1315(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1316(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1625(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1626(.a(gate441inter0), .b(s_154), .O(gate441inter1));
  and2  gate1627(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1628(.a(s_154), .O(gate441inter3));
  inv1  gate1629(.a(s_155), .O(gate441inter4));
  nand2 gate1630(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1631(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1632(.a(G12), .O(gate441inter7));
  inv1  gate1633(.a(G1165), .O(gate441inter8));
  nand2 gate1634(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1635(.a(s_155), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1636(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1637(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1638(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2059(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2060(.a(gate445inter0), .b(s_216), .O(gate445inter1));
  and2  gate2061(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2062(.a(s_216), .O(gate445inter3));
  inv1  gate2063(.a(s_217), .O(gate445inter4));
  nand2 gate2064(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2065(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2066(.a(G14), .O(gate445inter7));
  inv1  gate2067(.a(G1171), .O(gate445inter8));
  nand2 gate2068(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2069(.a(s_217), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2070(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2071(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2072(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1401(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1402(.a(gate447inter0), .b(s_122), .O(gate447inter1));
  and2  gate1403(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1404(.a(s_122), .O(gate447inter3));
  inv1  gate1405(.a(s_123), .O(gate447inter4));
  nand2 gate1406(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1407(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1408(.a(G15), .O(gate447inter7));
  inv1  gate1409(.a(G1174), .O(gate447inter8));
  nand2 gate1410(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1411(.a(s_123), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1412(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1413(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1414(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1219(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1220(.a(gate449inter0), .b(s_96), .O(gate449inter1));
  and2  gate1221(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1222(.a(s_96), .O(gate449inter3));
  inv1  gate1223(.a(s_97), .O(gate449inter4));
  nand2 gate1224(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1225(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1226(.a(G16), .O(gate449inter7));
  inv1  gate1227(.a(G1177), .O(gate449inter8));
  nand2 gate1228(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1229(.a(s_97), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1230(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1231(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1232(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1121(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1122(.a(gate455inter0), .b(s_82), .O(gate455inter1));
  and2  gate1123(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1124(.a(s_82), .O(gate455inter3));
  inv1  gate1125(.a(s_83), .O(gate455inter4));
  nand2 gate1126(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1127(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1128(.a(G19), .O(gate455inter7));
  inv1  gate1129(.a(G1186), .O(gate455inter8));
  nand2 gate1130(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1131(.a(s_83), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1132(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1133(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1134(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate687(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate688(.a(gate457inter0), .b(s_20), .O(gate457inter1));
  and2  gate689(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate690(.a(s_20), .O(gate457inter3));
  inv1  gate691(.a(s_21), .O(gate457inter4));
  nand2 gate692(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate693(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate694(.a(G20), .O(gate457inter7));
  inv1  gate695(.a(G1189), .O(gate457inter8));
  nand2 gate696(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate697(.a(s_21), .b(gate457inter3), .O(gate457inter10));
  nor2  gate698(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate699(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate700(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate785(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate786(.a(gate459inter0), .b(s_34), .O(gate459inter1));
  and2  gate787(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate788(.a(s_34), .O(gate459inter3));
  inv1  gate789(.a(s_35), .O(gate459inter4));
  nand2 gate790(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate791(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate792(.a(G21), .O(gate459inter7));
  inv1  gate793(.a(G1192), .O(gate459inter8));
  nand2 gate794(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate795(.a(s_35), .b(gate459inter3), .O(gate459inter10));
  nor2  gate796(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate797(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate798(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2395(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2396(.a(gate464inter0), .b(s_264), .O(gate464inter1));
  and2  gate2397(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2398(.a(s_264), .O(gate464inter3));
  inv1  gate2399(.a(s_265), .O(gate464inter4));
  nand2 gate2400(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2401(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2402(.a(G1102), .O(gate464inter7));
  inv1  gate2403(.a(G1198), .O(gate464inter8));
  nand2 gate2404(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2405(.a(s_265), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2406(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2407(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2408(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate925(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate926(.a(gate465inter0), .b(s_54), .O(gate465inter1));
  and2  gate927(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate928(.a(s_54), .O(gate465inter3));
  inv1  gate929(.a(s_55), .O(gate465inter4));
  nand2 gate930(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate931(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate932(.a(G24), .O(gate465inter7));
  inv1  gate933(.a(G1201), .O(gate465inter8));
  nand2 gate934(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate935(.a(s_55), .b(gate465inter3), .O(gate465inter10));
  nor2  gate936(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate937(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate938(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1821(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1822(.a(gate466inter0), .b(s_182), .O(gate466inter1));
  and2  gate1823(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1824(.a(s_182), .O(gate466inter3));
  inv1  gate1825(.a(s_183), .O(gate466inter4));
  nand2 gate1826(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1827(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1828(.a(G1105), .O(gate466inter7));
  inv1  gate1829(.a(G1201), .O(gate466inter8));
  nand2 gate1830(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1831(.a(s_183), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1832(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1833(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1834(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2451(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2452(.a(gate472inter0), .b(s_272), .O(gate472inter1));
  and2  gate2453(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2454(.a(s_272), .O(gate472inter3));
  inv1  gate2455(.a(s_273), .O(gate472inter4));
  nand2 gate2456(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2457(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2458(.a(G1114), .O(gate472inter7));
  inv1  gate2459(.a(G1210), .O(gate472inter8));
  nand2 gate2460(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2461(.a(s_273), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2462(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2463(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2464(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1765(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1766(.a(gate474inter0), .b(s_174), .O(gate474inter1));
  and2  gate1767(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1768(.a(s_174), .O(gate474inter3));
  inv1  gate1769(.a(s_175), .O(gate474inter4));
  nand2 gate1770(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1771(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1772(.a(G1117), .O(gate474inter7));
  inv1  gate1773(.a(G1213), .O(gate474inter8));
  nand2 gate1774(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1775(.a(s_175), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1776(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1777(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1778(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2479(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2480(.a(gate476inter0), .b(s_276), .O(gate476inter1));
  and2  gate2481(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2482(.a(s_276), .O(gate476inter3));
  inv1  gate2483(.a(s_277), .O(gate476inter4));
  nand2 gate2484(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2485(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2486(.a(G1120), .O(gate476inter7));
  inv1  gate2487(.a(G1216), .O(gate476inter8));
  nand2 gate2488(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2489(.a(s_277), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2490(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2491(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2492(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2549(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2550(.a(gate480inter0), .b(s_286), .O(gate480inter1));
  and2  gate2551(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2552(.a(s_286), .O(gate480inter3));
  inv1  gate2553(.a(s_287), .O(gate480inter4));
  nand2 gate2554(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2555(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2556(.a(G1126), .O(gate480inter7));
  inv1  gate2557(.a(G1222), .O(gate480inter8));
  nand2 gate2558(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2559(.a(s_287), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2560(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2561(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2562(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1457(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1458(.a(gate482inter0), .b(s_130), .O(gate482inter1));
  and2  gate1459(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1460(.a(s_130), .O(gate482inter3));
  inv1  gate1461(.a(s_131), .O(gate482inter4));
  nand2 gate1462(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1463(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1464(.a(G1129), .O(gate482inter7));
  inv1  gate1465(.a(G1225), .O(gate482inter8));
  nand2 gate1466(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1467(.a(s_131), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1468(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1469(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1470(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate2129(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2130(.a(gate484inter0), .b(s_226), .O(gate484inter1));
  and2  gate2131(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2132(.a(s_226), .O(gate484inter3));
  inv1  gate2133(.a(s_227), .O(gate484inter4));
  nand2 gate2134(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2135(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2136(.a(G1230), .O(gate484inter7));
  inv1  gate2137(.a(G1231), .O(gate484inter8));
  nand2 gate2138(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2139(.a(s_227), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2140(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2141(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2142(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1919(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1920(.a(gate485inter0), .b(s_196), .O(gate485inter1));
  and2  gate1921(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1922(.a(s_196), .O(gate485inter3));
  inv1  gate1923(.a(s_197), .O(gate485inter4));
  nand2 gate1924(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1925(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1926(.a(G1232), .O(gate485inter7));
  inv1  gate1927(.a(G1233), .O(gate485inter8));
  nand2 gate1928(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1929(.a(s_197), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1930(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1931(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1932(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2437(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2438(.a(gate488inter0), .b(s_270), .O(gate488inter1));
  and2  gate2439(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2440(.a(s_270), .O(gate488inter3));
  inv1  gate2441(.a(s_271), .O(gate488inter4));
  nand2 gate2442(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2443(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2444(.a(G1238), .O(gate488inter7));
  inv1  gate2445(.a(G1239), .O(gate488inter8));
  nand2 gate2446(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2447(.a(s_271), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2448(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2449(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2450(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1793(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1794(.a(gate489inter0), .b(s_178), .O(gate489inter1));
  and2  gate1795(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1796(.a(s_178), .O(gate489inter3));
  inv1  gate1797(.a(s_179), .O(gate489inter4));
  nand2 gate1798(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1799(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1800(.a(G1240), .O(gate489inter7));
  inv1  gate1801(.a(G1241), .O(gate489inter8));
  nand2 gate1802(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1803(.a(s_179), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1804(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1805(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1806(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2325(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2326(.a(gate491inter0), .b(s_254), .O(gate491inter1));
  and2  gate2327(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2328(.a(s_254), .O(gate491inter3));
  inv1  gate2329(.a(s_255), .O(gate491inter4));
  nand2 gate2330(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2331(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2332(.a(G1244), .O(gate491inter7));
  inv1  gate2333(.a(G1245), .O(gate491inter8));
  nand2 gate2334(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2335(.a(s_255), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2336(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2337(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2338(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2185(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2186(.a(gate497inter0), .b(s_234), .O(gate497inter1));
  and2  gate2187(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2188(.a(s_234), .O(gate497inter3));
  inv1  gate2189(.a(s_235), .O(gate497inter4));
  nand2 gate2190(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2191(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2192(.a(G1256), .O(gate497inter7));
  inv1  gate2193(.a(G1257), .O(gate497inter8));
  nand2 gate2194(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2195(.a(s_235), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2196(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2197(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2198(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate589(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate590(.a(gate500inter0), .b(s_6), .O(gate500inter1));
  and2  gate591(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate592(.a(s_6), .O(gate500inter3));
  inv1  gate593(.a(s_7), .O(gate500inter4));
  nand2 gate594(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate595(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate596(.a(G1262), .O(gate500inter7));
  inv1  gate597(.a(G1263), .O(gate500inter8));
  nand2 gate598(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate599(.a(s_7), .b(gate500inter3), .O(gate500inter10));
  nor2  gate600(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate601(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate602(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1233(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1234(.a(gate501inter0), .b(s_98), .O(gate501inter1));
  and2  gate1235(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1236(.a(s_98), .O(gate501inter3));
  inv1  gate1237(.a(s_99), .O(gate501inter4));
  nand2 gate1238(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1239(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1240(.a(G1264), .O(gate501inter7));
  inv1  gate1241(.a(G1265), .O(gate501inter8));
  nand2 gate1242(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1243(.a(s_99), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1244(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1245(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1246(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2311(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2312(.a(gate503inter0), .b(s_252), .O(gate503inter1));
  and2  gate2313(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2314(.a(s_252), .O(gate503inter3));
  inv1  gate2315(.a(s_253), .O(gate503inter4));
  nand2 gate2316(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2317(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2318(.a(G1268), .O(gate503inter7));
  inv1  gate2319(.a(G1269), .O(gate503inter8));
  nand2 gate2320(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2321(.a(s_253), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2322(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2323(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2324(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate967(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate968(.a(gate505inter0), .b(s_60), .O(gate505inter1));
  and2  gate969(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate970(.a(s_60), .O(gate505inter3));
  inv1  gate971(.a(s_61), .O(gate505inter4));
  nand2 gate972(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate973(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate974(.a(G1272), .O(gate505inter7));
  inv1  gate975(.a(G1273), .O(gate505inter8));
  nand2 gate976(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate977(.a(s_61), .b(gate505inter3), .O(gate505inter10));
  nor2  gate978(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate979(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate980(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2339(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2340(.a(gate507inter0), .b(s_256), .O(gate507inter1));
  and2  gate2341(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2342(.a(s_256), .O(gate507inter3));
  inv1  gate2343(.a(s_257), .O(gate507inter4));
  nand2 gate2344(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2345(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2346(.a(G1276), .O(gate507inter7));
  inv1  gate2347(.a(G1277), .O(gate507inter8));
  nand2 gate2348(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2349(.a(s_257), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2350(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2351(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2352(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1877(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1878(.a(gate508inter0), .b(s_190), .O(gate508inter1));
  and2  gate1879(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1880(.a(s_190), .O(gate508inter3));
  inv1  gate1881(.a(s_191), .O(gate508inter4));
  nand2 gate1882(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1883(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1884(.a(G1278), .O(gate508inter7));
  inv1  gate1885(.a(G1279), .O(gate508inter8));
  nand2 gate1886(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1887(.a(s_191), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1888(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1889(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1890(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate827(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate828(.a(gate513inter0), .b(s_40), .O(gate513inter1));
  and2  gate829(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate830(.a(s_40), .O(gate513inter3));
  inv1  gate831(.a(s_41), .O(gate513inter4));
  nand2 gate832(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate833(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate834(.a(G1288), .O(gate513inter7));
  inv1  gate835(.a(G1289), .O(gate513inter8));
  nand2 gate836(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate837(.a(s_41), .b(gate513inter3), .O(gate513inter10));
  nor2  gate838(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate839(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate840(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule