module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate315(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate316(.a(gate19inter0), .b(s_22), .O(gate19inter1));
  and2  gate317(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate318(.a(s_22), .O(gate19inter3));
  inv1  gate319(.a(s_23), .O(gate19inter4));
  nand2 gate320(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate321(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate322(.a(N118), .O(gate19inter7));
  inv1  gate323(.a(N4), .O(gate19inter8));
  nand2 gate324(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate325(.a(s_23), .b(gate19inter3), .O(gate19inter10));
  nor2  gate326(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate327(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate328(.a(gate19inter12), .b(gate19inter1), .O(N154));
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate581(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate582(.a(gate29inter0), .b(s_60), .O(gate29inter1));
  and2  gate583(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate584(.a(s_60), .O(gate29inter3));
  inv1  gate585(.a(s_61), .O(gate29inter4));
  nand2 gate586(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate587(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate588(.a(N150), .O(gate29inter7));
  inv1  gate589(.a(N108), .O(gate29inter8));
  nand2 gate590(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate591(.a(s_61), .b(gate29inter3), .O(gate29inter10));
  nor2  gate592(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate593(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate594(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );

  xor2  gate189(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate190(.a(gate31inter0), .b(s_4), .O(gate31inter1));
  and2  gate191(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate192(.a(s_4), .O(gate31inter3));
  inv1  gate193(.a(s_5), .O(gate31inter4));
  nand2 gate194(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate195(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate196(.a(N27), .O(gate31inter7));
  inv1  gate197(.a(N123), .O(gate31inter8));
  nand2 gate198(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate199(.a(s_5), .b(gate31inter3), .O(gate31inter10));
  nor2  gate200(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate201(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate202(.a(gate31inter12), .b(gate31inter1), .O(N184));

  xor2  gate595(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate596(.a(gate32inter0), .b(s_62), .O(gate32inter1));
  and2  gate597(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate598(.a(s_62), .O(gate32inter3));
  inv1  gate599(.a(s_63), .O(gate32inter4));
  nand2 gate600(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate601(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate602(.a(N34), .O(gate32inter7));
  inv1  gate603(.a(N127), .O(gate32inter8));
  nand2 gate604(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate605(.a(s_63), .b(gate32inter3), .O(gate32inter10));
  nor2  gate606(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate607(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate608(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate413(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate414(.a(gate38inter0), .b(s_36), .O(gate38inter1));
  and2  gate415(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate416(.a(s_36), .O(gate38inter3));
  inv1  gate417(.a(s_37), .O(gate38inter4));
  nand2 gate418(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate419(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate420(.a(N73), .O(gate38inter7));
  inv1  gate421(.a(N139), .O(gate38inter8));
  nand2 gate422(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate423(.a(s_37), .b(gate38inter3), .O(gate38inter10));
  nor2  gate424(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate425(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate426(.a(gate38inter12), .b(gate38inter1), .O(N191));
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate427(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate428(.a(gate40inter0), .b(s_38), .O(gate40inter1));
  and2  gate429(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate430(.a(s_38), .O(gate40inter3));
  inv1  gate431(.a(s_39), .O(gate40inter4));
  nand2 gate432(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate433(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate434(.a(N86), .O(gate40inter7));
  inv1  gate435(.a(N143), .O(gate40inter8));
  nand2 gate436(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate437(.a(s_39), .b(gate40inter3), .O(gate40inter10));
  nor2  gate438(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate439(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate440(.a(gate40inter12), .b(gate40inter1), .O(N193));
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );

  xor2  gate455(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate456(.a(gate45inter0), .b(s_42), .O(gate45inter1));
  and2  gate457(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate458(.a(s_42), .O(gate45inter3));
  inv1  gate459(.a(s_43), .O(gate45inter4));
  nand2 gate460(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate461(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate462(.a(N115), .O(gate45inter7));
  inv1  gate463(.a(N151), .O(gate45inter8));
  nand2 gate464(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate465(.a(s_43), .b(gate45inter3), .O(gate45inter10));
  nor2  gate466(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate467(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate468(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );

  xor2  gate357(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate358(.a(gate51inter0), .b(s_28), .O(gate51inter1));
  and2  gate359(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate360(.a(s_28), .O(gate51inter3));
  inv1  gate361(.a(s_29), .O(gate51inter4));
  nand2 gate362(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate363(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate364(.a(N203), .O(gate51inter7));
  inv1  gate365(.a(N159), .O(gate51inter8));
  nand2 gate366(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate367(.a(s_29), .b(gate51inter3), .O(gate51inter10));
  nor2  gate368(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate369(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate370(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );

  xor2  gate441(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate442(.a(gate53inter0), .b(s_40), .O(gate53inter1));
  and2  gate443(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate444(.a(s_40), .O(gate53inter3));
  inv1  gate445(.a(s_41), .O(gate53inter4));
  nand2 gate446(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate447(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate448(.a(N203), .O(gate53inter7));
  inv1  gate449(.a(N165), .O(gate53inter8));
  nand2 gate450(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate451(.a(s_41), .b(gate53inter3), .O(gate53inter10));
  nor2  gate452(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate453(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate454(.a(gate53inter12), .b(gate53inter1), .O(N233));

  xor2  gate385(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate386(.a(gate54inter0), .b(s_32), .O(gate54inter1));
  and2  gate387(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate388(.a(s_32), .O(gate54inter3));
  inv1  gate389(.a(s_33), .O(gate54inter4));
  nand2 gate390(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate391(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate392(.a(N203), .O(gate54inter7));
  inv1  gate393(.a(N168), .O(gate54inter8));
  nand2 gate394(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate395(.a(s_33), .b(gate54inter3), .O(gate54inter10));
  nor2  gate396(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate397(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate398(.a(gate54inter12), .b(gate54inter1), .O(N236));
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate329(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate330(.a(gate57inter0), .b(s_24), .O(gate57inter1));
  and2  gate331(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate332(.a(s_24), .O(gate57inter3));
  inv1  gate333(.a(s_25), .O(gate57inter4));
  nand2 gate334(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate335(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate336(.a(N203), .O(gate57inter7));
  inv1  gate337(.a(N174), .O(gate57inter8));
  nand2 gate338(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate339(.a(s_25), .b(gate57inter3), .O(gate57inter10));
  nor2  gate340(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate341(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate342(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate301(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate302(.a(gate59inter0), .b(s_20), .O(gate59inter1));
  and2  gate303(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate304(.a(s_20), .O(gate59inter3));
  inv1  gate305(.a(s_21), .O(gate59inter4));
  nand2 gate306(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate307(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate308(.a(N203), .O(gate59inter7));
  inv1  gate309(.a(N177), .O(gate59inter8));
  nand2 gate310(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate311(.a(s_21), .b(gate59inter3), .O(gate59inter10));
  nor2  gate312(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate313(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate314(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );

  xor2  gate273(.a(N180), .b(N203), .O(gate61inter0));
  nand2 gate274(.a(gate61inter0), .b(s_16), .O(gate61inter1));
  and2  gate275(.a(N180), .b(N203), .O(gate61inter2));
  inv1  gate276(.a(s_16), .O(gate61inter3));
  inv1  gate277(.a(s_17), .O(gate61inter4));
  nand2 gate278(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate279(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate280(.a(N203), .O(gate61inter7));
  inv1  gate281(.a(N180), .O(gate61inter8));
  nand2 gate282(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate283(.a(s_17), .b(gate61inter3), .O(gate61inter10));
  nor2  gate284(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate285(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate286(.a(gate61inter12), .b(gate61inter1), .O(N251));

  xor2  gate511(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate512(.a(gate62inter0), .b(s_50), .O(gate62inter1));
  and2  gate513(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate514(.a(s_50), .O(gate62inter3));
  inv1  gate515(.a(s_51), .O(gate62inter4));
  nand2 gate516(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate517(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate518(.a(N213), .O(gate62inter7));
  inv1  gate519(.a(N37), .O(gate62inter8));
  nand2 gate520(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate521(.a(s_51), .b(gate62inter3), .O(gate62inter10));
  nor2  gate522(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate523(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate524(.a(gate62inter12), .b(gate62inter1), .O(N254));

  xor2  gate203(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate204(.a(gate63inter0), .b(s_6), .O(gate63inter1));
  and2  gate205(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate206(.a(s_6), .O(gate63inter3));
  inv1  gate207(.a(s_7), .O(gate63inter4));
  nand2 gate208(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate209(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate210(.a(N213), .O(gate63inter7));
  inv1  gate211(.a(N50), .O(gate63inter8));
  nand2 gate212(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate213(.a(s_7), .b(gate63inter3), .O(gate63inter10));
  nor2  gate214(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate215(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate216(.a(gate63inter12), .b(gate63inter1), .O(N255));
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate609(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate610(.a(gate65inter0), .b(s_64), .O(gate65inter1));
  and2  gate611(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate612(.a(s_64), .O(gate65inter3));
  inv1  gate613(.a(s_65), .O(gate65inter4));
  nand2 gate614(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate615(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate616(.a(N213), .O(gate65inter7));
  inv1  gate617(.a(N76), .O(gate65inter8));
  nand2 gate618(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate619(.a(s_65), .b(gate65inter3), .O(gate65inter10));
  nor2  gate620(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate621(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate622(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );

  xor2  gate371(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate372(.a(gate69inter0), .b(s_30), .O(gate69inter1));
  and2  gate373(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate374(.a(s_30), .O(gate69inter3));
  inv1  gate375(.a(s_31), .O(gate69inter4));
  nand2 gate376(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate377(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate378(.a(N224), .O(gate69inter7));
  inv1  gate379(.a(N158), .O(gate69inter8));
  nand2 gate380(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate381(.a(s_31), .b(gate69inter3), .O(gate69inter10));
  nor2  gate382(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate383(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate384(.a(gate69inter12), .b(gate69inter1), .O(N263));

  xor2  gate399(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate400(.a(gate70inter0), .b(s_34), .O(gate70inter1));
  and2  gate401(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate402(.a(s_34), .O(gate70inter3));
  inv1  gate403(.a(s_35), .O(gate70inter4));
  nand2 gate404(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate405(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate406(.a(N227), .O(gate70inter7));
  inv1  gate407(.a(N183), .O(gate70inter8));
  nand2 gate408(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate409(.a(s_35), .b(gate70inter3), .O(gate70inter10));
  nor2  gate410(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate411(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate412(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate483(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate484(.a(gate72inter0), .b(s_46), .O(gate72inter1));
  and2  gate485(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate486(.a(s_46), .O(gate72inter3));
  inv1  gate487(.a(s_47), .O(gate72inter4));
  nand2 gate488(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate489(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate490(.a(N233), .O(gate72inter7));
  inv1  gate491(.a(N187), .O(gate72inter8));
  nand2 gate492(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate493(.a(s_47), .b(gate72inter3), .O(gate72inter10));
  nor2  gate494(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate495(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate496(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );

  xor2  gate175(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate176(.a(gate74inter0), .b(s_2), .O(gate74inter1));
  and2  gate177(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate178(.a(s_2), .O(gate74inter3));
  inv1  gate179(.a(s_3), .O(gate74inter4));
  nand2 gate180(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate181(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate182(.a(N239), .O(gate74inter7));
  inv1  gate183(.a(N191), .O(gate74inter8));
  nand2 gate184(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate185(.a(s_3), .b(gate74inter3), .O(gate74inter10));
  nor2  gate186(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate187(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate188(.a(gate74inter12), .b(gate74inter1), .O(N276));

  xor2  gate553(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate554(.a(gate75inter0), .b(s_56), .O(gate75inter1));
  and2  gate555(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate556(.a(s_56), .O(gate75inter3));
  inv1  gate557(.a(s_57), .O(gate75inter4));
  nand2 gate558(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate559(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate560(.a(N243), .O(gate75inter7));
  inv1  gate561(.a(N193), .O(gate75inter8));
  nand2 gate562(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate563(.a(s_57), .b(gate75inter3), .O(gate75inter10));
  nor2  gate564(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate565(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate566(.a(gate75inter12), .b(gate75inter1), .O(N279));

  xor2  gate343(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate344(.a(gate76inter0), .b(s_26), .O(gate76inter1));
  and2  gate345(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate346(.a(s_26), .O(gate76inter3));
  inv1  gate347(.a(s_27), .O(gate76inter4));
  nand2 gate348(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate349(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate350(.a(N247), .O(gate76inter7));
  inv1  gate351(.a(N195), .O(gate76inter8));
  nand2 gate352(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate353(.a(s_27), .b(gate76inter3), .O(gate76inter10));
  nor2  gate354(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate355(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate356(.a(gate76inter12), .b(gate76inter1), .O(N282));
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );

  xor2  gate525(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate526(.a(gate101inter0), .b(s_52), .O(gate101inter1));
  and2  gate527(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate528(.a(s_52), .O(gate101inter3));
  inv1  gate529(.a(s_53), .O(gate101inter4));
  nand2 gate530(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate531(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate532(.a(N309), .O(gate101inter7));
  inv1  gate533(.a(N267), .O(gate101inter8));
  nand2 gate534(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate535(.a(s_53), .b(gate101inter3), .O(gate101inter10));
  nor2  gate536(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate537(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate538(.a(gate101inter12), .b(gate101inter1), .O(N332));

  xor2  gate287(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate288(.a(gate102inter0), .b(s_18), .O(gate102inter1));
  and2  gate289(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate290(.a(s_18), .O(gate102inter3));
  inv1  gate291(.a(s_19), .O(gate102inter4));
  nand2 gate292(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate293(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate294(.a(N309), .O(gate102inter7));
  inv1  gate295(.a(N270), .O(gate102inter8));
  nand2 gate296(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate297(.a(s_19), .b(gate102inter3), .O(gate102inter10));
  nor2  gate298(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate299(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate300(.a(gate102inter12), .b(gate102inter1), .O(N333));

  xor2  gate567(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate568(.a(gate103inter0), .b(s_58), .O(gate103inter1));
  and2  gate569(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate570(.a(s_58), .O(gate103inter3));
  inv1  gate571(.a(s_59), .O(gate103inter4));
  nand2 gate572(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate573(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate574(.a(N8), .O(gate103inter7));
  inv1  gate575(.a(N319), .O(gate103inter8));
  nand2 gate576(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate577(.a(s_59), .b(gate103inter3), .O(gate103inter10));
  nor2  gate578(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate579(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate580(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );

  xor2  gate245(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate246(.a(gate106inter0), .b(s_12), .O(gate106inter1));
  and2  gate247(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate248(.a(s_12), .O(gate106inter3));
  inv1  gate249(.a(s_13), .O(gate106inter4));
  nand2 gate250(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate251(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate252(.a(N309), .O(gate106inter7));
  inv1  gate253(.a(N276), .O(gate106inter8));
  nand2 gate254(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate255(.a(s_13), .b(gate106inter3), .O(gate106inter10));
  nor2  gate256(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate257(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate258(.a(gate106inter12), .b(gate106inter1), .O(N337));

  xor2  gate469(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate470(.a(gate107inter0), .b(s_44), .O(gate107inter1));
  and2  gate471(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate472(.a(s_44), .O(gate107inter3));
  inv1  gate473(.a(s_45), .O(gate107inter4));
  nand2 gate474(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate475(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate476(.a(N319), .O(gate107inter7));
  inv1  gate477(.a(N34), .O(gate107inter8));
  nand2 gate478(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate479(.a(s_45), .b(gate107inter3), .O(gate107inter10));
  nor2  gate480(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate481(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate482(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );

  xor2  gate497(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate498(.a(gate109inter0), .b(s_48), .O(gate109inter1));
  and2  gate499(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate500(.a(s_48), .O(gate109inter3));
  inv1  gate501(.a(s_49), .O(gate109inter4));
  nand2 gate502(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate503(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate504(.a(N319), .O(gate109inter7));
  inv1  gate505(.a(N47), .O(gate109inter8));
  nand2 gate506(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate507(.a(s_49), .b(gate109inter3), .O(gate109inter10));
  nor2  gate508(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate509(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate510(.a(gate109inter12), .b(gate109inter1), .O(N340));
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate259(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate260(.a(gate113inter0), .b(s_14), .O(gate113inter1));
  and2  gate261(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate262(.a(s_14), .O(gate113inter3));
  inv1  gate263(.a(s_15), .O(gate113inter4));
  nand2 gate264(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate265(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate266(.a(N319), .O(gate113inter7));
  inv1  gate267(.a(N73), .O(gate113inter8));
  nand2 gate268(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate269(.a(s_15), .b(gate113inter3), .O(gate113inter10));
  nor2  gate270(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate271(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate272(.a(gate113inter12), .b(gate113inter1), .O(N344));

  xor2  gate161(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate162(.a(gate114inter0), .b(s_0), .O(gate114inter1));
  and2  gate163(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate164(.a(s_0), .O(gate114inter3));
  inv1  gate165(.a(s_1), .O(gate114inter4));
  nand2 gate166(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate167(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate168(.a(N319), .O(gate114inter7));
  inv1  gate169(.a(N86), .O(gate114inter8));
  nand2 gate170(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate171(.a(s_1), .b(gate114inter3), .O(gate114inter10));
  nor2  gate172(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate173(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate174(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate217(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate218(.a(gate120inter0), .b(s_8), .O(gate120inter1));
  and2  gate219(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate220(.a(s_8), .O(gate120inter3));
  inv1  gate221(.a(s_9), .O(gate120inter4));
  nand2 gate222(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate223(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate224(.a(N333), .O(gate120inter7));
  inv1  gate225(.a(N303), .O(gate120inter8));
  nand2 gate226(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate227(.a(s_9), .b(gate120inter3), .O(gate120inter10));
  nor2  gate228(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate229(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate230(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate623(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate624(.a(gate129inter0), .b(s_66), .O(gate129inter1));
  and2  gate625(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate626(.a(s_66), .O(gate129inter3));
  inv1  gate627(.a(s_67), .O(gate129inter4));
  nand2 gate628(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate629(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate630(.a(N14), .O(gate129inter7));
  inv1  gate631(.a(N360), .O(gate129inter8));
  nand2 gate632(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate633(.a(s_67), .b(gate129inter3), .O(gate129inter10));
  nor2  gate634(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate635(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate636(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate637(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate638(.a(gate132inter0), .b(s_68), .O(gate132inter1));
  and2  gate639(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate640(.a(s_68), .O(gate132inter3));
  inv1  gate641(.a(s_69), .O(gate132inter4));
  nand2 gate642(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate643(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate644(.a(N360), .O(gate132inter7));
  inv1  gate645(.a(N53), .O(gate132inter8));
  nand2 gate646(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate647(.a(s_69), .b(gate132inter3), .O(gate132inter10));
  nor2  gate648(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate649(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate650(.a(gate132inter12), .b(gate132inter1), .O(N374));

  xor2  gate231(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate232(.a(gate133inter0), .b(s_10), .O(gate133inter1));
  and2  gate233(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate234(.a(s_10), .O(gate133inter3));
  inv1  gate235(.a(s_11), .O(gate133inter4));
  nand2 gate236(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate237(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate238(.a(N360), .O(gate133inter7));
  inv1  gate239(.a(N66), .O(gate133inter8));
  nand2 gate240(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate241(.a(s_11), .b(gate133inter3), .O(gate133inter10));
  nor2  gate242(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate243(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate244(.a(gate133inter12), .b(gate133inter1), .O(N375));
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate651(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate652(.a(gate136inter0), .b(s_70), .O(gate136inter1));
  and2  gate653(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate654(.a(s_70), .O(gate136inter3));
  inv1  gate655(.a(s_71), .O(gate136inter4));
  nand2 gate656(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate657(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate658(.a(N360), .O(gate136inter7));
  inv1  gate659(.a(N105), .O(gate136inter8));
  nand2 gate660(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate661(.a(s_71), .b(gate136inter3), .O(gate136inter10));
  nor2  gate662(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate663(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate664(.a(gate136inter12), .b(gate136inter1), .O(N378));

  xor2  gate539(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate540(.a(gate137inter0), .b(s_54), .O(gate137inter1));
  and2  gate541(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate542(.a(s_54), .O(gate137inter3));
  inv1  gate543(.a(s_55), .O(gate137inter4));
  nand2 gate544(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate545(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate546(.a(N360), .O(gate137inter7));
  inv1  gate547(.a(N115), .O(gate137inter8));
  nand2 gate548(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate549(.a(s_55), .b(gate137inter3), .O(gate137inter10));
  nor2  gate550(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate551(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate552(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule