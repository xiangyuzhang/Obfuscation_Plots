module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );

  xor2  gate595(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate596(.a(gate20inter0), .b(s_62), .O(gate20inter1));
  and2  gate597(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate598(.a(s_62), .O(gate20inter3));
  inv1  gate599(.a(s_63), .O(gate20inter4));
  nand2 gate600(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate601(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate602(.a(N8), .O(gate20inter7));
  inv1  gate603(.a(N119), .O(gate20inter8));
  nand2 gate604(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate605(.a(s_63), .b(gate20inter3), .O(gate20inter10));
  nor2  gate606(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate607(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate608(.a(gate20inter12), .b(gate20inter1), .O(N157));

  xor2  gate315(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate316(.a(gate21inter0), .b(s_22), .O(gate21inter1));
  and2  gate317(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate318(.a(s_22), .O(gate21inter3));
  inv1  gate319(.a(s_23), .O(gate21inter4));
  nand2 gate320(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate321(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate322(.a(N14), .O(gate21inter7));
  inv1  gate323(.a(N119), .O(gate21inter8));
  nand2 gate324(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate325(.a(s_23), .b(gate21inter3), .O(gate21inter10));
  nor2  gate326(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate327(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate328(.a(gate21inter12), .b(gate21inter1), .O(N158));
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate231(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate232(.a(gate24inter0), .b(s_10), .O(gate24inter1));
  and2  gate233(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate234(.a(s_10), .O(gate24inter3));
  inv1  gate235(.a(s_11), .O(gate24inter4));
  nand2 gate236(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate237(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate238(.a(N130), .O(gate24inter7));
  inv1  gate239(.a(N43), .O(gate24inter8));
  nand2 gate240(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate241(.a(s_11), .b(gate24inter3), .O(gate24inter10));
  nor2  gate242(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate243(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate244(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate245(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate246(.a(gate27inter0), .b(s_12), .O(gate27inter1));
  and2  gate247(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate248(.a(s_12), .O(gate27inter3));
  inv1  gate249(.a(s_13), .O(gate27inter4));
  nand2 gate250(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate251(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate252(.a(N142), .O(gate27inter7));
  inv1  gate253(.a(N82), .O(gate27inter8));
  nand2 gate254(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate255(.a(s_13), .b(gate27inter3), .O(gate27inter10));
  nor2  gate256(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate257(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate258(.a(gate27inter12), .b(gate27inter1), .O(N174));

  xor2  gate483(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate484(.a(gate28inter0), .b(s_46), .O(gate28inter1));
  and2  gate485(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate486(.a(s_46), .O(gate28inter3));
  inv1  gate487(.a(s_47), .O(gate28inter4));
  nand2 gate488(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate489(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate490(.a(N146), .O(gate28inter7));
  inv1  gate491(.a(N95), .O(gate28inter8));
  nand2 gate492(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate493(.a(s_47), .b(gate28inter3), .O(gate28inter10));
  nor2  gate494(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate495(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate496(.a(gate28inter12), .b(gate28inter1), .O(N177));

  xor2  gate553(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate554(.a(gate29inter0), .b(s_56), .O(gate29inter1));
  and2  gate555(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate556(.a(s_56), .O(gate29inter3));
  inv1  gate557(.a(s_57), .O(gate29inter4));
  nand2 gate558(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate559(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate560(.a(N150), .O(gate29inter7));
  inv1  gate561(.a(N108), .O(gate29inter8));
  nand2 gate562(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate563(.a(s_57), .b(gate29inter3), .O(gate29inter10));
  nor2  gate564(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate565(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate566(.a(gate29inter12), .b(gate29inter1), .O(N180));

  xor2  gate791(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate792(.a(gate30inter0), .b(s_90), .O(gate30inter1));
  and2  gate793(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate794(.a(s_90), .O(gate30inter3));
  inv1  gate795(.a(s_91), .O(gate30inter4));
  nand2 gate796(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate797(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate798(.a(N21), .O(gate30inter7));
  inv1  gate799(.a(N123), .O(gate30inter8));
  nand2 gate800(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate801(.a(s_91), .b(gate30inter3), .O(gate30inter10));
  nor2  gate802(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate803(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate804(.a(gate30inter12), .b(gate30inter1), .O(N183));
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate497(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate498(.a(gate34inter0), .b(s_48), .O(gate34inter1));
  and2  gate499(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate500(.a(s_48), .O(gate34inter3));
  inv1  gate501(.a(s_49), .O(gate34inter4));
  nand2 gate502(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate503(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate504(.a(N47), .O(gate34inter7));
  inv1  gate505(.a(N131), .O(gate34inter8));
  nand2 gate506(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate507(.a(s_49), .b(gate34inter3), .O(gate34inter10));
  nor2  gate508(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate509(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate510(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate287(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate288(.a(gate35inter0), .b(s_18), .O(gate35inter1));
  and2  gate289(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate290(.a(s_18), .O(gate35inter3));
  inv1  gate291(.a(s_19), .O(gate35inter4));
  nand2 gate292(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate293(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate294(.a(N53), .O(gate35inter7));
  inv1  gate295(.a(N131), .O(gate35inter8));
  nand2 gate296(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate297(.a(s_19), .b(gate35inter3), .O(gate35inter10));
  nor2  gate298(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate299(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate300(.a(gate35inter12), .b(gate35inter1), .O(N188));

  xor2  gate749(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate750(.a(gate36inter0), .b(s_84), .O(gate36inter1));
  and2  gate751(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate752(.a(s_84), .O(gate36inter3));
  inv1  gate753(.a(s_85), .O(gate36inter4));
  nand2 gate754(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate755(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate756(.a(N60), .O(gate36inter7));
  inv1  gate757(.a(N135), .O(gate36inter8));
  nand2 gate758(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate759(.a(s_85), .b(gate36inter3), .O(gate36inter10));
  nor2  gate760(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate761(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate762(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate175(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate176(.a(gate40inter0), .b(s_2), .O(gate40inter1));
  and2  gate177(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate178(.a(s_2), .O(gate40inter3));
  inv1  gate179(.a(s_3), .O(gate40inter4));
  nand2 gate180(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate181(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate182(.a(N86), .O(gate40inter7));
  inv1  gate183(.a(N143), .O(gate40inter8));
  nand2 gate184(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate185(.a(s_3), .b(gate40inter3), .O(gate40inter10));
  nor2  gate186(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate187(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate188(.a(gate40inter12), .b(gate40inter1), .O(N193));

  xor2  gate525(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate526(.a(gate41inter0), .b(s_52), .O(gate41inter1));
  and2  gate527(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate528(.a(s_52), .O(gate41inter3));
  inv1  gate529(.a(s_53), .O(gate41inter4));
  nand2 gate530(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate531(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate532(.a(N92), .O(gate41inter7));
  inv1  gate533(.a(N143), .O(gate41inter8));
  nand2 gate534(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate535(.a(s_53), .b(gate41inter3), .O(gate41inter10));
  nor2  gate536(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate537(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate538(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate637(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate638(.a(gate43inter0), .b(s_68), .O(gate43inter1));
  and2  gate639(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate640(.a(s_68), .O(gate43inter3));
  inv1  gate641(.a(s_69), .O(gate43inter4));
  nand2 gate642(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate643(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate644(.a(N105), .O(gate43inter7));
  inv1  gate645(.a(N147), .O(gate43inter8));
  nand2 gate646(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate647(.a(s_69), .b(gate43inter3), .O(gate43inter10));
  nor2  gate648(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate649(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate650(.a(gate43inter12), .b(gate43inter1), .O(N196));

  xor2  gate217(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate218(.a(gate44inter0), .b(s_8), .O(gate44inter1));
  and2  gate219(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate220(.a(s_8), .O(gate44inter3));
  inv1  gate221(.a(s_9), .O(gate44inter4));
  nand2 gate222(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate223(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate224(.a(N112), .O(gate44inter7));
  inv1  gate225(.a(N151), .O(gate44inter8));
  nand2 gate226(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate227(.a(s_9), .b(gate44inter3), .O(gate44inter10));
  nor2  gate228(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate229(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate230(.a(gate44inter12), .b(gate44inter1), .O(N197));
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate763(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate764(.a(gate50inter0), .b(s_86), .O(gate50inter1));
  and2  gate765(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate766(.a(s_86), .O(gate50inter3));
  inv1  gate767(.a(s_87), .O(gate50inter4));
  nand2 gate768(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate769(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate770(.a(N203), .O(gate50inter7));
  inv1  gate771(.a(N154), .O(gate50inter8));
  nand2 gate772(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate773(.a(s_87), .b(gate50inter3), .O(gate50inter10));
  nor2  gate774(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate775(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate776(.a(gate50inter12), .b(gate50inter1), .O(N224));
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );

  xor2  gate413(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate414(.a(gate55inter0), .b(s_36), .O(gate55inter1));
  and2  gate415(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate416(.a(s_36), .O(gate55inter3));
  inv1  gate417(.a(s_37), .O(gate55inter4));
  nand2 gate418(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate419(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate420(.a(N203), .O(gate55inter7));
  inv1  gate421(.a(N171), .O(gate55inter8));
  nand2 gate422(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate423(.a(s_37), .b(gate55inter3), .O(gate55inter10));
  nor2  gate424(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate425(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate426(.a(gate55inter12), .b(gate55inter1), .O(N239));

  xor2  gate357(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate358(.a(gate56inter0), .b(s_28), .O(gate56inter1));
  and2  gate359(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate360(.a(s_28), .O(gate56inter3));
  inv1  gate361(.a(s_29), .O(gate56inter4));
  nand2 gate362(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate363(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate364(.a(N1), .O(gate56inter7));
  inv1  gate365(.a(N213), .O(gate56inter8));
  nand2 gate366(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate367(.a(s_29), .b(gate56inter3), .O(gate56inter10));
  nor2  gate368(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate369(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate370(.a(gate56inter12), .b(gate56inter1), .O(N242));

  xor2  gate427(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate428(.a(gate57inter0), .b(s_38), .O(gate57inter1));
  and2  gate429(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate430(.a(s_38), .O(gate57inter3));
  inv1  gate431(.a(s_39), .O(gate57inter4));
  nand2 gate432(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate433(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate434(.a(N203), .O(gate57inter7));
  inv1  gate435(.a(N174), .O(gate57inter8));
  nand2 gate436(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate437(.a(s_39), .b(gate57inter3), .O(gate57inter10));
  nor2  gate438(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate439(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate440(.a(gate57inter12), .b(gate57inter1), .O(N243));

  xor2  gate329(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate330(.a(gate58inter0), .b(s_24), .O(gate58inter1));
  and2  gate331(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate332(.a(s_24), .O(gate58inter3));
  inv1  gate333(.a(s_25), .O(gate58inter4));
  nand2 gate334(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate335(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate336(.a(N213), .O(gate58inter7));
  inv1  gate337(.a(N11), .O(gate58inter8));
  nand2 gate338(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate339(.a(s_25), .b(gate58inter3), .O(gate58inter10));
  nor2  gate340(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate341(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate342(.a(gate58inter12), .b(gate58inter1), .O(N246));

  xor2  gate189(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate190(.a(gate59inter0), .b(s_4), .O(gate59inter1));
  and2  gate191(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate192(.a(s_4), .O(gate59inter3));
  inv1  gate193(.a(s_5), .O(gate59inter4));
  nand2 gate194(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate195(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate196(.a(N203), .O(gate59inter7));
  inv1  gate197(.a(N177), .O(gate59inter8));
  nand2 gate198(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate199(.a(s_5), .b(gate59inter3), .O(gate59inter10));
  nor2  gate200(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate201(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate202(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );

  xor2  gate399(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate400(.a(gate64inter0), .b(s_34), .O(gate64inter1));
  and2  gate401(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate402(.a(s_34), .O(gate64inter3));
  inv1  gate403(.a(s_35), .O(gate64inter4));
  nand2 gate404(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate405(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate406(.a(N213), .O(gate64inter7));
  inv1  gate407(.a(N63), .O(gate64inter8));
  nand2 gate408(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate409(.a(s_35), .b(gate64inter3), .O(gate64inter10));
  nor2  gate410(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate411(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate412(.a(gate64inter12), .b(gate64inter1), .O(N256));
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate343(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate344(.a(gate68inter0), .b(s_26), .O(gate68inter1));
  and2  gate345(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate346(.a(s_26), .O(gate68inter3));
  inv1  gate347(.a(s_27), .O(gate68inter4));
  nand2 gate348(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate349(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate350(.a(N224), .O(gate68inter7));
  inv1  gate351(.a(N157), .O(gate68inter8));
  nand2 gate352(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate353(.a(s_27), .b(gate68inter3), .O(gate68inter10));
  nor2  gate354(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate355(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate356(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate777(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate778(.a(gate70inter0), .b(s_88), .O(gate70inter1));
  and2  gate779(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate780(.a(s_88), .O(gate70inter3));
  inv1  gate781(.a(s_89), .O(gate70inter4));
  nand2 gate782(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate783(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate784(.a(N227), .O(gate70inter7));
  inv1  gate785(.a(N183), .O(gate70inter8));
  nand2 gate786(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate787(.a(s_89), .b(gate70inter3), .O(gate70inter10));
  nor2  gate788(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate789(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate790(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate567(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate568(.a(gate73inter0), .b(s_58), .O(gate73inter1));
  and2  gate569(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate570(.a(s_58), .O(gate73inter3));
  inv1  gate571(.a(s_59), .O(gate73inter4));
  nand2 gate572(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate573(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate574(.a(N236), .O(gate73inter7));
  inv1  gate575(.a(N189), .O(gate73inter8));
  nand2 gate576(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate577(.a(s_59), .b(gate73inter3), .O(gate73inter10));
  nor2  gate578(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate579(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate580(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate581(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate582(.a(gate77inter0), .b(s_60), .O(gate77inter1));
  and2  gate583(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate584(.a(s_60), .O(gate77inter3));
  inv1  gate585(.a(s_61), .O(gate77inter4));
  nand2 gate586(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate587(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate588(.a(N251), .O(gate77inter7));
  inv1  gate589(.a(N197), .O(gate77inter8));
  nand2 gate590(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate591(.a(s_61), .b(gate77inter3), .O(gate77inter10));
  nor2  gate592(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate593(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate594(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate371(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate372(.a(gate80inter0), .b(s_30), .O(gate80inter1));
  and2  gate373(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate374(.a(s_30), .O(gate80inter3));
  inv1  gate375(.a(s_31), .O(gate80inter4));
  nand2 gate376(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate377(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate378(.a(N233), .O(gate80inter7));
  inv1  gate379(.a(N188), .O(gate80inter8));
  nand2 gate380(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate381(.a(s_31), .b(gate80inter3), .O(gate80inter10));
  nor2  gate382(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate383(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate384(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate259(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate260(.a(gate83inter0), .b(s_14), .O(gate83inter1));
  and2  gate261(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate262(.a(s_14), .O(gate83inter3));
  inv1  gate263(.a(s_15), .O(gate83inter4));
  nand2 gate264(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate265(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate266(.a(N243), .O(gate83inter7));
  inv1  gate267(.a(N194), .O(gate83inter8));
  nand2 gate268(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate269(.a(s_15), .b(gate83inter3), .O(gate83inter10));
  nor2  gate270(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate271(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate272(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );

  xor2  gate273(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate274(.a(gate102inter0), .b(s_16), .O(gate102inter1));
  and2  gate275(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate276(.a(s_16), .O(gate102inter3));
  inv1  gate277(.a(s_17), .O(gate102inter4));
  nand2 gate278(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate279(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate280(.a(N309), .O(gate102inter7));
  inv1  gate281(.a(N270), .O(gate102inter8));
  nand2 gate282(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate283(.a(s_17), .b(gate102inter3), .O(gate102inter10));
  nor2  gate284(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate285(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate286(.a(gate102inter12), .b(gate102inter1), .O(N333));

  xor2  gate441(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate442(.a(gate103inter0), .b(s_40), .O(gate103inter1));
  and2  gate443(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate444(.a(s_40), .O(gate103inter3));
  inv1  gate445(.a(s_41), .O(gate103inter4));
  nand2 gate446(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate447(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate448(.a(N8), .O(gate103inter7));
  inv1  gate449(.a(N319), .O(gate103inter8));
  nand2 gate450(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate451(.a(s_41), .b(gate103inter3), .O(gate103inter10));
  nor2  gate452(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate453(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate454(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate455(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate456(.a(gate105inter0), .b(s_42), .O(gate105inter1));
  and2  gate457(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate458(.a(s_42), .O(gate105inter3));
  inv1  gate459(.a(s_43), .O(gate105inter4));
  nand2 gate460(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate461(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate462(.a(N319), .O(gate105inter7));
  inv1  gate463(.a(N21), .O(gate105inter8));
  nand2 gate464(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate465(.a(s_43), .b(gate105inter3), .O(gate105inter10));
  nor2  gate466(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate467(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate468(.a(gate105inter12), .b(gate105inter1), .O(N336));

  xor2  gate735(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate736(.a(gate106inter0), .b(s_82), .O(gate106inter1));
  and2  gate737(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate738(.a(s_82), .O(gate106inter3));
  inv1  gate739(.a(s_83), .O(gate106inter4));
  nand2 gate740(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate741(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate742(.a(N309), .O(gate106inter7));
  inv1  gate743(.a(N276), .O(gate106inter8));
  nand2 gate744(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate745(.a(s_83), .b(gate106inter3), .O(gate106inter10));
  nor2  gate746(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate747(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate748(.a(gate106inter12), .b(gate106inter1), .O(N337));

  xor2  gate693(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate694(.a(gate107inter0), .b(s_76), .O(gate107inter1));
  and2  gate695(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate696(.a(s_76), .O(gate107inter3));
  inv1  gate697(.a(s_77), .O(gate107inter4));
  nand2 gate698(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate699(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate700(.a(N319), .O(gate107inter7));
  inv1  gate701(.a(N34), .O(gate107inter8));
  nand2 gate702(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate703(.a(s_77), .b(gate107inter3), .O(gate107inter10));
  nor2  gate704(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate705(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate706(.a(gate107inter12), .b(gate107inter1), .O(N338));

  xor2  gate161(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate162(.a(gate108inter0), .b(s_0), .O(gate108inter1));
  and2  gate163(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate164(.a(s_0), .O(gate108inter3));
  inv1  gate165(.a(s_1), .O(gate108inter4));
  nand2 gate166(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate167(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate168(.a(N309), .O(gate108inter7));
  inv1  gate169(.a(N279), .O(gate108inter8));
  nand2 gate170(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate171(.a(s_1), .b(gate108inter3), .O(gate108inter10));
  nor2  gate172(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate173(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate174(.a(gate108inter12), .b(gate108inter1), .O(N339));

  xor2  gate679(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate680(.a(gate109inter0), .b(s_74), .O(gate109inter1));
  and2  gate681(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate682(.a(s_74), .O(gate109inter3));
  inv1  gate683(.a(s_75), .O(gate109inter4));
  nand2 gate684(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate685(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate686(.a(N319), .O(gate109inter7));
  inv1  gate687(.a(N47), .O(gate109inter8));
  nand2 gate688(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate689(.a(s_75), .b(gate109inter3), .O(gate109inter10));
  nor2  gate690(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate691(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate692(.a(gate109inter12), .b(gate109inter1), .O(N340));
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate721(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate722(.a(gate111inter0), .b(s_80), .O(gate111inter1));
  and2  gate723(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate724(.a(s_80), .O(gate111inter3));
  inv1  gate725(.a(s_81), .O(gate111inter4));
  nand2 gate726(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate727(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate728(.a(N319), .O(gate111inter7));
  inv1  gate729(.a(N60), .O(gate111inter8));
  nand2 gate730(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate731(.a(s_81), .b(gate111inter3), .O(gate111inter10));
  nor2  gate732(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate733(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate734(.a(gate111inter12), .b(gate111inter1), .O(N342));

  xor2  gate609(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate610(.a(gate112inter0), .b(s_64), .O(gate112inter1));
  and2  gate611(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate612(.a(s_64), .O(gate112inter3));
  inv1  gate613(.a(s_65), .O(gate112inter4));
  nand2 gate614(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate615(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate616(.a(N309), .O(gate112inter7));
  inv1  gate617(.a(N285), .O(gate112inter8));
  nand2 gate618(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate619(.a(s_65), .b(gate112inter3), .O(gate112inter10));
  nor2  gate620(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate621(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate622(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );

  xor2  gate707(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate708(.a(gate114inter0), .b(s_78), .O(gate114inter1));
  and2  gate709(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate710(.a(s_78), .O(gate114inter3));
  inv1  gate711(.a(s_79), .O(gate114inter4));
  nand2 gate712(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate713(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate714(.a(N319), .O(gate114inter7));
  inv1  gate715(.a(N86), .O(gate114inter8));
  nand2 gate716(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate717(.a(s_79), .b(gate114inter3), .O(gate114inter10));
  nor2  gate718(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate719(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate720(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );

  xor2  gate301(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate302(.a(gate117inter0), .b(s_20), .O(gate117inter1));
  and2  gate303(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate304(.a(s_20), .O(gate117inter3));
  inv1  gate305(.a(s_21), .O(gate117inter4));
  nand2 gate306(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate307(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate308(.a(N330), .O(gate117inter7));
  inv1  gate309(.a(N300), .O(gate117inter8));
  nand2 gate310(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate311(.a(s_21), .b(gate117inter3), .O(gate117inter10));
  nor2  gate312(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate313(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate314(.a(gate117inter12), .b(gate117inter1), .O(N348));

  xor2  gate665(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate666(.a(gate118inter0), .b(s_72), .O(gate118inter1));
  and2  gate667(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate668(.a(s_72), .O(gate118inter3));
  inv1  gate669(.a(s_73), .O(gate118inter4));
  nand2 gate670(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate671(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate672(.a(N331), .O(gate118inter7));
  inv1  gate673(.a(N301), .O(gate118inter8));
  nand2 gate674(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate675(.a(s_73), .b(gate118inter3), .O(gate118inter10));
  nor2  gate676(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate677(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate678(.a(gate118inter12), .b(gate118inter1), .O(N349));

  xor2  gate651(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate652(.a(gate119inter0), .b(s_70), .O(gate119inter1));
  and2  gate653(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate654(.a(s_70), .O(gate119inter3));
  inv1  gate655(.a(s_71), .O(gate119inter4));
  nand2 gate656(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate657(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate658(.a(N332), .O(gate119inter7));
  inv1  gate659(.a(N302), .O(gate119inter8));
  nand2 gate660(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate661(.a(s_71), .b(gate119inter3), .O(gate119inter10));
  nor2  gate662(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate663(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate664(.a(gate119inter12), .b(gate119inter1), .O(N350));

  xor2  gate511(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate512(.a(gate120inter0), .b(s_50), .O(gate120inter1));
  and2  gate513(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate514(.a(s_50), .O(gate120inter3));
  inv1  gate515(.a(s_51), .O(gate120inter4));
  nand2 gate516(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate517(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate518(.a(N333), .O(gate120inter7));
  inv1  gate519(.a(N303), .O(gate120inter8));
  nand2 gate520(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate521(.a(s_51), .b(gate120inter3), .O(gate120inter10));
  nor2  gate522(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate523(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate524(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );

  xor2  gate203(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate204(.a(gate122inter0), .b(s_6), .O(gate122inter1));
  and2  gate205(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate206(.a(s_6), .O(gate122inter3));
  inv1  gate207(.a(s_7), .O(gate122inter4));
  nand2 gate208(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate209(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate210(.a(N337), .O(gate122inter7));
  inv1  gate211(.a(N305), .O(gate122inter8));
  nand2 gate212(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate213(.a(s_7), .b(gate122inter3), .O(gate122inter10));
  nor2  gate214(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate215(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate216(.a(gate122inter12), .b(gate122inter1), .O(N353));
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate623(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate624(.a(gate129inter0), .b(s_66), .O(gate129inter1));
  and2  gate625(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate626(.a(s_66), .O(gate129inter3));
  inv1  gate627(.a(s_67), .O(gate129inter4));
  nand2 gate628(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate629(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate630(.a(N14), .O(gate129inter7));
  inv1  gate631(.a(N360), .O(gate129inter8));
  nand2 gate632(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate633(.a(s_67), .b(gate129inter3), .O(gate129inter10));
  nor2  gate634(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate635(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate636(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate469(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate470(.a(gate131inter0), .b(s_44), .O(gate131inter1));
  and2  gate471(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate472(.a(s_44), .O(gate131inter3));
  inv1  gate473(.a(s_45), .O(gate131inter4));
  nand2 gate474(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate475(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate476(.a(N360), .O(gate131inter7));
  inv1  gate477(.a(N40), .O(gate131inter8));
  nand2 gate478(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate479(.a(s_45), .b(gate131inter3), .O(gate131inter10));
  nor2  gate480(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate481(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate482(.a(gate131inter12), .b(gate131inter1), .O(N373));

  xor2  gate385(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate386(.a(gate132inter0), .b(s_32), .O(gate132inter1));
  and2  gate387(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate388(.a(s_32), .O(gate132inter3));
  inv1  gate389(.a(s_33), .O(gate132inter4));
  nand2 gate390(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate391(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate392(.a(N360), .O(gate132inter7));
  inv1  gate393(.a(N53), .O(gate132inter8));
  nand2 gate394(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate395(.a(s_33), .b(gate132inter3), .O(gate132inter10));
  nor2  gate396(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate397(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate398(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );

  xor2  gate539(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate540(.a(gate137inter0), .b(s_54), .O(gate137inter1));
  and2  gate541(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate542(.a(s_54), .O(gate137inter3));
  inv1  gate543(.a(s_55), .O(gate137inter4));
  nand2 gate544(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate545(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate546(.a(N360), .O(gate137inter7));
  inv1  gate547(.a(N115), .O(gate137inter8));
  nand2 gate548(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate549(.a(s_55), .b(gate137inter3), .O(gate137inter10));
  nor2  gate550(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate551(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate552(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule