module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate967(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate968(.a(gate20inter0), .b(s_60), .O(gate20inter1));
  and2  gate969(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate970(.a(s_60), .O(gate20inter3));
  inv1  gate971(.a(s_61), .O(gate20inter4));
  nand2 gate972(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate973(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate974(.a(G23), .O(gate20inter7));
  inv1  gate975(.a(G24), .O(gate20inter8));
  nand2 gate976(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate977(.a(s_61), .b(gate20inter3), .O(gate20inter10));
  nor2  gate978(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate979(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate980(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1079(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1080(.a(gate25inter0), .b(s_76), .O(gate25inter1));
  and2  gate1081(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1082(.a(s_76), .O(gate25inter3));
  inv1  gate1083(.a(s_77), .O(gate25inter4));
  nand2 gate1084(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1085(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1086(.a(G1), .O(gate25inter7));
  inv1  gate1087(.a(G5), .O(gate25inter8));
  nand2 gate1088(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1089(.a(s_77), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1090(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1091(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1092(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate841(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate842(.a(gate26inter0), .b(s_42), .O(gate26inter1));
  and2  gate843(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate844(.a(s_42), .O(gate26inter3));
  inv1  gate845(.a(s_43), .O(gate26inter4));
  nand2 gate846(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate847(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate848(.a(G9), .O(gate26inter7));
  inv1  gate849(.a(G13), .O(gate26inter8));
  nand2 gate850(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate851(.a(s_43), .b(gate26inter3), .O(gate26inter10));
  nor2  gate852(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate853(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate854(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate659(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate660(.a(gate29inter0), .b(s_16), .O(gate29inter1));
  and2  gate661(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate662(.a(s_16), .O(gate29inter3));
  inv1  gate663(.a(s_17), .O(gate29inter4));
  nand2 gate664(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate665(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate666(.a(G3), .O(gate29inter7));
  inv1  gate667(.a(G7), .O(gate29inter8));
  nand2 gate668(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate669(.a(s_17), .b(gate29inter3), .O(gate29inter10));
  nor2  gate670(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate671(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate672(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1009(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1010(.a(gate30inter0), .b(s_66), .O(gate30inter1));
  and2  gate1011(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1012(.a(s_66), .O(gate30inter3));
  inv1  gate1013(.a(s_67), .O(gate30inter4));
  nand2 gate1014(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1015(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1016(.a(G11), .O(gate30inter7));
  inv1  gate1017(.a(G15), .O(gate30inter8));
  nand2 gate1018(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1019(.a(s_67), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1020(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1021(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1022(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate813(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate814(.a(gate48inter0), .b(s_38), .O(gate48inter1));
  and2  gate815(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate816(.a(s_38), .O(gate48inter3));
  inv1  gate817(.a(s_39), .O(gate48inter4));
  nand2 gate818(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate819(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate820(.a(G8), .O(gate48inter7));
  inv1  gate821(.a(G275), .O(gate48inter8));
  nand2 gate822(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate823(.a(s_39), .b(gate48inter3), .O(gate48inter10));
  nor2  gate824(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate825(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate826(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1107(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1108(.a(gate54inter0), .b(s_80), .O(gate54inter1));
  and2  gate1109(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1110(.a(s_80), .O(gate54inter3));
  inv1  gate1111(.a(s_81), .O(gate54inter4));
  nand2 gate1112(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1113(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1114(.a(G14), .O(gate54inter7));
  inv1  gate1115(.a(G284), .O(gate54inter8));
  nand2 gate1116(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1117(.a(s_81), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1118(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1119(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1120(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate827(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate828(.a(gate66inter0), .b(s_40), .O(gate66inter1));
  and2  gate829(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate830(.a(s_40), .O(gate66inter3));
  inv1  gate831(.a(s_41), .O(gate66inter4));
  nand2 gate832(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate833(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate834(.a(G26), .O(gate66inter7));
  inv1  gate835(.a(G302), .O(gate66inter8));
  nand2 gate836(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate837(.a(s_41), .b(gate66inter3), .O(gate66inter10));
  nor2  gate838(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate839(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate840(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1037(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1038(.a(gate67inter0), .b(s_70), .O(gate67inter1));
  and2  gate1039(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1040(.a(s_70), .O(gate67inter3));
  inv1  gate1041(.a(s_71), .O(gate67inter4));
  nand2 gate1042(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1043(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1044(.a(G27), .O(gate67inter7));
  inv1  gate1045(.a(G305), .O(gate67inter8));
  nand2 gate1046(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1047(.a(s_71), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1048(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1049(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1050(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate673(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate674(.a(gate75inter0), .b(s_18), .O(gate75inter1));
  and2  gate675(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate676(.a(s_18), .O(gate75inter3));
  inv1  gate677(.a(s_19), .O(gate75inter4));
  nand2 gate678(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate679(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate680(.a(G9), .O(gate75inter7));
  inv1  gate681(.a(G317), .O(gate75inter8));
  nand2 gate682(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate683(.a(s_19), .b(gate75inter3), .O(gate75inter10));
  nor2  gate684(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate685(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate686(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1219(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1220(.a(gate76inter0), .b(s_96), .O(gate76inter1));
  and2  gate1221(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1222(.a(s_96), .O(gate76inter3));
  inv1  gate1223(.a(s_97), .O(gate76inter4));
  nand2 gate1224(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1225(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1226(.a(G13), .O(gate76inter7));
  inv1  gate1227(.a(G317), .O(gate76inter8));
  nand2 gate1228(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1229(.a(s_97), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1230(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1231(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1232(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate869(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate870(.a(gate78inter0), .b(s_46), .O(gate78inter1));
  and2  gate871(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate872(.a(s_46), .O(gate78inter3));
  inv1  gate873(.a(s_47), .O(gate78inter4));
  nand2 gate874(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate875(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate876(.a(G6), .O(gate78inter7));
  inv1  gate877(.a(G320), .O(gate78inter8));
  nand2 gate878(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate879(.a(s_47), .b(gate78inter3), .O(gate78inter10));
  nor2  gate880(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate881(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate882(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1065(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1066(.a(gate87inter0), .b(s_74), .O(gate87inter1));
  and2  gate1067(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1068(.a(s_74), .O(gate87inter3));
  inv1  gate1069(.a(s_75), .O(gate87inter4));
  nand2 gate1070(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1071(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1072(.a(G12), .O(gate87inter7));
  inv1  gate1073(.a(G335), .O(gate87inter8));
  nand2 gate1074(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1075(.a(s_75), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1076(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1077(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1078(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate771(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate772(.a(gate89inter0), .b(s_32), .O(gate89inter1));
  and2  gate773(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate774(.a(s_32), .O(gate89inter3));
  inv1  gate775(.a(s_33), .O(gate89inter4));
  nand2 gate776(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate777(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate778(.a(G17), .O(gate89inter7));
  inv1  gate779(.a(G338), .O(gate89inter8));
  nand2 gate780(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate781(.a(s_33), .b(gate89inter3), .O(gate89inter10));
  nor2  gate782(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate783(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate784(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate995(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate996(.a(gate96inter0), .b(s_64), .O(gate96inter1));
  and2  gate997(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate998(.a(s_64), .O(gate96inter3));
  inv1  gate999(.a(s_65), .O(gate96inter4));
  nand2 gate1000(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1001(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1002(.a(G30), .O(gate96inter7));
  inv1  gate1003(.a(G347), .O(gate96inter8));
  nand2 gate1004(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1005(.a(s_65), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1006(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1007(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1008(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate547(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate548(.a(gate116inter0), .b(s_0), .O(gate116inter1));
  and2  gate549(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate550(.a(s_0), .O(gate116inter3));
  inv1  gate551(.a(s_1), .O(gate116inter4));
  nand2 gate552(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate553(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate554(.a(G384), .O(gate116inter7));
  inv1  gate555(.a(G385), .O(gate116inter8));
  nand2 gate556(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate557(.a(s_1), .b(gate116inter3), .O(gate116inter10));
  nor2  gate558(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate559(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate560(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate575(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate576(.a(gate117inter0), .b(s_4), .O(gate117inter1));
  and2  gate577(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate578(.a(s_4), .O(gate117inter3));
  inv1  gate579(.a(s_5), .O(gate117inter4));
  nand2 gate580(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate581(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate582(.a(G386), .O(gate117inter7));
  inv1  gate583(.a(G387), .O(gate117inter8));
  nand2 gate584(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate585(.a(s_5), .b(gate117inter3), .O(gate117inter10));
  nor2  gate586(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate587(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate588(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate589(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate590(.a(gate138inter0), .b(s_6), .O(gate138inter1));
  and2  gate591(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate592(.a(s_6), .O(gate138inter3));
  inv1  gate593(.a(s_7), .O(gate138inter4));
  nand2 gate594(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate595(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate596(.a(G432), .O(gate138inter7));
  inv1  gate597(.a(G435), .O(gate138inter8));
  nand2 gate598(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate599(.a(s_7), .b(gate138inter3), .O(gate138inter10));
  nor2  gate600(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate601(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate602(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1093(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1094(.a(gate143inter0), .b(s_78), .O(gate143inter1));
  and2  gate1095(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1096(.a(s_78), .O(gate143inter3));
  inv1  gate1097(.a(s_79), .O(gate143inter4));
  nand2 gate1098(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1099(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1100(.a(G462), .O(gate143inter7));
  inv1  gate1101(.a(G465), .O(gate143inter8));
  nand2 gate1102(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1103(.a(s_79), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1104(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1105(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1106(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate561(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate562(.a(gate147inter0), .b(s_2), .O(gate147inter1));
  and2  gate563(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate564(.a(s_2), .O(gate147inter3));
  inv1  gate565(.a(s_3), .O(gate147inter4));
  nand2 gate566(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate567(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate568(.a(G486), .O(gate147inter7));
  inv1  gate569(.a(G489), .O(gate147inter8));
  nand2 gate570(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate571(.a(s_3), .b(gate147inter3), .O(gate147inter10));
  nor2  gate572(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate573(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate574(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate925(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate926(.a(gate150inter0), .b(s_54), .O(gate150inter1));
  and2  gate927(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate928(.a(s_54), .O(gate150inter3));
  inv1  gate929(.a(s_55), .O(gate150inter4));
  nand2 gate930(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate931(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate932(.a(G504), .O(gate150inter7));
  inv1  gate933(.a(G507), .O(gate150inter8));
  nand2 gate934(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate935(.a(s_55), .b(gate150inter3), .O(gate150inter10));
  nor2  gate936(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate937(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate938(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1023(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1024(.a(gate155inter0), .b(s_68), .O(gate155inter1));
  and2  gate1025(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1026(.a(s_68), .O(gate155inter3));
  inv1  gate1027(.a(s_69), .O(gate155inter4));
  nand2 gate1028(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1029(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1030(.a(G432), .O(gate155inter7));
  inv1  gate1031(.a(G525), .O(gate155inter8));
  nand2 gate1032(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1033(.a(s_69), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1034(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1035(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1036(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate911(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate912(.a(gate169inter0), .b(s_52), .O(gate169inter1));
  and2  gate913(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate914(.a(s_52), .O(gate169inter3));
  inv1  gate915(.a(s_53), .O(gate169inter4));
  nand2 gate916(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate917(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate918(.a(G474), .O(gate169inter7));
  inv1  gate919(.a(G546), .O(gate169inter8));
  nand2 gate920(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate921(.a(s_53), .b(gate169inter3), .O(gate169inter10));
  nor2  gate922(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate923(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate924(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate757(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate758(.a(gate170inter0), .b(s_30), .O(gate170inter1));
  and2  gate759(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate760(.a(s_30), .O(gate170inter3));
  inv1  gate761(.a(s_31), .O(gate170inter4));
  nand2 gate762(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate763(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate764(.a(G477), .O(gate170inter7));
  inv1  gate765(.a(G546), .O(gate170inter8));
  nand2 gate766(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate767(.a(s_31), .b(gate170inter3), .O(gate170inter10));
  nor2  gate768(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate769(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate770(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate743(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate744(.a(gate171inter0), .b(s_28), .O(gate171inter1));
  and2  gate745(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate746(.a(s_28), .O(gate171inter3));
  inv1  gate747(.a(s_29), .O(gate171inter4));
  nand2 gate748(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate749(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate750(.a(G480), .O(gate171inter7));
  inv1  gate751(.a(G549), .O(gate171inter8));
  nand2 gate752(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate753(.a(s_29), .b(gate171inter3), .O(gate171inter10));
  nor2  gate754(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate755(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate756(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate701(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate702(.a(gate218inter0), .b(s_22), .O(gate218inter1));
  and2  gate703(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate704(.a(s_22), .O(gate218inter3));
  inv1  gate705(.a(s_23), .O(gate218inter4));
  nand2 gate706(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate707(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate708(.a(G627), .O(gate218inter7));
  inv1  gate709(.a(G678), .O(gate218inter8));
  nand2 gate710(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate711(.a(s_23), .b(gate218inter3), .O(gate218inter10));
  nor2  gate712(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate713(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate714(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1247(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1248(.a(gate227inter0), .b(s_100), .O(gate227inter1));
  and2  gate1249(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1250(.a(s_100), .O(gate227inter3));
  inv1  gate1251(.a(s_101), .O(gate227inter4));
  nand2 gate1252(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1253(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1254(.a(G694), .O(gate227inter7));
  inv1  gate1255(.a(G695), .O(gate227inter8));
  nand2 gate1256(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1257(.a(s_101), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1258(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1259(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1260(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1163(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1164(.a(gate238inter0), .b(s_88), .O(gate238inter1));
  and2  gate1165(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1166(.a(s_88), .O(gate238inter3));
  inv1  gate1167(.a(s_89), .O(gate238inter4));
  nand2 gate1168(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1169(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1170(.a(G257), .O(gate238inter7));
  inv1  gate1171(.a(G709), .O(gate238inter8));
  nand2 gate1172(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1173(.a(s_89), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1174(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1175(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1176(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate897(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate898(.a(gate263inter0), .b(s_50), .O(gate263inter1));
  and2  gate899(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate900(.a(s_50), .O(gate263inter3));
  inv1  gate901(.a(s_51), .O(gate263inter4));
  nand2 gate902(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate903(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate904(.a(G766), .O(gate263inter7));
  inv1  gate905(.a(G767), .O(gate263inter8));
  nand2 gate906(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate907(.a(s_51), .b(gate263inter3), .O(gate263inter10));
  nor2  gate908(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate909(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate910(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate953(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate954(.a(gate265inter0), .b(s_58), .O(gate265inter1));
  and2  gate955(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate956(.a(s_58), .O(gate265inter3));
  inv1  gate957(.a(s_59), .O(gate265inter4));
  nand2 gate958(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate959(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate960(.a(G642), .O(gate265inter7));
  inv1  gate961(.a(G770), .O(gate265inter8));
  nand2 gate962(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate963(.a(s_59), .b(gate265inter3), .O(gate265inter10));
  nor2  gate964(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate965(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate966(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1121(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1122(.a(gate269inter0), .b(s_82), .O(gate269inter1));
  and2  gate1123(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1124(.a(s_82), .O(gate269inter3));
  inv1  gate1125(.a(s_83), .O(gate269inter4));
  nand2 gate1126(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1127(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1128(.a(G654), .O(gate269inter7));
  inv1  gate1129(.a(G782), .O(gate269inter8));
  nand2 gate1130(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1131(.a(s_83), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1132(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1133(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1134(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate631(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate632(.a(gate278inter0), .b(s_12), .O(gate278inter1));
  and2  gate633(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate634(.a(s_12), .O(gate278inter3));
  inv1  gate635(.a(s_13), .O(gate278inter4));
  nand2 gate636(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate637(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate638(.a(G776), .O(gate278inter7));
  inv1  gate639(.a(G800), .O(gate278inter8));
  nand2 gate640(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate641(.a(s_13), .b(gate278inter3), .O(gate278inter10));
  nor2  gate642(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate643(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate644(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate645(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate646(.a(gate279inter0), .b(s_14), .O(gate279inter1));
  and2  gate647(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate648(.a(s_14), .O(gate279inter3));
  inv1  gate649(.a(s_15), .O(gate279inter4));
  nand2 gate650(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate651(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate652(.a(G651), .O(gate279inter7));
  inv1  gate653(.a(G803), .O(gate279inter8));
  nand2 gate654(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate655(.a(s_15), .b(gate279inter3), .O(gate279inter10));
  nor2  gate656(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate657(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate658(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1191(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1192(.a(gate285inter0), .b(s_92), .O(gate285inter1));
  and2  gate1193(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1194(.a(s_92), .O(gate285inter3));
  inv1  gate1195(.a(s_93), .O(gate285inter4));
  nand2 gate1196(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1197(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1198(.a(G660), .O(gate285inter7));
  inv1  gate1199(.a(G812), .O(gate285inter8));
  nand2 gate1200(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1201(.a(s_93), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1202(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1203(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1204(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate981(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate982(.a(gate296inter0), .b(s_62), .O(gate296inter1));
  and2  gate983(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate984(.a(s_62), .O(gate296inter3));
  inv1  gate985(.a(s_63), .O(gate296inter4));
  nand2 gate986(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate987(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate988(.a(G826), .O(gate296inter7));
  inv1  gate989(.a(G827), .O(gate296inter8));
  nand2 gate990(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate991(.a(s_63), .b(gate296inter3), .O(gate296inter10));
  nor2  gate992(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate993(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate994(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1177(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1178(.a(gate392inter0), .b(s_90), .O(gate392inter1));
  and2  gate1179(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1180(.a(s_90), .O(gate392inter3));
  inv1  gate1181(.a(s_91), .O(gate392inter4));
  nand2 gate1182(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1183(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1184(.a(G6), .O(gate392inter7));
  inv1  gate1185(.a(G1051), .O(gate392inter8));
  nand2 gate1186(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1187(.a(s_91), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1188(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1189(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1190(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate799(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate800(.a(gate394inter0), .b(s_36), .O(gate394inter1));
  and2  gate801(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate802(.a(s_36), .O(gate394inter3));
  inv1  gate803(.a(s_37), .O(gate394inter4));
  nand2 gate804(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate805(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate806(.a(G8), .O(gate394inter7));
  inv1  gate807(.a(G1057), .O(gate394inter8));
  nand2 gate808(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate809(.a(s_37), .b(gate394inter3), .O(gate394inter10));
  nor2  gate810(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate811(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate812(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1051(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1052(.a(gate399inter0), .b(s_72), .O(gate399inter1));
  and2  gate1053(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1054(.a(s_72), .O(gate399inter3));
  inv1  gate1055(.a(s_73), .O(gate399inter4));
  nand2 gate1056(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1057(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1058(.a(G13), .O(gate399inter7));
  inv1  gate1059(.a(G1072), .O(gate399inter8));
  nand2 gate1060(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1061(.a(s_73), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1062(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1063(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1064(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate729(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate730(.a(gate409inter0), .b(s_26), .O(gate409inter1));
  and2  gate731(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate732(.a(s_26), .O(gate409inter3));
  inv1  gate733(.a(s_27), .O(gate409inter4));
  nand2 gate734(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate735(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate736(.a(G23), .O(gate409inter7));
  inv1  gate737(.a(G1102), .O(gate409inter8));
  nand2 gate738(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate739(.a(s_27), .b(gate409inter3), .O(gate409inter10));
  nor2  gate740(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate741(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate742(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate855(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate856(.a(gate420inter0), .b(s_44), .O(gate420inter1));
  and2  gate857(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate858(.a(s_44), .O(gate420inter3));
  inv1  gate859(.a(s_45), .O(gate420inter4));
  nand2 gate860(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate861(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate862(.a(G1036), .O(gate420inter7));
  inv1  gate863(.a(G1132), .O(gate420inter8));
  nand2 gate864(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate865(.a(s_45), .b(gate420inter3), .O(gate420inter10));
  nor2  gate866(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate867(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate868(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate785(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate786(.a(gate422inter0), .b(s_34), .O(gate422inter1));
  and2  gate787(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate788(.a(s_34), .O(gate422inter3));
  inv1  gate789(.a(s_35), .O(gate422inter4));
  nand2 gate790(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate791(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate792(.a(G1039), .O(gate422inter7));
  inv1  gate793(.a(G1135), .O(gate422inter8));
  nand2 gate794(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate795(.a(s_35), .b(gate422inter3), .O(gate422inter10));
  nor2  gate796(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate797(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate798(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1149(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1150(.a(gate430inter0), .b(s_86), .O(gate430inter1));
  and2  gate1151(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1152(.a(s_86), .O(gate430inter3));
  inv1  gate1153(.a(s_87), .O(gate430inter4));
  nand2 gate1154(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1155(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1156(.a(G1051), .O(gate430inter7));
  inv1  gate1157(.a(G1147), .O(gate430inter8));
  nand2 gate1158(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1159(.a(s_87), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1160(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1161(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1162(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1233(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1234(.a(gate433inter0), .b(s_98), .O(gate433inter1));
  and2  gate1235(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1236(.a(s_98), .O(gate433inter3));
  inv1  gate1237(.a(s_99), .O(gate433inter4));
  nand2 gate1238(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1239(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1240(.a(G8), .O(gate433inter7));
  inv1  gate1241(.a(G1153), .O(gate433inter8));
  nand2 gate1242(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1243(.a(s_99), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1244(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1245(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1246(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1205(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1206(.a(gate457inter0), .b(s_94), .O(gate457inter1));
  and2  gate1207(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1208(.a(s_94), .O(gate457inter3));
  inv1  gate1209(.a(s_95), .O(gate457inter4));
  nand2 gate1210(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1211(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1212(.a(G20), .O(gate457inter7));
  inv1  gate1213(.a(G1189), .O(gate457inter8));
  nand2 gate1214(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1215(.a(s_95), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1216(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1217(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1218(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate687(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate688(.a(gate473inter0), .b(s_20), .O(gate473inter1));
  and2  gate689(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate690(.a(s_20), .O(gate473inter3));
  inv1  gate691(.a(s_21), .O(gate473inter4));
  nand2 gate692(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate693(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate694(.a(G28), .O(gate473inter7));
  inv1  gate695(.a(G1213), .O(gate473inter8));
  nand2 gate696(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate697(.a(s_21), .b(gate473inter3), .O(gate473inter10));
  nor2  gate698(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate699(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate700(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1135(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1136(.a(gate494inter0), .b(s_84), .O(gate494inter1));
  and2  gate1137(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1138(.a(s_84), .O(gate494inter3));
  inv1  gate1139(.a(s_85), .O(gate494inter4));
  nand2 gate1140(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1141(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1142(.a(G1250), .O(gate494inter7));
  inv1  gate1143(.a(G1251), .O(gate494inter8));
  nand2 gate1144(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1145(.a(s_85), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1146(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1147(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1148(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate617(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate618(.a(gate505inter0), .b(s_10), .O(gate505inter1));
  and2  gate619(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate620(.a(s_10), .O(gate505inter3));
  inv1  gate621(.a(s_11), .O(gate505inter4));
  nand2 gate622(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate623(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate624(.a(G1272), .O(gate505inter7));
  inv1  gate625(.a(G1273), .O(gate505inter8));
  nand2 gate626(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate627(.a(s_11), .b(gate505inter3), .O(gate505inter10));
  nor2  gate628(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate629(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate630(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate715(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate716(.a(gate508inter0), .b(s_24), .O(gate508inter1));
  and2  gate717(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate718(.a(s_24), .O(gate508inter3));
  inv1  gate719(.a(s_25), .O(gate508inter4));
  nand2 gate720(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate721(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate722(.a(G1278), .O(gate508inter7));
  inv1  gate723(.a(G1279), .O(gate508inter8));
  nand2 gate724(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate725(.a(s_25), .b(gate508inter3), .O(gate508inter10));
  nor2  gate726(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate727(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate728(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate603(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate604(.a(gate510inter0), .b(s_8), .O(gate510inter1));
  and2  gate605(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate606(.a(s_8), .O(gate510inter3));
  inv1  gate607(.a(s_9), .O(gate510inter4));
  nand2 gate608(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate609(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate610(.a(G1282), .O(gate510inter7));
  inv1  gate611(.a(G1283), .O(gate510inter8));
  nand2 gate612(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate613(.a(s_9), .b(gate510inter3), .O(gate510inter10));
  nor2  gate614(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate615(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate616(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate883(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate884(.a(gate512inter0), .b(s_48), .O(gate512inter1));
  and2  gate885(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate886(.a(s_48), .O(gate512inter3));
  inv1  gate887(.a(s_49), .O(gate512inter4));
  nand2 gate888(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate889(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate890(.a(G1286), .O(gate512inter7));
  inv1  gate891(.a(G1287), .O(gate512inter8));
  nand2 gate892(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate893(.a(s_49), .b(gate512inter3), .O(gate512inter10));
  nor2  gate894(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate895(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate896(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate939(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate940(.a(gate513inter0), .b(s_56), .O(gate513inter1));
  and2  gate941(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate942(.a(s_56), .O(gate513inter3));
  inv1  gate943(.a(s_57), .O(gate513inter4));
  nand2 gate944(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate945(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate946(.a(G1288), .O(gate513inter7));
  inv1  gate947(.a(G1289), .O(gate513inter8));
  nand2 gate948(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate949(.a(s_57), .b(gate513inter3), .O(gate513inter10));
  nor2  gate950(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate951(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate952(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule