module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate497(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate498(.a(gate19inter0), .b(s_48), .O(gate19inter1));
  and2  gate499(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate500(.a(s_48), .O(gate19inter3));
  inv1  gate501(.a(s_49), .O(gate19inter4));
  nand2 gate502(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate503(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate504(.a(N118), .O(gate19inter7));
  inv1  gate505(.a(N4), .O(gate19inter8));
  nand2 gate506(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate507(.a(s_49), .b(gate19inter3), .O(gate19inter10));
  nor2  gate508(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate509(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate510(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate203(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate204(.a(gate20inter0), .b(s_6), .O(gate20inter1));
  and2  gate205(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate206(.a(s_6), .O(gate20inter3));
  inv1  gate207(.a(s_7), .O(gate20inter4));
  nand2 gate208(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate209(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate210(.a(N8), .O(gate20inter7));
  inv1  gate211(.a(N119), .O(gate20inter8));
  nand2 gate212(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate213(.a(s_7), .b(gate20inter3), .O(gate20inter10));
  nor2  gate214(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate215(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate216(.a(gate20inter12), .b(gate20inter1), .O(N157));

  xor2  gate595(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate596(.a(gate21inter0), .b(s_62), .O(gate21inter1));
  and2  gate597(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate598(.a(s_62), .O(gate21inter3));
  inv1  gate599(.a(s_63), .O(gate21inter4));
  nand2 gate600(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate601(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate602(.a(N14), .O(gate21inter7));
  inv1  gate603(.a(N119), .O(gate21inter8));
  nand2 gate604(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate605(.a(s_63), .b(gate21inter3), .O(gate21inter10));
  nor2  gate606(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate607(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate608(.a(gate21inter12), .b(gate21inter1), .O(N158));

  xor2  gate301(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate302(.a(gate22inter0), .b(s_20), .O(gate22inter1));
  and2  gate303(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate304(.a(s_20), .O(gate22inter3));
  inv1  gate305(.a(s_21), .O(gate22inter4));
  nand2 gate306(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate307(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate308(.a(N122), .O(gate22inter7));
  inv1  gate309(.a(N17), .O(gate22inter8));
  nand2 gate310(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate311(.a(s_21), .b(gate22inter3), .O(gate22inter10));
  nor2  gate312(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate313(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate314(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );

  xor2  gate651(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate652(.a(gate26inter0), .b(s_70), .O(gate26inter1));
  and2  gate653(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate654(.a(s_70), .O(gate26inter3));
  inv1  gate655(.a(s_71), .O(gate26inter4));
  nand2 gate656(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate657(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate658(.a(N138), .O(gate26inter7));
  inv1  gate659(.a(N69), .O(gate26inter8));
  nand2 gate660(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate661(.a(s_71), .b(gate26inter3), .O(gate26inter10));
  nor2  gate662(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate663(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate664(.a(gate26inter12), .b(gate26inter1), .O(N171));
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate287(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate288(.a(gate29inter0), .b(s_18), .O(gate29inter1));
  and2  gate289(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate290(.a(s_18), .O(gate29inter3));
  inv1  gate291(.a(s_19), .O(gate29inter4));
  nand2 gate292(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate293(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate294(.a(N150), .O(gate29inter7));
  inv1  gate295(.a(N108), .O(gate29inter8));
  nand2 gate296(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate297(.a(s_19), .b(gate29inter3), .O(gate29inter10));
  nor2  gate298(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate299(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate300(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate273(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate274(.a(gate32inter0), .b(s_16), .O(gate32inter1));
  and2  gate275(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate276(.a(s_16), .O(gate32inter3));
  inv1  gate277(.a(s_17), .O(gate32inter4));
  nand2 gate278(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate279(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate280(.a(N34), .O(gate32inter7));
  inv1  gate281(.a(N127), .O(gate32inter8));
  nand2 gate282(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate283(.a(s_17), .b(gate32inter3), .O(gate32inter10));
  nor2  gate284(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate285(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate286(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate665(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate666(.a(gate36inter0), .b(s_72), .O(gate36inter1));
  and2  gate667(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate668(.a(s_72), .O(gate36inter3));
  inv1  gate669(.a(s_73), .O(gate36inter4));
  nand2 gate670(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate671(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate672(.a(N60), .O(gate36inter7));
  inv1  gate673(.a(N135), .O(gate36inter8));
  nand2 gate674(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate675(.a(s_73), .b(gate36inter3), .O(gate36inter10));
  nor2  gate676(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate677(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate678(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate175(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate176(.a(gate41inter0), .b(s_2), .O(gate41inter1));
  and2  gate177(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate178(.a(s_2), .O(gate41inter3));
  inv1  gate179(.a(s_3), .O(gate41inter4));
  nand2 gate180(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate181(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate182(.a(N92), .O(gate41inter7));
  inv1  gate183(.a(N143), .O(gate41inter8));
  nand2 gate184(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate185(.a(s_3), .b(gate41inter3), .O(gate41inter10));
  nor2  gate186(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate187(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate188(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate637(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate638(.a(gate43inter0), .b(s_68), .O(gate43inter1));
  and2  gate639(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate640(.a(s_68), .O(gate43inter3));
  inv1  gate641(.a(s_69), .O(gate43inter4));
  nand2 gate642(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate643(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate644(.a(N105), .O(gate43inter7));
  inv1  gate645(.a(N147), .O(gate43inter8));
  nand2 gate646(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate647(.a(s_69), .b(gate43inter3), .O(gate43inter10));
  nor2  gate648(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate649(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate650(.a(gate43inter12), .b(gate43inter1), .O(N196));

  xor2  gate259(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate260(.a(gate44inter0), .b(s_14), .O(gate44inter1));
  and2  gate261(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate262(.a(s_14), .O(gate44inter3));
  inv1  gate263(.a(s_15), .O(gate44inter4));
  nand2 gate264(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate265(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate266(.a(N112), .O(gate44inter7));
  inv1  gate267(.a(N151), .O(gate44inter8));
  nand2 gate268(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate269(.a(s_15), .b(gate44inter3), .O(gate44inter10));
  nor2  gate270(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate271(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate272(.a(gate44inter12), .b(gate44inter1), .O(N197));
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate469(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate470(.a(gate52inter0), .b(s_44), .O(gate52inter1));
  and2  gate471(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate472(.a(s_44), .O(gate52inter3));
  inv1  gate473(.a(s_45), .O(gate52inter4));
  nand2 gate474(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate475(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate476(.a(N203), .O(gate52inter7));
  inv1  gate477(.a(N162), .O(gate52inter8));
  nand2 gate478(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate479(.a(s_45), .b(gate52inter3), .O(gate52inter10));
  nor2  gate480(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate481(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate482(.a(gate52inter12), .b(gate52inter1), .O(N230));

  xor2  gate623(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate624(.a(gate53inter0), .b(s_66), .O(gate53inter1));
  and2  gate625(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate626(.a(s_66), .O(gate53inter3));
  inv1  gate627(.a(s_67), .O(gate53inter4));
  nand2 gate628(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate629(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate630(.a(N203), .O(gate53inter7));
  inv1  gate631(.a(N165), .O(gate53inter8));
  nand2 gate632(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate633(.a(s_67), .b(gate53inter3), .O(gate53inter10));
  nor2  gate634(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate635(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate636(.a(gate53inter12), .b(gate53inter1), .O(N233));

  xor2  gate357(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate358(.a(gate54inter0), .b(s_28), .O(gate54inter1));
  and2  gate359(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate360(.a(s_28), .O(gate54inter3));
  inv1  gate361(.a(s_29), .O(gate54inter4));
  nand2 gate362(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate363(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate364(.a(N203), .O(gate54inter7));
  inv1  gate365(.a(N168), .O(gate54inter8));
  nand2 gate366(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate367(.a(s_29), .b(gate54inter3), .O(gate54inter10));
  nor2  gate368(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate369(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate370(.a(gate54inter12), .b(gate54inter1), .O(N236));
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate693(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate694(.a(gate57inter0), .b(s_76), .O(gate57inter1));
  and2  gate695(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate696(.a(s_76), .O(gate57inter3));
  inv1  gate697(.a(s_77), .O(gate57inter4));
  nand2 gate698(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate699(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate700(.a(N203), .O(gate57inter7));
  inv1  gate701(.a(N174), .O(gate57inter8));
  nand2 gate702(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate703(.a(s_77), .b(gate57inter3), .O(gate57inter10));
  nor2  gate704(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate705(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate706(.a(gate57inter12), .b(gate57inter1), .O(N243));

  xor2  gate161(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate162(.a(gate58inter0), .b(s_0), .O(gate58inter1));
  and2  gate163(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate164(.a(s_0), .O(gate58inter3));
  inv1  gate165(.a(s_1), .O(gate58inter4));
  nand2 gate166(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate167(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate168(.a(N213), .O(gate58inter7));
  inv1  gate169(.a(N11), .O(gate58inter8));
  nand2 gate170(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate171(.a(s_1), .b(gate58inter3), .O(gate58inter10));
  nor2  gate172(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate173(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate174(.a(gate58inter12), .b(gate58inter1), .O(N246));
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate539(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate540(.a(gate60inter0), .b(s_54), .O(gate60inter1));
  and2  gate541(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate542(.a(s_54), .O(gate60inter3));
  inv1  gate543(.a(s_55), .O(gate60inter4));
  nand2 gate544(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate545(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate546(.a(N213), .O(gate60inter7));
  inv1  gate547(.a(N24), .O(gate60inter8));
  nand2 gate548(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate549(.a(s_55), .b(gate60inter3), .O(gate60inter10));
  nor2  gate550(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate551(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate552(.a(gate60inter12), .b(gate60inter1), .O(N250));
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate343(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate344(.a(gate62inter0), .b(s_26), .O(gate62inter1));
  and2  gate345(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate346(.a(s_26), .O(gate62inter3));
  inv1  gate347(.a(s_27), .O(gate62inter4));
  nand2 gate348(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate349(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate350(.a(N213), .O(gate62inter7));
  inv1  gate351(.a(N37), .O(gate62inter8));
  nand2 gate352(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate353(.a(s_27), .b(gate62inter3), .O(gate62inter10));
  nor2  gate354(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate355(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate356(.a(gate62inter12), .b(gate62inter1), .O(N254));
nand2 gate63( .a(N213), .b(N50), .O(N255) );

  xor2  gate511(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate512(.a(gate64inter0), .b(s_50), .O(gate64inter1));
  and2  gate513(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate514(.a(s_50), .O(gate64inter3));
  inv1  gate515(.a(s_51), .O(gate64inter4));
  nand2 gate516(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate517(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate518(.a(N213), .O(gate64inter7));
  inv1  gate519(.a(N63), .O(gate64inter8));
  nand2 gate520(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate521(.a(s_51), .b(gate64inter3), .O(gate64inter10));
  nor2  gate522(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate523(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate524(.a(gate64inter12), .b(gate64inter1), .O(N256));
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate567(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate568(.a(gate73inter0), .b(s_58), .O(gate73inter1));
  and2  gate569(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate570(.a(s_58), .O(gate73inter3));
  inv1  gate571(.a(s_59), .O(gate73inter4));
  nand2 gate572(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate573(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate574(.a(N236), .O(gate73inter7));
  inv1  gate575(.a(N189), .O(gate73inter8));
  nand2 gate576(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate577(.a(s_59), .b(gate73inter3), .O(gate73inter10));
  nor2  gate578(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate579(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate580(.a(gate73inter12), .b(gate73inter1), .O(N273));

  xor2  gate679(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate680(.a(gate74inter0), .b(s_74), .O(gate74inter1));
  and2  gate681(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate682(.a(s_74), .O(gate74inter3));
  inv1  gate683(.a(s_75), .O(gate74inter4));
  nand2 gate684(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate685(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate686(.a(N239), .O(gate74inter7));
  inv1  gate687(.a(N191), .O(gate74inter8));
  nand2 gate688(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate689(.a(s_75), .b(gate74inter3), .O(gate74inter10));
  nor2  gate690(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate691(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate692(.a(gate74inter12), .b(gate74inter1), .O(N276));

  xor2  gate707(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate708(.a(gate75inter0), .b(s_78), .O(gate75inter1));
  and2  gate709(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate710(.a(s_78), .O(gate75inter3));
  inv1  gate711(.a(s_79), .O(gate75inter4));
  nand2 gate712(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate713(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate714(.a(N243), .O(gate75inter7));
  inv1  gate715(.a(N193), .O(gate75inter8));
  nand2 gate716(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate717(.a(s_79), .b(gate75inter3), .O(gate75inter10));
  nor2  gate718(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate719(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate720(.a(gate75inter12), .b(gate75inter1), .O(N279));

  xor2  gate217(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate218(.a(gate76inter0), .b(s_8), .O(gate76inter1));
  and2  gate219(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate220(.a(s_8), .O(gate76inter3));
  inv1  gate221(.a(s_9), .O(gate76inter4));
  nand2 gate222(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate223(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate224(.a(N247), .O(gate76inter7));
  inv1  gate225(.a(N195), .O(gate76inter8));
  nand2 gate226(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate227(.a(s_9), .b(gate76inter3), .O(gate76inter10));
  nor2  gate228(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate229(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate230(.a(gate76inter12), .b(gate76inter1), .O(N282));
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate721(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate722(.a(gate80inter0), .b(s_80), .O(gate80inter1));
  and2  gate723(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate724(.a(s_80), .O(gate80inter3));
  inv1  gate725(.a(s_81), .O(gate80inter4));
  nand2 gate726(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate727(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate728(.a(N233), .O(gate80inter7));
  inv1  gate729(.a(N188), .O(gate80inter8));
  nand2 gate730(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate731(.a(s_81), .b(gate80inter3), .O(gate80inter10));
  nor2  gate732(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate733(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate734(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );

  xor2  gate581(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate582(.a(gate82inter0), .b(s_60), .O(gate82inter1));
  and2  gate583(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate584(.a(s_60), .O(gate82inter3));
  inv1  gate585(.a(s_61), .O(gate82inter4));
  nand2 gate586(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate587(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate588(.a(N239), .O(gate82inter7));
  inv1  gate589(.a(N192), .O(gate82inter8));
  nand2 gate590(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate591(.a(s_61), .b(gate82inter3), .O(gate82inter10));
  nor2  gate592(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate593(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate594(.a(gate82inter12), .b(gate82inter1), .O(N292));

  xor2  gate371(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate372(.a(gate83inter0), .b(s_30), .O(gate83inter1));
  and2  gate373(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate374(.a(s_30), .O(gate83inter3));
  inv1  gate375(.a(s_31), .O(gate83inter4));
  nand2 gate376(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate377(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate378(.a(N243), .O(gate83inter7));
  inv1  gate379(.a(N194), .O(gate83inter8));
  nand2 gate380(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate381(.a(s_31), .b(gate83inter3), .O(gate83inter10));
  nor2  gate382(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate383(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate384(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );

  xor2  gate609(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate610(.a(gate101inter0), .b(s_64), .O(gate101inter1));
  and2  gate611(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate612(.a(s_64), .O(gate101inter3));
  inv1  gate613(.a(s_65), .O(gate101inter4));
  nand2 gate614(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate615(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate616(.a(N309), .O(gate101inter7));
  inv1  gate617(.a(N267), .O(gate101inter8));
  nand2 gate618(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate619(.a(s_65), .b(gate101inter3), .O(gate101inter10));
  nor2  gate620(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate621(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate622(.a(gate101inter12), .b(gate101inter1), .O(N332));
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate315(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate316(.a(gate103inter0), .b(s_22), .O(gate103inter1));
  and2  gate317(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate318(.a(s_22), .O(gate103inter3));
  inv1  gate319(.a(s_23), .O(gate103inter4));
  nand2 gate320(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate321(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate322(.a(N8), .O(gate103inter7));
  inv1  gate323(.a(N319), .O(gate103inter8));
  nand2 gate324(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate325(.a(s_23), .b(gate103inter3), .O(gate103inter10));
  nor2  gate326(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate327(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate328(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate441(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate442(.a(gate105inter0), .b(s_40), .O(gate105inter1));
  and2  gate443(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate444(.a(s_40), .O(gate105inter3));
  inv1  gate445(.a(s_41), .O(gate105inter4));
  nand2 gate446(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate447(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate448(.a(N319), .O(gate105inter7));
  inv1  gate449(.a(N21), .O(gate105inter8));
  nand2 gate450(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate451(.a(s_41), .b(gate105inter3), .O(gate105inter10));
  nor2  gate452(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate453(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate454(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );

  xor2  gate329(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate330(.a(gate109inter0), .b(s_24), .O(gate109inter1));
  and2  gate331(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate332(.a(s_24), .O(gate109inter3));
  inv1  gate333(.a(s_25), .O(gate109inter4));
  nand2 gate334(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate335(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate336(.a(N319), .O(gate109inter7));
  inv1  gate337(.a(N47), .O(gate109inter8));
  nand2 gate338(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate339(.a(s_25), .b(gate109inter3), .O(gate109inter10));
  nor2  gate340(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate341(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate342(.a(gate109inter12), .b(gate109inter1), .O(N340));

  xor2  gate189(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate190(.a(gate110inter0), .b(s_4), .O(gate110inter1));
  and2  gate191(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate192(.a(s_4), .O(gate110inter3));
  inv1  gate193(.a(s_5), .O(gate110inter4));
  nand2 gate194(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate195(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate196(.a(N309), .O(gate110inter7));
  inv1  gate197(.a(N282), .O(gate110inter8));
  nand2 gate198(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate199(.a(s_5), .b(gate110inter3), .O(gate110inter10));
  nor2  gate200(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate201(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate202(.a(gate110inter12), .b(gate110inter1), .O(N341));

  xor2  gate427(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate428(.a(gate111inter0), .b(s_38), .O(gate111inter1));
  and2  gate429(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate430(.a(s_38), .O(gate111inter3));
  inv1  gate431(.a(s_39), .O(gate111inter4));
  nand2 gate432(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate433(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate434(.a(N319), .O(gate111inter7));
  inv1  gate435(.a(N60), .O(gate111inter8));
  nand2 gate436(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate437(.a(s_39), .b(gate111inter3), .O(gate111inter10));
  nor2  gate438(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate439(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate440(.a(gate111inter12), .b(gate111inter1), .O(N342));

  xor2  gate455(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate456(.a(gate112inter0), .b(s_42), .O(gate112inter1));
  and2  gate457(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate458(.a(s_42), .O(gate112inter3));
  inv1  gate459(.a(s_43), .O(gate112inter4));
  nand2 gate460(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate461(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate462(.a(N309), .O(gate112inter7));
  inv1  gate463(.a(N285), .O(gate112inter8));
  nand2 gate464(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate465(.a(s_43), .b(gate112inter3), .O(gate112inter10));
  nor2  gate466(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate467(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate468(.a(gate112inter12), .b(gate112inter1), .O(N343));

  xor2  gate525(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate526(.a(gate113inter0), .b(s_52), .O(gate113inter1));
  and2  gate527(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate528(.a(s_52), .O(gate113inter3));
  inv1  gate529(.a(s_53), .O(gate113inter4));
  nand2 gate530(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate531(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate532(.a(N319), .O(gate113inter7));
  inv1  gate533(.a(N73), .O(gate113inter8));
  nand2 gate534(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate535(.a(s_53), .b(gate113inter3), .O(gate113inter10));
  nor2  gate536(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate537(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate538(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );

  xor2  gate245(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate246(.a(gate122inter0), .b(s_12), .O(gate122inter1));
  and2  gate247(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate248(.a(s_12), .O(gate122inter3));
  inv1  gate249(.a(s_13), .O(gate122inter4));
  nand2 gate250(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate251(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate252(.a(N337), .O(gate122inter7));
  inv1  gate253(.a(N305), .O(gate122inter8));
  nand2 gate254(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate255(.a(s_13), .b(gate122inter3), .O(gate122inter10));
  nor2  gate256(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate257(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate258(.a(gate122inter12), .b(gate122inter1), .O(N353));

  xor2  gate385(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate386(.a(gate123inter0), .b(s_32), .O(gate123inter1));
  and2  gate387(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate388(.a(s_32), .O(gate123inter3));
  inv1  gate389(.a(s_33), .O(gate123inter4));
  nand2 gate390(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate391(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate392(.a(N339), .O(gate123inter7));
  inv1  gate393(.a(N306), .O(gate123inter8));
  nand2 gate394(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate395(.a(s_33), .b(gate123inter3), .O(gate123inter10));
  nor2  gate396(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate397(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate398(.a(gate123inter12), .b(gate123inter1), .O(N354));

  xor2  gate413(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate414(.a(gate124inter0), .b(s_36), .O(gate124inter1));
  and2  gate415(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate416(.a(s_36), .O(gate124inter3));
  inv1  gate417(.a(s_37), .O(gate124inter4));
  nand2 gate418(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate419(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate420(.a(N341), .O(gate124inter7));
  inv1  gate421(.a(N307), .O(gate124inter8));
  nand2 gate422(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate423(.a(s_37), .b(gate124inter3), .O(gate124inter10));
  nor2  gate424(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate425(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate426(.a(gate124inter12), .b(gate124inter1), .O(N355));

  xor2  gate553(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate554(.a(gate125inter0), .b(s_56), .O(gate125inter1));
  and2  gate555(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate556(.a(s_56), .O(gate125inter3));
  inv1  gate557(.a(s_57), .O(gate125inter4));
  nand2 gate558(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate559(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate560(.a(N343), .O(gate125inter7));
  inv1  gate561(.a(N308), .O(gate125inter8));
  nand2 gate562(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate563(.a(s_57), .b(gate125inter3), .O(gate125inter10));
  nor2  gate564(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate565(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate566(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate483(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate484(.a(gate129inter0), .b(s_46), .O(gate129inter1));
  and2  gate485(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate486(.a(s_46), .O(gate129inter3));
  inv1  gate487(.a(s_47), .O(gate129inter4));
  nand2 gate488(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate489(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate490(.a(N14), .O(gate129inter7));
  inv1  gate491(.a(N360), .O(gate129inter8));
  nand2 gate492(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate493(.a(s_47), .b(gate129inter3), .O(gate129inter10));
  nor2  gate494(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate495(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate496(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );

  xor2  gate399(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate400(.a(gate134inter0), .b(s_34), .O(gate134inter1));
  and2  gate401(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate402(.a(s_34), .O(gate134inter3));
  inv1  gate403(.a(s_35), .O(gate134inter4));
  nand2 gate404(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate405(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate406(.a(N360), .O(gate134inter7));
  inv1  gate407(.a(N79), .O(gate134inter8));
  nand2 gate408(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate409(.a(s_35), .b(gate134inter3), .O(gate134inter10));
  nor2  gate410(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate411(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate412(.a(gate134inter12), .b(gate134inter1), .O(N376));

  xor2  gate231(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate232(.a(gate135inter0), .b(s_10), .O(gate135inter1));
  and2  gate233(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate234(.a(s_10), .O(gate135inter3));
  inv1  gate235(.a(s_11), .O(gate135inter4));
  nand2 gate236(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate237(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate238(.a(N360), .O(gate135inter7));
  inv1  gate239(.a(N92), .O(gate135inter8));
  nand2 gate240(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate241(.a(s_11), .b(gate135inter3), .O(gate135inter10));
  nor2  gate242(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate243(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate244(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule