module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate953(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate954(.a(gate11inter0), .b(s_58), .O(gate11inter1));
  and2  gate955(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate956(.a(s_58), .O(gate11inter3));
  inv1  gate957(.a(s_59), .O(gate11inter4));
  nand2 gate958(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate959(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate960(.a(G5), .O(gate11inter7));
  inv1  gate961(.a(G6), .O(gate11inter8));
  nand2 gate962(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate963(.a(s_59), .b(gate11inter3), .O(gate11inter10));
  nor2  gate964(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate965(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate966(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2115(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2116(.a(gate14inter0), .b(s_224), .O(gate14inter1));
  and2  gate2117(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2118(.a(s_224), .O(gate14inter3));
  inv1  gate2119(.a(s_225), .O(gate14inter4));
  nand2 gate2120(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2121(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2122(.a(G11), .O(gate14inter7));
  inv1  gate2123(.a(G12), .O(gate14inter8));
  nand2 gate2124(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2125(.a(s_225), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2126(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2127(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2128(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate575(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate576(.a(gate18inter0), .b(s_4), .O(gate18inter1));
  and2  gate577(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate578(.a(s_4), .O(gate18inter3));
  inv1  gate579(.a(s_5), .O(gate18inter4));
  nand2 gate580(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate581(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate582(.a(G19), .O(gate18inter7));
  inv1  gate583(.a(G20), .O(gate18inter8));
  nand2 gate584(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate585(.a(s_5), .b(gate18inter3), .O(gate18inter10));
  nor2  gate586(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate587(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate588(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2227(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2228(.a(gate19inter0), .b(s_240), .O(gate19inter1));
  and2  gate2229(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2230(.a(s_240), .O(gate19inter3));
  inv1  gate2231(.a(s_241), .O(gate19inter4));
  nand2 gate2232(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2233(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2234(.a(G21), .O(gate19inter7));
  inv1  gate2235(.a(G22), .O(gate19inter8));
  nand2 gate2236(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2237(.a(s_241), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2238(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2239(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2240(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2283(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2284(.a(gate21inter0), .b(s_248), .O(gate21inter1));
  and2  gate2285(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2286(.a(s_248), .O(gate21inter3));
  inv1  gate2287(.a(s_249), .O(gate21inter4));
  nand2 gate2288(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2289(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2290(.a(G25), .O(gate21inter7));
  inv1  gate2291(.a(G26), .O(gate21inter8));
  nand2 gate2292(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2293(.a(s_249), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2294(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2295(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2296(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1401(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1402(.a(gate28inter0), .b(s_122), .O(gate28inter1));
  and2  gate1403(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1404(.a(s_122), .O(gate28inter3));
  inv1  gate1405(.a(s_123), .O(gate28inter4));
  nand2 gate1406(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1407(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1408(.a(G10), .O(gate28inter7));
  inv1  gate1409(.a(G14), .O(gate28inter8));
  nand2 gate1410(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1411(.a(s_123), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1412(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1413(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1414(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate631(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate632(.a(gate37inter0), .b(s_12), .O(gate37inter1));
  and2  gate633(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate634(.a(s_12), .O(gate37inter3));
  inv1  gate635(.a(s_13), .O(gate37inter4));
  nand2 gate636(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate637(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate638(.a(G19), .O(gate37inter7));
  inv1  gate639(.a(G23), .O(gate37inter8));
  nand2 gate640(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate641(.a(s_13), .b(gate37inter3), .O(gate37inter10));
  nor2  gate642(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate643(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate644(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate799(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate800(.a(gate39inter0), .b(s_36), .O(gate39inter1));
  and2  gate801(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate802(.a(s_36), .O(gate39inter3));
  inv1  gate803(.a(s_37), .O(gate39inter4));
  nand2 gate804(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate805(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate806(.a(G20), .O(gate39inter7));
  inv1  gate807(.a(G24), .O(gate39inter8));
  nand2 gate808(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate809(.a(s_37), .b(gate39inter3), .O(gate39inter10));
  nor2  gate810(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate811(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate812(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate981(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate982(.a(gate40inter0), .b(s_62), .O(gate40inter1));
  and2  gate983(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate984(.a(s_62), .O(gate40inter3));
  inv1  gate985(.a(s_63), .O(gate40inter4));
  nand2 gate986(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate987(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate988(.a(G28), .O(gate40inter7));
  inv1  gate989(.a(G32), .O(gate40inter8));
  nand2 gate990(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate991(.a(s_63), .b(gate40inter3), .O(gate40inter10));
  nor2  gate992(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate993(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate994(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1933(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1934(.a(gate43inter0), .b(s_198), .O(gate43inter1));
  and2  gate1935(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1936(.a(s_198), .O(gate43inter3));
  inv1  gate1937(.a(s_199), .O(gate43inter4));
  nand2 gate1938(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1939(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1940(.a(G3), .O(gate43inter7));
  inv1  gate1941(.a(G269), .O(gate43inter8));
  nand2 gate1942(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1943(.a(s_199), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1944(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1945(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1946(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1471(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1472(.a(gate48inter0), .b(s_132), .O(gate48inter1));
  and2  gate1473(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1474(.a(s_132), .O(gate48inter3));
  inv1  gate1475(.a(s_133), .O(gate48inter4));
  nand2 gate1476(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1477(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1478(.a(G8), .O(gate48inter7));
  inv1  gate1479(.a(G275), .O(gate48inter8));
  nand2 gate1480(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1481(.a(s_133), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1482(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1483(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1484(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1023(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1024(.a(gate50inter0), .b(s_68), .O(gate50inter1));
  and2  gate1025(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1026(.a(s_68), .O(gate50inter3));
  inv1  gate1027(.a(s_69), .O(gate50inter4));
  nand2 gate1028(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1029(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1030(.a(G10), .O(gate50inter7));
  inv1  gate1031(.a(G278), .O(gate50inter8));
  nand2 gate1032(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1033(.a(s_69), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1034(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1035(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1036(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1919(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1920(.a(gate52inter0), .b(s_196), .O(gate52inter1));
  and2  gate1921(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1922(.a(s_196), .O(gate52inter3));
  inv1  gate1923(.a(s_197), .O(gate52inter4));
  nand2 gate1924(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1925(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1926(.a(G12), .O(gate52inter7));
  inv1  gate1927(.a(G281), .O(gate52inter8));
  nand2 gate1928(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1929(.a(s_197), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1930(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1931(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1932(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1527(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1528(.a(gate53inter0), .b(s_140), .O(gate53inter1));
  and2  gate1529(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1530(.a(s_140), .O(gate53inter3));
  inv1  gate1531(.a(s_141), .O(gate53inter4));
  nand2 gate1532(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1533(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1534(.a(G13), .O(gate53inter7));
  inv1  gate1535(.a(G284), .O(gate53inter8));
  nand2 gate1536(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1537(.a(s_141), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1538(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1539(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1540(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1135(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1136(.a(gate54inter0), .b(s_84), .O(gate54inter1));
  and2  gate1137(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1138(.a(s_84), .O(gate54inter3));
  inv1  gate1139(.a(s_85), .O(gate54inter4));
  nand2 gate1140(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1141(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1142(.a(G14), .O(gate54inter7));
  inv1  gate1143(.a(G284), .O(gate54inter8));
  nand2 gate1144(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1145(.a(s_85), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1146(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1147(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1148(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate911(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate912(.a(gate55inter0), .b(s_52), .O(gate55inter1));
  and2  gate913(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate914(.a(s_52), .O(gate55inter3));
  inv1  gate915(.a(s_53), .O(gate55inter4));
  nand2 gate916(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate917(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate918(.a(G15), .O(gate55inter7));
  inv1  gate919(.a(G287), .O(gate55inter8));
  nand2 gate920(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate921(.a(s_53), .b(gate55inter3), .O(gate55inter10));
  nor2  gate922(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate923(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate924(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1779(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1780(.a(gate59inter0), .b(s_176), .O(gate59inter1));
  and2  gate1781(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1782(.a(s_176), .O(gate59inter3));
  inv1  gate1783(.a(s_177), .O(gate59inter4));
  nand2 gate1784(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1785(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1786(.a(G19), .O(gate59inter7));
  inv1  gate1787(.a(G293), .O(gate59inter8));
  nand2 gate1788(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1789(.a(s_177), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1790(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1791(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1792(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate603(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate604(.a(gate62inter0), .b(s_8), .O(gate62inter1));
  and2  gate605(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate606(.a(s_8), .O(gate62inter3));
  inv1  gate607(.a(s_9), .O(gate62inter4));
  nand2 gate608(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate609(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate610(.a(G22), .O(gate62inter7));
  inv1  gate611(.a(G296), .O(gate62inter8));
  nand2 gate612(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate613(.a(s_9), .b(gate62inter3), .O(gate62inter10));
  nor2  gate614(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate615(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate616(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1555(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1556(.a(gate65inter0), .b(s_144), .O(gate65inter1));
  and2  gate1557(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1558(.a(s_144), .O(gate65inter3));
  inv1  gate1559(.a(s_145), .O(gate65inter4));
  nand2 gate1560(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1561(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1562(.a(G25), .O(gate65inter7));
  inv1  gate1563(.a(G302), .O(gate65inter8));
  nand2 gate1564(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1565(.a(s_145), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1566(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1567(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1568(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate743(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate744(.a(gate69inter0), .b(s_28), .O(gate69inter1));
  and2  gate745(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate746(.a(s_28), .O(gate69inter3));
  inv1  gate747(.a(s_29), .O(gate69inter4));
  nand2 gate748(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate749(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate750(.a(G29), .O(gate69inter7));
  inv1  gate751(.a(G308), .O(gate69inter8));
  nand2 gate752(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate753(.a(s_29), .b(gate69inter3), .O(gate69inter10));
  nor2  gate754(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate755(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate756(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2143(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2144(.a(gate71inter0), .b(s_228), .O(gate71inter1));
  and2  gate2145(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2146(.a(s_228), .O(gate71inter3));
  inv1  gate2147(.a(s_229), .O(gate71inter4));
  nand2 gate2148(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2149(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2150(.a(G31), .O(gate71inter7));
  inv1  gate2151(.a(G311), .O(gate71inter8));
  nand2 gate2152(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2153(.a(s_229), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2154(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2155(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2156(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1289(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1290(.a(gate74inter0), .b(s_106), .O(gate74inter1));
  and2  gate1291(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1292(.a(s_106), .O(gate74inter3));
  inv1  gate1293(.a(s_107), .O(gate74inter4));
  nand2 gate1294(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1295(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1296(.a(G5), .O(gate74inter7));
  inv1  gate1297(.a(G314), .O(gate74inter8));
  nand2 gate1298(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1299(.a(s_107), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1300(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1301(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1302(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1751(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1752(.a(gate80inter0), .b(s_172), .O(gate80inter1));
  and2  gate1753(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1754(.a(s_172), .O(gate80inter3));
  inv1  gate1755(.a(s_173), .O(gate80inter4));
  nand2 gate1756(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1757(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1758(.a(G14), .O(gate80inter7));
  inv1  gate1759(.a(G323), .O(gate80inter8));
  nand2 gate1760(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1761(.a(s_173), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1762(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1763(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1764(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate2185(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2186(.a(gate83inter0), .b(s_234), .O(gate83inter1));
  and2  gate2187(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2188(.a(s_234), .O(gate83inter3));
  inv1  gate2189(.a(s_235), .O(gate83inter4));
  nand2 gate2190(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2191(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2192(.a(G11), .O(gate83inter7));
  inv1  gate2193(.a(G329), .O(gate83inter8));
  nand2 gate2194(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2195(.a(s_235), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2196(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2197(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2198(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1359(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1360(.a(gate85inter0), .b(s_116), .O(gate85inter1));
  and2  gate1361(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1362(.a(s_116), .O(gate85inter3));
  inv1  gate1363(.a(s_117), .O(gate85inter4));
  nand2 gate1364(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1365(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1366(.a(G4), .O(gate85inter7));
  inv1  gate1367(.a(G332), .O(gate85inter8));
  nand2 gate1368(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1369(.a(s_117), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1370(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1371(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1372(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate2031(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2032(.a(gate86inter0), .b(s_212), .O(gate86inter1));
  and2  gate2033(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2034(.a(s_212), .O(gate86inter3));
  inv1  gate2035(.a(s_213), .O(gate86inter4));
  nand2 gate2036(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2037(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2038(.a(G8), .O(gate86inter7));
  inv1  gate2039(.a(G332), .O(gate86inter8));
  nand2 gate2040(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2041(.a(s_213), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2042(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2043(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2044(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1597(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1598(.a(gate87inter0), .b(s_150), .O(gate87inter1));
  and2  gate1599(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1600(.a(s_150), .O(gate87inter3));
  inv1  gate1601(.a(s_151), .O(gate87inter4));
  nand2 gate1602(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1603(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1604(.a(G12), .O(gate87inter7));
  inv1  gate1605(.a(G335), .O(gate87inter8));
  nand2 gate1606(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1607(.a(s_151), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1608(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1609(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1610(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2101(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2102(.a(gate92inter0), .b(s_222), .O(gate92inter1));
  and2  gate2103(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2104(.a(s_222), .O(gate92inter3));
  inv1  gate2105(.a(s_223), .O(gate92inter4));
  nand2 gate2106(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2107(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2108(.a(G29), .O(gate92inter7));
  inv1  gate2109(.a(G341), .O(gate92inter8));
  nand2 gate2110(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2111(.a(s_223), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2112(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2113(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2114(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1093(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1094(.a(gate93inter0), .b(s_78), .O(gate93inter1));
  and2  gate1095(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1096(.a(s_78), .O(gate93inter3));
  inv1  gate1097(.a(s_79), .O(gate93inter4));
  nand2 gate1098(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1099(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1100(.a(G18), .O(gate93inter7));
  inv1  gate1101(.a(G344), .O(gate93inter8));
  nand2 gate1102(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1103(.a(s_79), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1104(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1105(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1106(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2241(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2242(.a(gate95inter0), .b(s_242), .O(gate95inter1));
  and2  gate2243(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2244(.a(s_242), .O(gate95inter3));
  inv1  gate2245(.a(s_243), .O(gate95inter4));
  nand2 gate2246(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2247(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2248(.a(G26), .O(gate95inter7));
  inv1  gate2249(.a(G347), .O(gate95inter8));
  nand2 gate2250(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2251(.a(s_243), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2252(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2253(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2254(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate827(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate828(.a(gate96inter0), .b(s_40), .O(gate96inter1));
  and2  gate829(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate830(.a(s_40), .O(gate96inter3));
  inv1  gate831(.a(s_41), .O(gate96inter4));
  nand2 gate832(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate833(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate834(.a(G30), .O(gate96inter7));
  inv1  gate835(.a(G347), .O(gate96inter8));
  nand2 gate836(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate837(.a(s_41), .b(gate96inter3), .O(gate96inter10));
  nor2  gate838(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate839(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate840(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1709(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1710(.a(gate97inter0), .b(s_166), .O(gate97inter1));
  and2  gate1711(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1712(.a(s_166), .O(gate97inter3));
  inv1  gate1713(.a(s_167), .O(gate97inter4));
  nand2 gate1714(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1715(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1716(.a(G19), .O(gate97inter7));
  inv1  gate1717(.a(G350), .O(gate97inter8));
  nand2 gate1718(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1719(.a(s_167), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1720(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1721(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1722(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1247(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1248(.a(gate98inter0), .b(s_100), .O(gate98inter1));
  and2  gate1249(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1250(.a(s_100), .O(gate98inter3));
  inv1  gate1251(.a(s_101), .O(gate98inter4));
  nand2 gate1252(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1253(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1254(.a(G23), .O(gate98inter7));
  inv1  gate1255(.a(G350), .O(gate98inter8));
  nand2 gate1256(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1257(.a(s_101), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1258(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1259(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1260(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2213(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2214(.a(gate100inter0), .b(s_238), .O(gate100inter1));
  and2  gate2215(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2216(.a(s_238), .O(gate100inter3));
  inv1  gate2217(.a(s_239), .O(gate100inter4));
  nand2 gate2218(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2219(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2220(.a(G31), .O(gate100inter7));
  inv1  gate2221(.a(G353), .O(gate100inter8));
  nand2 gate2222(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2223(.a(s_239), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2224(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2225(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2226(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate589(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate590(.a(gate102inter0), .b(s_6), .O(gate102inter1));
  and2  gate591(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate592(.a(s_6), .O(gate102inter3));
  inv1  gate593(.a(s_7), .O(gate102inter4));
  nand2 gate594(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate595(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate596(.a(G24), .O(gate102inter7));
  inv1  gate597(.a(G356), .O(gate102inter8));
  nand2 gate598(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate599(.a(s_7), .b(gate102inter3), .O(gate102inter10));
  nor2  gate600(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate601(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate602(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate883(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate884(.a(gate105inter0), .b(s_48), .O(gate105inter1));
  and2  gate885(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate886(.a(s_48), .O(gate105inter3));
  inv1  gate887(.a(s_49), .O(gate105inter4));
  nand2 gate888(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate889(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate890(.a(G362), .O(gate105inter7));
  inv1  gate891(.a(G363), .O(gate105inter8));
  nand2 gate892(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate893(.a(s_49), .b(gate105inter3), .O(gate105inter10));
  nor2  gate894(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate895(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate896(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1009(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1010(.a(gate110inter0), .b(s_66), .O(gate110inter1));
  and2  gate1011(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1012(.a(s_66), .O(gate110inter3));
  inv1  gate1013(.a(s_67), .O(gate110inter4));
  nand2 gate1014(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1015(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1016(.a(G372), .O(gate110inter7));
  inv1  gate1017(.a(G373), .O(gate110inter8));
  nand2 gate1018(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1019(.a(s_67), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1020(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1021(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1022(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1219(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1220(.a(gate113inter0), .b(s_96), .O(gate113inter1));
  and2  gate1221(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1222(.a(s_96), .O(gate113inter3));
  inv1  gate1223(.a(s_97), .O(gate113inter4));
  nand2 gate1224(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1225(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1226(.a(G378), .O(gate113inter7));
  inv1  gate1227(.a(G379), .O(gate113inter8));
  nand2 gate1228(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1229(.a(s_97), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1230(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1231(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1232(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1513(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1514(.a(gate115inter0), .b(s_138), .O(gate115inter1));
  and2  gate1515(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1516(.a(s_138), .O(gate115inter3));
  inv1  gate1517(.a(s_139), .O(gate115inter4));
  nand2 gate1518(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1519(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1520(.a(G382), .O(gate115inter7));
  inv1  gate1521(.a(G383), .O(gate115inter8));
  nand2 gate1522(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1523(.a(s_139), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1524(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1525(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1526(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1429(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1430(.a(gate116inter0), .b(s_126), .O(gate116inter1));
  and2  gate1431(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1432(.a(s_126), .O(gate116inter3));
  inv1  gate1433(.a(s_127), .O(gate116inter4));
  nand2 gate1434(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1435(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1436(.a(G384), .O(gate116inter7));
  inv1  gate1437(.a(G385), .O(gate116inter8));
  nand2 gate1438(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1439(.a(s_127), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1440(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1441(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1442(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1947(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1948(.a(gate118inter0), .b(s_200), .O(gate118inter1));
  and2  gate1949(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1950(.a(s_200), .O(gate118inter3));
  inv1  gate1951(.a(s_201), .O(gate118inter4));
  nand2 gate1952(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1953(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1954(.a(G388), .O(gate118inter7));
  inv1  gate1955(.a(G389), .O(gate118inter8));
  nand2 gate1956(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1957(.a(s_201), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1958(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1959(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1960(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate561(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate562(.a(gate123inter0), .b(s_2), .O(gate123inter1));
  and2  gate563(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate564(.a(s_2), .O(gate123inter3));
  inv1  gate565(.a(s_3), .O(gate123inter4));
  nand2 gate566(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate567(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate568(.a(G398), .O(gate123inter7));
  inv1  gate569(.a(G399), .O(gate123inter8));
  nand2 gate570(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate571(.a(s_3), .b(gate123inter3), .O(gate123inter10));
  nor2  gate572(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate573(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate574(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1051(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1052(.a(gate125inter0), .b(s_72), .O(gate125inter1));
  and2  gate1053(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1054(.a(s_72), .O(gate125inter3));
  inv1  gate1055(.a(s_73), .O(gate125inter4));
  nand2 gate1056(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1057(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1058(.a(G402), .O(gate125inter7));
  inv1  gate1059(.a(G403), .O(gate125inter8));
  nand2 gate1060(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1061(.a(s_73), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1062(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1063(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1064(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1107(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1108(.a(gate128inter0), .b(s_80), .O(gate128inter1));
  and2  gate1109(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1110(.a(s_80), .O(gate128inter3));
  inv1  gate1111(.a(s_81), .O(gate128inter4));
  nand2 gate1112(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1113(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1114(.a(G408), .O(gate128inter7));
  inv1  gate1115(.a(G409), .O(gate128inter8));
  nand2 gate1116(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1117(.a(s_81), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1118(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1119(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1120(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1485(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1486(.a(gate130inter0), .b(s_134), .O(gate130inter1));
  and2  gate1487(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1488(.a(s_134), .O(gate130inter3));
  inv1  gate1489(.a(s_135), .O(gate130inter4));
  nand2 gate1490(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1491(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1492(.a(G412), .O(gate130inter7));
  inv1  gate1493(.a(G413), .O(gate130inter8));
  nand2 gate1494(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1495(.a(s_135), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1496(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1497(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1498(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate771(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate772(.a(gate131inter0), .b(s_32), .O(gate131inter1));
  and2  gate773(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate774(.a(s_32), .O(gate131inter3));
  inv1  gate775(.a(s_33), .O(gate131inter4));
  nand2 gate776(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate777(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate778(.a(G414), .O(gate131inter7));
  inv1  gate779(.a(G415), .O(gate131inter8));
  nand2 gate780(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate781(.a(s_33), .b(gate131inter3), .O(gate131inter10));
  nor2  gate782(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate783(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate784(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate645(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate646(.a(gate132inter0), .b(s_14), .O(gate132inter1));
  and2  gate647(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate648(.a(s_14), .O(gate132inter3));
  inv1  gate649(.a(s_15), .O(gate132inter4));
  nand2 gate650(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate651(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate652(.a(G416), .O(gate132inter7));
  inv1  gate653(.a(G417), .O(gate132inter8));
  nand2 gate654(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate655(.a(s_15), .b(gate132inter3), .O(gate132inter10));
  nor2  gate656(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate657(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate658(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1793(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1794(.a(gate134inter0), .b(s_178), .O(gate134inter1));
  and2  gate1795(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1796(.a(s_178), .O(gate134inter3));
  inv1  gate1797(.a(s_179), .O(gate134inter4));
  nand2 gate1798(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1799(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1800(.a(G420), .O(gate134inter7));
  inv1  gate1801(.a(G421), .O(gate134inter8));
  nand2 gate1802(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1803(.a(s_179), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1804(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1805(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1806(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1569(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1570(.a(gate137inter0), .b(s_146), .O(gate137inter1));
  and2  gate1571(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1572(.a(s_146), .O(gate137inter3));
  inv1  gate1573(.a(s_147), .O(gate137inter4));
  nand2 gate1574(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1575(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1576(.a(G426), .O(gate137inter7));
  inv1  gate1577(.a(G429), .O(gate137inter8));
  nand2 gate1578(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1579(.a(s_147), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1580(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1581(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1582(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1639(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1640(.a(gate139inter0), .b(s_156), .O(gate139inter1));
  and2  gate1641(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1642(.a(s_156), .O(gate139inter3));
  inv1  gate1643(.a(s_157), .O(gate139inter4));
  nand2 gate1644(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1645(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1646(.a(G438), .O(gate139inter7));
  inv1  gate1647(.a(G441), .O(gate139inter8));
  nand2 gate1648(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1649(.a(s_157), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1650(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1651(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1652(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate995(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate996(.a(gate143inter0), .b(s_64), .O(gate143inter1));
  and2  gate997(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate998(.a(s_64), .O(gate143inter3));
  inv1  gate999(.a(s_65), .O(gate143inter4));
  nand2 gate1000(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1001(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1002(.a(G462), .O(gate143inter7));
  inv1  gate1003(.a(G465), .O(gate143inter8));
  nand2 gate1004(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1005(.a(s_65), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1006(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1007(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1008(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1373(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1374(.a(gate145inter0), .b(s_118), .O(gate145inter1));
  and2  gate1375(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1376(.a(s_118), .O(gate145inter3));
  inv1  gate1377(.a(s_119), .O(gate145inter4));
  nand2 gate1378(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1379(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1380(.a(G474), .O(gate145inter7));
  inv1  gate1381(.a(G477), .O(gate145inter8));
  nand2 gate1382(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1383(.a(s_119), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1384(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1385(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1386(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate855(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate856(.a(gate147inter0), .b(s_44), .O(gate147inter1));
  and2  gate857(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate858(.a(s_44), .O(gate147inter3));
  inv1  gate859(.a(s_45), .O(gate147inter4));
  nand2 gate860(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate861(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate862(.a(G486), .O(gate147inter7));
  inv1  gate863(.a(G489), .O(gate147inter8));
  nand2 gate864(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate865(.a(s_45), .b(gate147inter3), .O(gate147inter10));
  nor2  gate866(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate867(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate868(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1457(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1458(.a(gate148inter0), .b(s_130), .O(gate148inter1));
  and2  gate1459(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1460(.a(s_130), .O(gate148inter3));
  inv1  gate1461(.a(s_131), .O(gate148inter4));
  nand2 gate1462(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1463(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1464(.a(G492), .O(gate148inter7));
  inv1  gate1465(.a(G495), .O(gate148inter8));
  nand2 gate1466(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1467(.a(s_131), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1468(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1469(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1470(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate2367(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2368(.a(gate149inter0), .b(s_260), .O(gate149inter1));
  and2  gate2369(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2370(.a(s_260), .O(gate149inter3));
  inv1  gate2371(.a(s_261), .O(gate149inter4));
  nand2 gate2372(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2373(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2374(.a(G498), .O(gate149inter7));
  inv1  gate2375(.a(G501), .O(gate149inter8));
  nand2 gate2376(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2377(.a(s_261), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2378(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2379(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2380(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2311(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2312(.a(gate150inter0), .b(s_252), .O(gate150inter1));
  and2  gate2313(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2314(.a(s_252), .O(gate150inter3));
  inv1  gate2315(.a(s_253), .O(gate150inter4));
  nand2 gate2316(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2317(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2318(.a(G504), .O(gate150inter7));
  inv1  gate2319(.a(G507), .O(gate150inter8));
  nand2 gate2320(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2321(.a(s_253), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2322(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2323(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2324(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1205(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1206(.a(gate154inter0), .b(s_94), .O(gate154inter1));
  and2  gate1207(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1208(.a(s_94), .O(gate154inter3));
  inv1  gate1209(.a(s_95), .O(gate154inter4));
  nand2 gate1210(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1211(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1212(.a(G429), .O(gate154inter7));
  inv1  gate1213(.a(G522), .O(gate154inter8));
  nand2 gate1214(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1215(.a(s_95), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1216(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1217(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1218(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate757(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate758(.a(gate160inter0), .b(s_30), .O(gate160inter1));
  and2  gate759(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate760(.a(s_30), .O(gate160inter3));
  inv1  gate761(.a(s_31), .O(gate160inter4));
  nand2 gate762(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate763(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate764(.a(G447), .O(gate160inter7));
  inv1  gate765(.a(G531), .O(gate160inter8));
  nand2 gate766(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate767(.a(s_31), .b(gate160inter3), .O(gate160inter10));
  nor2  gate768(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate769(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate770(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate547(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate548(.a(gate163inter0), .b(s_0), .O(gate163inter1));
  and2  gate549(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate550(.a(s_0), .O(gate163inter3));
  inv1  gate551(.a(s_1), .O(gate163inter4));
  nand2 gate552(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate553(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate554(.a(G456), .O(gate163inter7));
  inv1  gate555(.a(G537), .O(gate163inter8));
  nand2 gate556(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate557(.a(s_1), .b(gate163inter3), .O(gate163inter10));
  nor2  gate558(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate559(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate560(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1065(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1066(.a(gate177inter0), .b(s_74), .O(gate177inter1));
  and2  gate1067(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1068(.a(s_74), .O(gate177inter3));
  inv1  gate1069(.a(s_75), .O(gate177inter4));
  nand2 gate1070(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1071(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1072(.a(G498), .O(gate177inter7));
  inv1  gate1073(.a(G558), .O(gate177inter8));
  nand2 gate1074(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1075(.a(s_75), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1076(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1077(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1078(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate897(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate898(.a(gate179inter0), .b(s_50), .O(gate179inter1));
  and2  gate899(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate900(.a(s_50), .O(gate179inter3));
  inv1  gate901(.a(s_51), .O(gate179inter4));
  nand2 gate902(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate903(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate904(.a(G504), .O(gate179inter7));
  inv1  gate905(.a(G561), .O(gate179inter8));
  nand2 gate906(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate907(.a(s_51), .b(gate179inter3), .O(gate179inter10));
  nor2  gate908(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate909(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate910(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1317(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1318(.a(gate182inter0), .b(s_110), .O(gate182inter1));
  and2  gate1319(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1320(.a(s_110), .O(gate182inter3));
  inv1  gate1321(.a(s_111), .O(gate182inter4));
  nand2 gate1322(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1323(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1324(.a(G513), .O(gate182inter7));
  inv1  gate1325(.a(G564), .O(gate182inter8));
  nand2 gate1326(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1327(.a(s_111), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1328(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1329(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1330(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1499(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1500(.a(gate185inter0), .b(s_136), .O(gate185inter1));
  and2  gate1501(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1502(.a(s_136), .O(gate185inter3));
  inv1  gate1503(.a(s_137), .O(gate185inter4));
  nand2 gate1504(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1505(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1506(.a(G570), .O(gate185inter7));
  inv1  gate1507(.a(G571), .O(gate185inter8));
  nand2 gate1508(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1509(.a(s_137), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1510(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1511(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1512(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1387(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1388(.a(gate186inter0), .b(s_120), .O(gate186inter1));
  and2  gate1389(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1390(.a(s_120), .O(gate186inter3));
  inv1  gate1391(.a(s_121), .O(gate186inter4));
  nand2 gate1392(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1393(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1394(.a(G572), .O(gate186inter7));
  inv1  gate1395(.a(G573), .O(gate186inter8));
  nand2 gate1396(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1397(.a(s_121), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1398(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1399(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1400(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1345(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1346(.a(gate194inter0), .b(s_114), .O(gate194inter1));
  and2  gate1347(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1348(.a(s_114), .O(gate194inter3));
  inv1  gate1349(.a(s_115), .O(gate194inter4));
  nand2 gate1350(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1351(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1352(.a(G588), .O(gate194inter7));
  inv1  gate1353(.a(G589), .O(gate194inter8));
  nand2 gate1354(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1355(.a(s_115), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1356(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1357(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1358(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1275(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1276(.a(gate196inter0), .b(s_104), .O(gate196inter1));
  and2  gate1277(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1278(.a(s_104), .O(gate196inter3));
  inv1  gate1279(.a(s_105), .O(gate196inter4));
  nand2 gate1280(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1281(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1282(.a(G592), .O(gate196inter7));
  inv1  gate1283(.a(G593), .O(gate196inter8));
  nand2 gate1284(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1285(.a(s_105), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1286(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1287(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1288(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2353(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2354(.a(gate200inter0), .b(s_258), .O(gate200inter1));
  and2  gate2355(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2356(.a(s_258), .O(gate200inter3));
  inv1  gate2357(.a(s_259), .O(gate200inter4));
  nand2 gate2358(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2359(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2360(.a(G600), .O(gate200inter7));
  inv1  gate2361(.a(G601), .O(gate200inter8));
  nand2 gate2362(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2363(.a(s_259), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2364(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2365(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2366(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1233(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1234(.a(gate205inter0), .b(s_98), .O(gate205inter1));
  and2  gate1235(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1236(.a(s_98), .O(gate205inter3));
  inv1  gate1237(.a(s_99), .O(gate205inter4));
  nand2 gate1238(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1239(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1240(.a(G622), .O(gate205inter7));
  inv1  gate1241(.a(G627), .O(gate205inter8));
  nand2 gate1242(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1243(.a(s_99), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1244(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1245(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1246(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1975(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1976(.a(gate208inter0), .b(s_204), .O(gate208inter1));
  and2  gate1977(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1978(.a(s_204), .O(gate208inter3));
  inv1  gate1979(.a(s_205), .O(gate208inter4));
  nand2 gate1980(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1981(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1982(.a(G627), .O(gate208inter7));
  inv1  gate1983(.a(G637), .O(gate208inter8));
  nand2 gate1984(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1985(.a(s_205), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1986(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1987(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1988(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1863(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1864(.a(gate209inter0), .b(s_188), .O(gate209inter1));
  and2  gate1865(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1866(.a(s_188), .O(gate209inter3));
  inv1  gate1867(.a(s_189), .O(gate209inter4));
  nand2 gate1868(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1869(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1870(.a(G602), .O(gate209inter7));
  inv1  gate1871(.a(G666), .O(gate209inter8));
  nand2 gate1872(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1873(.a(s_189), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1874(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1875(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1876(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1443(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1444(.a(gate210inter0), .b(s_128), .O(gate210inter1));
  and2  gate1445(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1446(.a(s_128), .O(gate210inter3));
  inv1  gate1447(.a(s_129), .O(gate210inter4));
  nand2 gate1448(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1449(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1450(.a(G607), .O(gate210inter7));
  inv1  gate1451(.a(G666), .O(gate210inter8));
  nand2 gate1452(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1453(.a(s_129), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1454(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1455(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1456(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate841(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate842(.a(gate211inter0), .b(s_42), .O(gate211inter1));
  and2  gate843(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate844(.a(s_42), .O(gate211inter3));
  inv1  gate845(.a(s_43), .O(gate211inter4));
  nand2 gate846(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate847(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate848(.a(G612), .O(gate211inter7));
  inv1  gate849(.a(G669), .O(gate211inter8));
  nand2 gate850(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate851(.a(s_43), .b(gate211inter3), .O(gate211inter10));
  nor2  gate852(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate853(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate854(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1737(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1738(.a(gate215inter0), .b(s_170), .O(gate215inter1));
  and2  gate1739(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1740(.a(s_170), .O(gate215inter3));
  inv1  gate1741(.a(s_171), .O(gate215inter4));
  nand2 gate1742(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1743(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1744(.a(G607), .O(gate215inter7));
  inv1  gate1745(.a(G675), .O(gate215inter8));
  nand2 gate1746(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1747(.a(s_171), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1748(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1749(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1750(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1303(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1304(.a(gate222inter0), .b(s_108), .O(gate222inter1));
  and2  gate1305(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1306(.a(s_108), .O(gate222inter3));
  inv1  gate1307(.a(s_109), .O(gate222inter4));
  nand2 gate1308(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1309(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1310(.a(G632), .O(gate222inter7));
  inv1  gate1311(.a(G684), .O(gate222inter8));
  nand2 gate1312(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1313(.a(s_109), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1314(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1315(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1316(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate715(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate716(.a(gate230inter0), .b(s_24), .O(gate230inter1));
  and2  gate717(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate718(.a(s_24), .O(gate230inter3));
  inv1  gate719(.a(s_25), .O(gate230inter4));
  nand2 gate720(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate721(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate722(.a(G700), .O(gate230inter7));
  inv1  gate723(.a(G701), .O(gate230inter8));
  nand2 gate724(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate725(.a(s_25), .b(gate230inter3), .O(gate230inter10));
  nor2  gate726(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate727(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate728(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1989(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1990(.a(gate234inter0), .b(s_206), .O(gate234inter1));
  and2  gate1991(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1992(.a(s_206), .O(gate234inter3));
  inv1  gate1993(.a(s_207), .O(gate234inter4));
  nand2 gate1994(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1995(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1996(.a(G245), .O(gate234inter7));
  inv1  gate1997(.a(G721), .O(gate234inter8));
  nand2 gate1998(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1999(.a(s_207), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2000(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2001(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2002(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2045(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2046(.a(gate236inter0), .b(s_214), .O(gate236inter1));
  and2  gate2047(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2048(.a(s_214), .O(gate236inter3));
  inv1  gate2049(.a(s_215), .O(gate236inter4));
  nand2 gate2050(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2051(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2052(.a(G251), .O(gate236inter7));
  inv1  gate2053(.a(G727), .O(gate236inter8));
  nand2 gate2054(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2055(.a(s_215), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2056(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2057(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2058(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate617(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate618(.a(gate237inter0), .b(s_10), .O(gate237inter1));
  and2  gate619(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate620(.a(s_10), .O(gate237inter3));
  inv1  gate621(.a(s_11), .O(gate237inter4));
  nand2 gate622(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate623(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate624(.a(G254), .O(gate237inter7));
  inv1  gate625(.a(G706), .O(gate237inter8));
  nand2 gate626(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate627(.a(s_11), .b(gate237inter3), .O(gate237inter10));
  nor2  gate628(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate629(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate630(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1163(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1164(.a(gate248inter0), .b(s_88), .O(gate248inter1));
  and2  gate1165(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1166(.a(s_88), .O(gate248inter3));
  inv1  gate1167(.a(s_89), .O(gate248inter4));
  nand2 gate1168(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1169(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1170(.a(G727), .O(gate248inter7));
  inv1  gate1171(.a(G739), .O(gate248inter8));
  nand2 gate1172(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1173(.a(s_89), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1174(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1175(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1176(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1625(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1626(.a(gate252inter0), .b(s_154), .O(gate252inter1));
  and2  gate1627(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1628(.a(s_154), .O(gate252inter3));
  inv1  gate1629(.a(s_155), .O(gate252inter4));
  nand2 gate1630(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1631(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1632(.a(G709), .O(gate252inter7));
  inv1  gate1633(.a(G745), .O(gate252inter8));
  nand2 gate1634(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1635(.a(s_155), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1636(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1637(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1638(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate925(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate926(.a(gate253inter0), .b(s_54), .O(gate253inter1));
  and2  gate927(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate928(.a(s_54), .O(gate253inter3));
  inv1  gate929(.a(s_55), .O(gate253inter4));
  nand2 gate930(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate931(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate932(.a(G260), .O(gate253inter7));
  inv1  gate933(.a(G748), .O(gate253inter8));
  nand2 gate934(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate935(.a(s_55), .b(gate253inter3), .O(gate253inter10));
  nor2  gate936(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate937(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate938(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1653(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1654(.a(gate256inter0), .b(s_158), .O(gate256inter1));
  and2  gate1655(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1656(.a(s_158), .O(gate256inter3));
  inv1  gate1657(.a(s_159), .O(gate256inter4));
  nand2 gate1658(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1659(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1660(.a(G715), .O(gate256inter7));
  inv1  gate1661(.a(G751), .O(gate256inter8));
  nand2 gate1662(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1663(.a(s_159), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1664(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1665(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1666(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1849(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1850(.a(gate257inter0), .b(s_186), .O(gate257inter1));
  and2  gate1851(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1852(.a(s_186), .O(gate257inter3));
  inv1  gate1853(.a(s_187), .O(gate257inter4));
  nand2 gate1854(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1855(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1856(.a(G754), .O(gate257inter7));
  inv1  gate1857(.a(G755), .O(gate257inter8));
  nand2 gate1858(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1859(.a(s_187), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1860(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1861(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1862(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1331(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1332(.a(gate260inter0), .b(s_112), .O(gate260inter1));
  and2  gate1333(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1334(.a(s_112), .O(gate260inter3));
  inv1  gate1335(.a(s_113), .O(gate260inter4));
  nand2 gate1336(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1337(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1338(.a(G760), .O(gate260inter7));
  inv1  gate1339(.a(G761), .O(gate260inter8));
  nand2 gate1340(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1341(.a(s_113), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1342(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1343(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1344(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1191(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1192(.a(gate263inter0), .b(s_92), .O(gate263inter1));
  and2  gate1193(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1194(.a(s_92), .O(gate263inter3));
  inv1  gate1195(.a(s_93), .O(gate263inter4));
  nand2 gate1196(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1197(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1198(.a(G766), .O(gate263inter7));
  inv1  gate1199(.a(G767), .O(gate263inter8));
  nand2 gate1200(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1201(.a(s_93), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1202(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1203(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1204(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2129(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2130(.a(gate265inter0), .b(s_226), .O(gate265inter1));
  and2  gate2131(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2132(.a(s_226), .O(gate265inter3));
  inv1  gate2133(.a(s_227), .O(gate265inter4));
  nand2 gate2134(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2135(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2136(.a(G642), .O(gate265inter7));
  inv1  gate2137(.a(G770), .O(gate265inter8));
  nand2 gate2138(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2139(.a(s_227), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2140(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2141(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2142(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1261(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1262(.a(gate268inter0), .b(s_102), .O(gate268inter1));
  and2  gate1263(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1264(.a(s_102), .O(gate268inter3));
  inv1  gate1265(.a(s_103), .O(gate268inter4));
  nand2 gate1266(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1267(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1268(.a(G651), .O(gate268inter7));
  inv1  gate1269(.a(G779), .O(gate268inter8));
  nand2 gate1270(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1271(.a(s_103), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1272(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1273(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1274(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1681(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1682(.a(gate269inter0), .b(s_162), .O(gate269inter1));
  and2  gate1683(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1684(.a(s_162), .O(gate269inter3));
  inv1  gate1685(.a(s_163), .O(gate269inter4));
  nand2 gate1686(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1687(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1688(.a(G654), .O(gate269inter7));
  inv1  gate1689(.a(G782), .O(gate269inter8));
  nand2 gate1690(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1691(.a(s_163), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1692(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1693(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1694(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate1723(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1724(.a(gate270inter0), .b(s_168), .O(gate270inter1));
  and2  gate1725(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1726(.a(s_168), .O(gate270inter3));
  inv1  gate1727(.a(s_169), .O(gate270inter4));
  nand2 gate1728(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1729(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1730(.a(G657), .O(gate270inter7));
  inv1  gate1731(.a(G785), .O(gate270inter8));
  nand2 gate1732(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1733(.a(s_169), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1734(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1735(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1736(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1695(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1696(.a(gate280inter0), .b(s_164), .O(gate280inter1));
  and2  gate1697(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1698(.a(s_164), .O(gate280inter3));
  inv1  gate1699(.a(s_165), .O(gate280inter4));
  nand2 gate1700(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1701(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1702(.a(G779), .O(gate280inter7));
  inv1  gate1703(.a(G803), .O(gate280inter8));
  nand2 gate1704(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1705(.a(s_165), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1706(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1707(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1708(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1583(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1584(.a(gate281inter0), .b(s_148), .O(gate281inter1));
  and2  gate1585(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1586(.a(s_148), .O(gate281inter3));
  inv1  gate1587(.a(s_149), .O(gate281inter4));
  nand2 gate1588(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1589(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1590(.a(G654), .O(gate281inter7));
  inv1  gate1591(.a(G806), .O(gate281inter8));
  nand2 gate1592(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1593(.a(s_149), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1594(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1595(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1596(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate967(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate968(.a(gate287inter0), .b(s_60), .O(gate287inter1));
  and2  gate969(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate970(.a(s_60), .O(gate287inter3));
  inv1  gate971(.a(s_61), .O(gate287inter4));
  nand2 gate972(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate973(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate974(.a(G663), .O(gate287inter7));
  inv1  gate975(.a(G815), .O(gate287inter8));
  nand2 gate976(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate977(.a(s_61), .b(gate287inter3), .O(gate287inter10));
  nor2  gate978(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate979(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate980(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2017(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2018(.a(gate291inter0), .b(s_210), .O(gate291inter1));
  and2  gate2019(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2020(.a(s_210), .O(gate291inter3));
  inv1  gate2021(.a(s_211), .O(gate291inter4));
  nand2 gate2022(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2023(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2024(.a(G822), .O(gate291inter7));
  inv1  gate2025(.a(G823), .O(gate291inter8));
  nand2 gate2026(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2027(.a(s_211), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2028(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2029(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2030(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1891(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1892(.a(gate292inter0), .b(s_192), .O(gate292inter1));
  and2  gate1893(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1894(.a(s_192), .O(gate292inter3));
  inv1  gate1895(.a(s_193), .O(gate292inter4));
  nand2 gate1896(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1897(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1898(.a(G824), .O(gate292inter7));
  inv1  gate1899(.a(G825), .O(gate292inter8));
  nand2 gate1900(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1901(.a(s_193), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1902(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1903(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1904(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1541(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1542(.a(gate294inter0), .b(s_142), .O(gate294inter1));
  and2  gate1543(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1544(.a(s_142), .O(gate294inter3));
  inv1  gate1545(.a(s_143), .O(gate294inter4));
  nand2 gate1546(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1547(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1548(.a(G832), .O(gate294inter7));
  inv1  gate1549(.a(G833), .O(gate294inter8));
  nand2 gate1550(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1551(.a(s_143), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1552(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1553(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1554(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1807(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1808(.a(gate296inter0), .b(s_180), .O(gate296inter1));
  and2  gate1809(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1810(.a(s_180), .O(gate296inter3));
  inv1  gate1811(.a(s_181), .O(gate296inter4));
  nand2 gate1812(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1813(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1814(.a(G826), .O(gate296inter7));
  inv1  gate1815(.a(G827), .O(gate296inter8));
  nand2 gate1816(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1817(.a(s_181), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1818(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1819(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1820(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1765(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1766(.a(gate388inter0), .b(s_174), .O(gate388inter1));
  and2  gate1767(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1768(.a(s_174), .O(gate388inter3));
  inv1  gate1769(.a(s_175), .O(gate388inter4));
  nand2 gate1770(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1771(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1772(.a(G2), .O(gate388inter7));
  inv1  gate1773(.a(G1039), .O(gate388inter8));
  nand2 gate1774(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1775(.a(s_175), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1776(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1777(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1778(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate869(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate870(.a(gate389inter0), .b(s_46), .O(gate389inter1));
  and2  gate871(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate872(.a(s_46), .O(gate389inter3));
  inv1  gate873(.a(s_47), .O(gate389inter4));
  nand2 gate874(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate875(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate876(.a(G3), .O(gate389inter7));
  inv1  gate877(.a(G1042), .O(gate389inter8));
  nand2 gate878(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate879(.a(s_47), .b(gate389inter3), .O(gate389inter10));
  nor2  gate880(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate881(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate882(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate2059(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2060(.a(gate390inter0), .b(s_216), .O(gate390inter1));
  and2  gate2061(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2062(.a(s_216), .O(gate390inter3));
  inv1  gate2063(.a(s_217), .O(gate390inter4));
  nand2 gate2064(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2065(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2066(.a(G4), .O(gate390inter7));
  inv1  gate2067(.a(G1045), .O(gate390inter8));
  nand2 gate2068(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2069(.a(s_217), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2070(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2071(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2072(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2073(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2074(.a(gate396inter0), .b(s_218), .O(gate396inter1));
  and2  gate2075(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2076(.a(s_218), .O(gate396inter3));
  inv1  gate2077(.a(s_219), .O(gate396inter4));
  nand2 gate2078(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2079(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2080(.a(G10), .O(gate396inter7));
  inv1  gate2081(.a(G1063), .O(gate396inter8));
  nand2 gate2082(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2083(.a(s_219), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2084(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2085(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2086(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1121(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1122(.a(gate406inter0), .b(s_82), .O(gate406inter1));
  and2  gate1123(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1124(.a(s_82), .O(gate406inter3));
  inv1  gate1125(.a(s_83), .O(gate406inter4));
  nand2 gate1126(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1127(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1128(.a(G20), .O(gate406inter7));
  inv1  gate1129(.a(G1093), .O(gate406inter8));
  nand2 gate1130(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1131(.a(s_83), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1132(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1133(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1134(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1415(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1416(.a(gate408inter0), .b(s_124), .O(gate408inter1));
  and2  gate1417(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1418(.a(s_124), .O(gate408inter3));
  inv1  gate1419(.a(s_125), .O(gate408inter4));
  nand2 gate1420(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1421(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1422(.a(G22), .O(gate408inter7));
  inv1  gate1423(.a(G1099), .O(gate408inter8));
  nand2 gate1424(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1425(.a(s_125), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1426(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1427(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1428(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1905(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1906(.a(gate409inter0), .b(s_194), .O(gate409inter1));
  and2  gate1907(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1908(.a(s_194), .O(gate409inter3));
  inv1  gate1909(.a(s_195), .O(gate409inter4));
  nand2 gate1910(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1911(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1912(.a(G23), .O(gate409inter7));
  inv1  gate1913(.a(G1102), .O(gate409inter8));
  nand2 gate1914(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1915(.a(s_195), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1916(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1917(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1918(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1667(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1668(.a(gate411inter0), .b(s_160), .O(gate411inter1));
  and2  gate1669(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1670(.a(s_160), .O(gate411inter3));
  inv1  gate1671(.a(s_161), .O(gate411inter4));
  nand2 gate1672(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1673(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1674(.a(G25), .O(gate411inter7));
  inv1  gate1675(.a(G1108), .O(gate411inter8));
  nand2 gate1676(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1677(.a(s_161), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1678(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1679(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1680(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2003(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2004(.a(gate416inter0), .b(s_208), .O(gate416inter1));
  and2  gate2005(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2006(.a(s_208), .O(gate416inter3));
  inv1  gate2007(.a(s_209), .O(gate416inter4));
  nand2 gate2008(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2009(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2010(.a(G30), .O(gate416inter7));
  inv1  gate2011(.a(G1123), .O(gate416inter8));
  nand2 gate2012(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2013(.a(s_209), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2014(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2015(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2016(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1877(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1878(.a(gate418inter0), .b(s_190), .O(gate418inter1));
  and2  gate1879(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1880(.a(s_190), .O(gate418inter3));
  inv1  gate1881(.a(s_191), .O(gate418inter4));
  nand2 gate1882(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1883(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1884(.a(G32), .O(gate418inter7));
  inv1  gate1885(.a(G1129), .O(gate418inter8));
  nand2 gate1886(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1887(.a(s_191), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1888(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1889(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1890(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate939(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate940(.a(gate422inter0), .b(s_56), .O(gate422inter1));
  and2  gate941(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate942(.a(s_56), .O(gate422inter3));
  inv1  gate943(.a(s_57), .O(gate422inter4));
  nand2 gate944(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate945(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate946(.a(G1039), .O(gate422inter7));
  inv1  gate947(.a(G1135), .O(gate422inter8));
  nand2 gate948(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate949(.a(s_57), .b(gate422inter3), .O(gate422inter10));
  nor2  gate950(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate951(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate952(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2339(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2340(.a(gate428inter0), .b(s_256), .O(gate428inter1));
  and2  gate2341(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2342(.a(s_256), .O(gate428inter3));
  inv1  gate2343(.a(s_257), .O(gate428inter4));
  nand2 gate2344(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2345(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2346(.a(G1048), .O(gate428inter7));
  inv1  gate2347(.a(G1144), .O(gate428inter8));
  nand2 gate2348(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2349(.a(s_257), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2350(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2351(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2352(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2199(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2200(.a(gate430inter0), .b(s_236), .O(gate430inter1));
  and2  gate2201(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2202(.a(s_236), .O(gate430inter3));
  inv1  gate2203(.a(s_237), .O(gate430inter4));
  nand2 gate2204(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2205(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2206(.a(G1051), .O(gate430inter7));
  inv1  gate2207(.a(G1147), .O(gate430inter8));
  nand2 gate2208(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2209(.a(s_237), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2210(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2211(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2212(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate785(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate786(.a(gate434inter0), .b(s_34), .O(gate434inter1));
  and2  gate787(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate788(.a(s_34), .O(gate434inter3));
  inv1  gate789(.a(s_35), .O(gate434inter4));
  nand2 gate790(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate791(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate792(.a(G1057), .O(gate434inter7));
  inv1  gate793(.a(G1153), .O(gate434inter8));
  nand2 gate794(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate795(.a(s_35), .b(gate434inter3), .O(gate434inter10));
  nor2  gate796(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate797(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate798(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2297(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2298(.a(gate439inter0), .b(s_250), .O(gate439inter1));
  and2  gate2299(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2300(.a(s_250), .O(gate439inter3));
  inv1  gate2301(.a(s_251), .O(gate439inter4));
  nand2 gate2302(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2303(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2304(.a(G11), .O(gate439inter7));
  inv1  gate2305(.a(G1162), .O(gate439inter8));
  nand2 gate2306(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2307(.a(s_251), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2308(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2309(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2310(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate729(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate730(.a(gate443inter0), .b(s_26), .O(gate443inter1));
  and2  gate731(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate732(.a(s_26), .O(gate443inter3));
  inv1  gate733(.a(s_27), .O(gate443inter4));
  nand2 gate734(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate735(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate736(.a(G13), .O(gate443inter7));
  inv1  gate737(.a(G1168), .O(gate443inter8));
  nand2 gate738(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate739(.a(s_27), .b(gate443inter3), .O(gate443inter10));
  nor2  gate740(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate741(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate742(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1079(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1080(.a(gate447inter0), .b(s_76), .O(gate447inter1));
  and2  gate1081(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1082(.a(s_76), .O(gate447inter3));
  inv1  gate1083(.a(s_77), .O(gate447inter4));
  nand2 gate1084(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1085(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1086(.a(G15), .O(gate447inter7));
  inv1  gate1087(.a(G1174), .O(gate447inter8));
  nand2 gate1088(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1089(.a(s_77), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1090(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1091(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1092(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2255(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2256(.a(gate448inter0), .b(s_244), .O(gate448inter1));
  and2  gate2257(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2258(.a(s_244), .O(gate448inter3));
  inv1  gate2259(.a(s_245), .O(gate448inter4));
  nand2 gate2260(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2261(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2262(.a(G1078), .O(gate448inter7));
  inv1  gate2263(.a(G1174), .O(gate448inter8));
  nand2 gate2264(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2265(.a(s_245), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2266(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2267(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2268(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2171(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2172(.a(gate449inter0), .b(s_232), .O(gate449inter1));
  and2  gate2173(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2174(.a(s_232), .O(gate449inter3));
  inv1  gate2175(.a(s_233), .O(gate449inter4));
  nand2 gate2176(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2177(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2178(.a(G16), .O(gate449inter7));
  inv1  gate2179(.a(G1177), .O(gate449inter8));
  nand2 gate2180(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2181(.a(s_233), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2182(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2183(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2184(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2087(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2088(.a(gate458inter0), .b(s_220), .O(gate458inter1));
  and2  gate2089(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2090(.a(s_220), .O(gate458inter3));
  inv1  gate2091(.a(s_221), .O(gate458inter4));
  nand2 gate2092(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2093(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2094(.a(G1093), .O(gate458inter7));
  inv1  gate2095(.a(G1189), .O(gate458inter8));
  nand2 gate2096(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2097(.a(s_221), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2098(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2099(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2100(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate813(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate814(.a(gate467inter0), .b(s_38), .O(gate467inter1));
  and2  gate815(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate816(.a(s_38), .O(gate467inter3));
  inv1  gate817(.a(s_39), .O(gate467inter4));
  nand2 gate818(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate819(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate820(.a(G25), .O(gate467inter7));
  inv1  gate821(.a(G1204), .O(gate467inter8));
  nand2 gate822(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate823(.a(s_39), .b(gate467inter3), .O(gate467inter10));
  nor2  gate824(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate825(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate826(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate2269(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2270(.a(gate468inter0), .b(s_246), .O(gate468inter1));
  and2  gate2271(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2272(.a(s_246), .O(gate468inter3));
  inv1  gate2273(.a(s_247), .O(gate468inter4));
  nand2 gate2274(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2275(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2276(.a(G1108), .O(gate468inter7));
  inv1  gate2277(.a(G1204), .O(gate468inter8));
  nand2 gate2278(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2279(.a(s_247), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2280(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2281(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2282(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2157(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2158(.a(gate474inter0), .b(s_230), .O(gate474inter1));
  and2  gate2159(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2160(.a(s_230), .O(gate474inter3));
  inv1  gate2161(.a(s_231), .O(gate474inter4));
  nand2 gate2162(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2163(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2164(.a(G1117), .O(gate474inter7));
  inv1  gate2165(.a(G1213), .O(gate474inter8));
  nand2 gate2166(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2167(.a(s_231), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2168(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2169(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2170(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate659(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate660(.a(gate476inter0), .b(s_16), .O(gate476inter1));
  and2  gate661(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate662(.a(s_16), .O(gate476inter3));
  inv1  gate663(.a(s_17), .O(gate476inter4));
  nand2 gate664(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate665(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate666(.a(G1120), .O(gate476inter7));
  inv1  gate667(.a(G1216), .O(gate476inter8));
  nand2 gate668(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate669(.a(s_17), .b(gate476inter3), .O(gate476inter10));
  nor2  gate670(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate671(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate672(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2325(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2326(.a(gate478inter0), .b(s_254), .O(gate478inter1));
  and2  gate2327(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2328(.a(s_254), .O(gate478inter3));
  inv1  gate2329(.a(s_255), .O(gate478inter4));
  nand2 gate2330(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2331(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2332(.a(G1123), .O(gate478inter7));
  inv1  gate2333(.a(G1219), .O(gate478inter8));
  nand2 gate2334(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2335(.a(s_255), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2336(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2337(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2338(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1961(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1962(.a(gate480inter0), .b(s_202), .O(gate480inter1));
  and2  gate1963(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1964(.a(s_202), .O(gate480inter3));
  inv1  gate1965(.a(s_203), .O(gate480inter4));
  nand2 gate1966(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1967(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1968(.a(G1126), .O(gate480inter7));
  inv1  gate1969(.a(G1222), .O(gate480inter8));
  nand2 gate1970(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1971(.a(s_203), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1972(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1973(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1974(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1177(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1178(.a(gate484inter0), .b(s_90), .O(gate484inter1));
  and2  gate1179(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1180(.a(s_90), .O(gate484inter3));
  inv1  gate1181(.a(s_91), .O(gate484inter4));
  nand2 gate1182(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1183(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1184(.a(G1230), .O(gate484inter7));
  inv1  gate1185(.a(G1231), .O(gate484inter8));
  nand2 gate1186(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1187(.a(s_91), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1188(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1189(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1190(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1835(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1836(.a(gate485inter0), .b(s_184), .O(gate485inter1));
  and2  gate1837(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1838(.a(s_184), .O(gate485inter3));
  inv1  gate1839(.a(s_185), .O(gate485inter4));
  nand2 gate1840(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1841(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1842(.a(G1232), .O(gate485inter7));
  inv1  gate1843(.a(G1233), .O(gate485inter8));
  nand2 gate1844(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1845(.a(s_185), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1846(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1847(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1848(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate701(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate702(.a(gate488inter0), .b(s_22), .O(gate488inter1));
  and2  gate703(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate704(.a(s_22), .O(gate488inter3));
  inv1  gate705(.a(s_23), .O(gate488inter4));
  nand2 gate706(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate707(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate708(.a(G1238), .O(gate488inter7));
  inv1  gate709(.a(G1239), .O(gate488inter8));
  nand2 gate710(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate711(.a(s_23), .b(gate488inter3), .O(gate488inter10));
  nor2  gate712(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate713(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate714(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1037(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1038(.a(gate496inter0), .b(s_70), .O(gate496inter1));
  and2  gate1039(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1040(.a(s_70), .O(gate496inter3));
  inv1  gate1041(.a(s_71), .O(gate496inter4));
  nand2 gate1042(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1043(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1044(.a(G1254), .O(gate496inter7));
  inv1  gate1045(.a(G1255), .O(gate496inter8));
  nand2 gate1046(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1047(.a(s_71), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1048(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1049(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1050(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate687(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate688(.a(gate497inter0), .b(s_20), .O(gate497inter1));
  and2  gate689(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate690(.a(s_20), .O(gate497inter3));
  inv1  gate691(.a(s_21), .O(gate497inter4));
  nand2 gate692(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate693(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate694(.a(G1256), .O(gate497inter7));
  inv1  gate695(.a(G1257), .O(gate497inter8));
  nand2 gate696(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate697(.a(s_21), .b(gate497inter3), .O(gate497inter10));
  nor2  gate698(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate699(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate700(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1149(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1150(.a(gate498inter0), .b(s_86), .O(gate498inter1));
  and2  gate1151(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1152(.a(s_86), .O(gate498inter3));
  inv1  gate1153(.a(s_87), .O(gate498inter4));
  nand2 gate1154(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1155(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1156(.a(G1258), .O(gate498inter7));
  inv1  gate1157(.a(G1259), .O(gate498inter8));
  nand2 gate1158(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1159(.a(s_87), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1160(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1161(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1162(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate673(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate674(.a(gate499inter0), .b(s_18), .O(gate499inter1));
  and2  gate675(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate676(.a(s_18), .O(gate499inter3));
  inv1  gate677(.a(s_19), .O(gate499inter4));
  nand2 gate678(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate679(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate680(.a(G1260), .O(gate499inter7));
  inv1  gate681(.a(G1261), .O(gate499inter8));
  nand2 gate682(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate683(.a(s_19), .b(gate499inter3), .O(gate499inter10));
  nor2  gate684(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate685(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate686(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1611(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1612(.a(gate503inter0), .b(s_152), .O(gate503inter1));
  and2  gate1613(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1614(.a(s_152), .O(gate503inter3));
  inv1  gate1615(.a(s_153), .O(gate503inter4));
  nand2 gate1616(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1617(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1618(.a(G1268), .O(gate503inter7));
  inv1  gate1619(.a(G1269), .O(gate503inter8));
  nand2 gate1620(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1621(.a(s_153), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1622(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1623(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1624(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1821(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1822(.a(gate510inter0), .b(s_182), .O(gate510inter1));
  and2  gate1823(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1824(.a(s_182), .O(gate510inter3));
  inv1  gate1825(.a(s_183), .O(gate510inter4));
  nand2 gate1826(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1827(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1828(.a(G1282), .O(gate510inter7));
  inv1  gate1829(.a(G1283), .O(gate510inter8));
  nand2 gate1830(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1831(.a(s_183), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1832(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1833(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1834(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule