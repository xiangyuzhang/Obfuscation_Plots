module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1261(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1262(.a(gate19inter0), .b(s_102), .O(gate19inter1));
  and2  gate1263(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1264(.a(s_102), .O(gate19inter3));
  inv1  gate1265(.a(s_103), .O(gate19inter4));
  nand2 gate1266(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1267(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1268(.a(G21), .O(gate19inter7));
  inv1  gate1269(.a(G22), .O(gate19inter8));
  nand2 gate1270(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1271(.a(s_103), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1272(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1273(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1274(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1723(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1724(.a(gate23inter0), .b(s_168), .O(gate23inter1));
  and2  gate1725(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1726(.a(s_168), .O(gate23inter3));
  inv1  gate1727(.a(s_169), .O(gate23inter4));
  nand2 gate1728(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1729(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1730(.a(G29), .O(gate23inter7));
  inv1  gate1731(.a(G30), .O(gate23inter8));
  nand2 gate1732(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1733(.a(s_169), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1734(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1735(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1736(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1611(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1612(.a(gate24inter0), .b(s_152), .O(gate24inter1));
  and2  gate1613(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1614(.a(s_152), .O(gate24inter3));
  inv1  gate1615(.a(s_153), .O(gate24inter4));
  nand2 gate1616(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1617(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1618(.a(G31), .O(gate24inter7));
  inv1  gate1619(.a(G32), .O(gate24inter8));
  nand2 gate1620(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1621(.a(s_153), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1622(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1623(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1624(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1177(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1178(.a(gate28inter0), .b(s_90), .O(gate28inter1));
  and2  gate1179(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1180(.a(s_90), .O(gate28inter3));
  inv1  gate1181(.a(s_91), .O(gate28inter4));
  nand2 gate1182(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1183(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1184(.a(G10), .O(gate28inter7));
  inv1  gate1185(.a(G14), .O(gate28inter8));
  nand2 gate1186(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1187(.a(s_91), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1188(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1189(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1190(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate673(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate674(.a(gate29inter0), .b(s_18), .O(gate29inter1));
  and2  gate675(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate676(.a(s_18), .O(gate29inter3));
  inv1  gate677(.a(s_19), .O(gate29inter4));
  nand2 gate678(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate679(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate680(.a(G3), .O(gate29inter7));
  inv1  gate681(.a(G7), .O(gate29inter8));
  nand2 gate682(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate683(.a(s_19), .b(gate29inter3), .O(gate29inter10));
  nor2  gate684(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate685(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate686(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1387(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1388(.a(gate32inter0), .b(s_120), .O(gate32inter1));
  and2  gate1389(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1390(.a(s_120), .O(gate32inter3));
  inv1  gate1391(.a(s_121), .O(gate32inter4));
  nand2 gate1392(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1393(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1394(.a(G12), .O(gate32inter7));
  inv1  gate1395(.a(G16), .O(gate32inter8));
  nand2 gate1396(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1397(.a(s_121), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1398(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1399(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1400(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1023(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1024(.a(gate36inter0), .b(s_68), .O(gate36inter1));
  and2  gate1025(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1026(.a(s_68), .O(gate36inter3));
  inv1  gate1027(.a(s_69), .O(gate36inter4));
  nand2 gate1028(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1029(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1030(.a(G26), .O(gate36inter7));
  inv1  gate1031(.a(G30), .O(gate36inter8));
  nand2 gate1032(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1033(.a(s_69), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1034(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1035(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1036(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1149(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1150(.a(gate42inter0), .b(s_86), .O(gate42inter1));
  and2  gate1151(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1152(.a(s_86), .O(gate42inter3));
  inv1  gate1153(.a(s_87), .O(gate42inter4));
  nand2 gate1154(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1155(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1156(.a(G2), .O(gate42inter7));
  inv1  gate1157(.a(G266), .O(gate42inter8));
  nand2 gate1158(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1159(.a(s_87), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1160(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1161(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1162(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate561(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate562(.a(gate47inter0), .b(s_2), .O(gate47inter1));
  and2  gate563(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate564(.a(s_2), .O(gate47inter3));
  inv1  gate565(.a(s_3), .O(gate47inter4));
  nand2 gate566(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate567(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate568(.a(G7), .O(gate47inter7));
  inv1  gate569(.a(G275), .O(gate47inter8));
  nand2 gate570(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate571(.a(s_3), .b(gate47inter3), .O(gate47inter10));
  nor2  gate572(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate573(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate574(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1065(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1066(.a(gate50inter0), .b(s_74), .O(gate50inter1));
  and2  gate1067(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1068(.a(s_74), .O(gate50inter3));
  inv1  gate1069(.a(s_75), .O(gate50inter4));
  nand2 gate1070(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1071(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1072(.a(G10), .O(gate50inter7));
  inv1  gate1073(.a(G278), .O(gate50inter8));
  nand2 gate1074(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1075(.a(s_75), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1076(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1077(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1078(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate855(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate856(.a(gate53inter0), .b(s_44), .O(gate53inter1));
  and2  gate857(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate858(.a(s_44), .O(gate53inter3));
  inv1  gate859(.a(s_45), .O(gate53inter4));
  nand2 gate860(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate861(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate862(.a(G13), .O(gate53inter7));
  inv1  gate863(.a(G284), .O(gate53inter8));
  nand2 gate864(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate865(.a(s_45), .b(gate53inter3), .O(gate53inter10));
  nor2  gate866(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate867(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate868(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1051(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1052(.a(gate57inter0), .b(s_72), .O(gate57inter1));
  and2  gate1053(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1054(.a(s_72), .O(gate57inter3));
  inv1  gate1055(.a(s_73), .O(gate57inter4));
  nand2 gate1056(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1057(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1058(.a(G17), .O(gate57inter7));
  inv1  gate1059(.a(G290), .O(gate57inter8));
  nand2 gate1060(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1061(.a(s_73), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1062(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1063(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1064(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1709(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1710(.a(gate62inter0), .b(s_166), .O(gate62inter1));
  and2  gate1711(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1712(.a(s_166), .O(gate62inter3));
  inv1  gate1713(.a(s_167), .O(gate62inter4));
  nand2 gate1714(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1715(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1716(.a(G22), .O(gate62inter7));
  inv1  gate1717(.a(G296), .O(gate62inter8));
  nand2 gate1718(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1719(.a(s_167), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1720(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1721(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1722(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate659(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate660(.a(gate66inter0), .b(s_16), .O(gate66inter1));
  and2  gate661(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate662(.a(s_16), .O(gate66inter3));
  inv1  gate663(.a(s_17), .O(gate66inter4));
  nand2 gate664(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate665(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate666(.a(G26), .O(gate66inter7));
  inv1  gate667(.a(G302), .O(gate66inter8));
  nand2 gate668(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate669(.a(s_17), .b(gate66inter3), .O(gate66inter10));
  nor2  gate670(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate671(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate672(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1429(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1430(.a(gate68inter0), .b(s_126), .O(gate68inter1));
  and2  gate1431(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1432(.a(s_126), .O(gate68inter3));
  inv1  gate1433(.a(s_127), .O(gate68inter4));
  nand2 gate1434(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1435(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1436(.a(G28), .O(gate68inter7));
  inv1  gate1437(.a(G305), .O(gate68inter8));
  nand2 gate1438(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1439(.a(s_127), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1440(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1441(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1442(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate771(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate772(.a(gate73inter0), .b(s_32), .O(gate73inter1));
  and2  gate773(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate774(.a(s_32), .O(gate73inter3));
  inv1  gate775(.a(s_33), .O(gate73inter4));
  nand2 gate776(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate777(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate778(.a(G1), .O(gate73inter7));
  inv1  gate779(.a(G314), .O(gate73inter8));
  nand2 gate780(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate781(.a(s_33), .b(gate73inter3), .O(gate73inter10));
  nor2  gate782(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate783(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate784(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1807(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1808(.a(gate76inter0), .b(s_180), .O(gate76inter1));
  and2  gate1809(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1810(.a(s_180), .O(gate76inter3));
  inv1  gate1811(.a(s_181), .O(gate76inter4));
  nand2 gate1812(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1813(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1814(.a(G13), .O(gate76inter7));
  inv1  gate1815(.a(G317), .O(gate76inter8));
  nand2 gate1816(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1817(.a(s_181), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1818(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1819(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1820(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1583(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1584(.a(gate77inter0), .b(s_148), .O(gate77inter1));
  and2  gate1585(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1586(.a(s_148), .O(gate77inter3));
  inv1  gate1587(.a(s_149), .O(gate77inter4));
  nand2 gate1588(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1589(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1590(.a(G2), .O(gate77inter7));
  inv1  gate1591(.a(G320), .O(gate77inter8));
  nand2 gate1592(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1593(.a(s_149), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1594(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1595(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1596(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1009(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1010(.a(gate79inter0), .b(s_66), .O(gate79inter1));
  and2  gate1011(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1012(.a(s_66), .O(gate79inter3));
  inv1  gate1013(.a(s_67), .O(gate79inter4));
  nand2 gate1014(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1015(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1016(.a(G10), .O(gate79inter7));
  inv1  gate1017(.a(G323), .O(gate79inter8));
  nand2 gate1018(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1019(.a(s_67), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1020(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1021(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1022(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1877(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1878(.a(gate85inter0), .b(s_190), .O(gate85inter1));
  and2  gate1879(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1880(.a(s_190), .O(gate85inter3));
  inv1  gate1881(.a(s_191), .O(gate85inter4));
  nand2 gate1882(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1883(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1884(.a(G4), .O(gate85inter7));
  inv1  gate1885(.a(G332), .O(gate85inter8));
  nand2 gate1886(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1887(.a(s_191), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1888(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1889(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1890(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate925(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate926(.a(gate88inter0), .b(s_54), .O(gate88inter1));
  and2  gate927(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate928(.a(s_54), .O(gate88inter3));
  inv1  gate929(.a(s_55), .O(gate88inter4));
  nand2 gate930(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate931(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate932(.a(G16), .O(gate88inter7));
  inv1  gate933(.a(G335), .O(gate88inter8));
  nand2 gate934(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate935(.a(s_55), .b(gate88inter3), .O(gate88inter10));
  nor2  gate936(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate937(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate938(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate939(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate940(.a(gate94inter0), .b(s_56), .O(gate94inter1));
  and2  gate941(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate942(.a(s_56), .O(gate94inter3));
  inv1  gate943(.a(s_57), .O(gate94inter4));
  nand2 gate944(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate945(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate946(.a(G22), .O(gate94inter7));
  inv1  gate947(.a(G344), .O(gate94inter8));
  nand2 gate948(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate949(.a(s_57), .b(gate94inter3), .O(gate94inter10));
  nor2  gate950(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate951(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate952(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate631(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate632(.a(gate97inter0), .b(s_12), .O(gate97inter1));
  and2  gate633(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate634(.a(s_12), .O(gate97inter3));
  inv1  gate635(.a(s_13), .O(gate97inter4));
  nand2 gate636(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate637(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate638(.a(G19), .O(gate97inter7));
  inv1  gate639(.a(G350), .O(gate97inter8));
  nand2 gate640(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate641(.a(s_13), .b(gate97inter3), .O(gate97inter10));
  nor2  gate642(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate643(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate644(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1835(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1836(.a(gate98inter0), .b(s_184), .O(gate98inter1));
  and2  gate1837(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1838(.a(s_184), .O(gate98inter3));
  inv1  gate1839(.a(s_185), .O(gate98inter4));
  nand2 gate1840(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1841(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1842(.a(G23), .O(gate98inter7));
  inv1  gate1843(.a(G350), .O(gate98inter8));
  nand2 gate1844(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1845(.a(s_185), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1846(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1847(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1848(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1037(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1038(.a(gate99inter0), .b(s_70), .O(gate99inter1));
  and2  gate1039(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1040(.a(s_70), .O(gate99inter3));
  inv1  gate1041(.a(s_71), .O(gate99inter4));
  nand2 gate1042(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1043(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1044(.a(G27), .O(gate99inter7));
  inv1  gate1045(.a(G353), .O(gate99inter8));
  nand2 gate1046(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1047(.a(s_71), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1048(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1049(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1050(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1317(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1318(.a(gate101inter0), .b(s_110), .O(gate101inter1));
  and2  gate1319(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1320(.a(s_110), .O(gate101inter3));
  inv1  gate1321(.a(s_111), .O(gate101inter4));
  nand2 gate1322(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1323(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1324(.a(G20), .O(gate101inter7));
  inv1  gate1325(.a(G356), .O(gate101inter8));
  nand2 gate1326(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1327(.a(s_111), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1328(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1329(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1330(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate589(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate590(.a(gate102inter0), .b(s_6), .O(gate102inter1));
  and2  gate591(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate592(.a(s_6), .O(gate102inter3));
  inv1  gate593(.a(s_7), .O(gate102inter4));
  nand2 gate594(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate595(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate596(.a(G24), .O(gate102inter7));
  inv1  gate597(.a(G356), .O(gate102inter8));
  nand2 gate598(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate599(.a(s_7), .b(gate102inter3), .O(gate102inter10));
  nor2  gate600(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate601(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate602(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate645(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate646(.a(gate108inter0), .b(s_14), .O(gate108inter1));
  and2  gate647(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate648(.a(s_14), .O(gate108inter3));
  inv1  gate649(.a(s_15), .O(gate108inter4));
  nand2 gate650(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate651(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate652(.a(G368), .O(gate108inter7));
  inv1  gate653(.a(G369), .O(gate108inter8));
  nand2 gate654(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate655(.a(s_15), .b(gate108inter3), .O(gate108inter10));
  nor2  gate656(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate657(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate658(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate813(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate814(.a(gate114inter0), .b(s_38), .O(gate114inter1));
  and2  gate815(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate816(.a(s_38), .O(gate114inter3));
  inv1  gate817(.a(s_39), .O(gate114inter4));
  nand2 gate818(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate819(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate820(.a(G380), .O(gate114inter7));
  inv1  gate821(.a(G381), .O(gate114inter8));
  nand2 gate822(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate823(.a(s_39), .b(gate114inter3), .O(gate114inter10));
  nor2  gate824(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate825(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate826(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1485(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1486(.a(gate119inter0), .b(s_134), .O(gate119inter1));
  and2  gate1487(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1488(.a(s_134), .O(gate119inter3));
  inv1  gate1489(.a(s_135), .O(gate119inter4));
  nand2 gate1490(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1491(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1492(.a(G390), .O(gate119inter7));
  inv1  gate1493(.a(G391), .O(gate119inter8));
  nand2 gate1494(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1495(.a(s_135), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1496(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1497(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1498(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate827(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate828(.a(gate125inter0), .b(s_40), .O(gate125inter1));
  and2  gate829(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate830(.a(s_40), .O(gate125inter3));
  inv1  gate831(.a(s_41), .O(gate125inter4));
  nand2 gate832(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate833(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate834(.a(G402), .O(gate125inter7));
  inv1  gate835(.a(G403), .O(gate125inter8));
  nand2 gate836(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate837(.a(s_41), .b(gate125inter3), .O(gate125inter10));
  nor2  gate838(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate839(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate840(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1289(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1290(.a(gate128inter0), .b(s_106), .O(gate128inter1));
  and2  gate1291(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1292(.a(s_106), .O(gate128inter3));
  inv1  gate1293(.a(s_107), .O(gate128inter4));
  nand2 gate1294(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1295(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1296(.a(G408), .O(gate128inter7));
  inv1  gate1297(.a(G409), .O(gate128inter8));
  nand2 gate1298(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1299(.a(s_107), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1300(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1301(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1302(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1233(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1234(.a(gate138inter0), .b(s_98), .O(gate138inter1));
  and2  gate1235(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1236(.a(s_98), .O(gate138inter3));
  inv1  gate1237(.a(s_99), .O(gate138inter4));
  nand2 gate1238(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1239(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1240(.a(G432), .O(gate138inter7));
  inv1  gate1241(.a(G435), .O(gate138inter8));
  nand2 gate1242(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1243(.a(s_99), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1244(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1245(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1246(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1079(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1080(.a(gate143inter0), .b(s_76), .O(gate143inter1));
  and2  gate1081(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1082(.a(s_76), .O(gate143inter3));
  inv1  gate1083(.a(s_77), .O(gate143inter4));
  nand2 gate1084(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1085(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1086(.a(G462), .O(gate143inter7));
  inv1  gate1087(.a(G465), .O(gate143inter8));
  nand2 gate1088(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1089(.a(s_77), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1090(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1091(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1092(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1681(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1682(.a(gate146inter0), .b(s_162), .O(gate146inter1));
  and2  gate1683(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1684(.a(s_162), .O(gate146inter3));
  inv1  gate1685(.a(s_163), .O(gate146inter4));
  nand2 gate1686(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1687(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1688(.a(G480), .O(gate146inter7));
  inv1  gate1689(.a(G483), .O(gate146inter8));
  nand2 gate1690(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1691(.a(s_163), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1692(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1693(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1694(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1457(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1458(.a(gate155inter0), .b(s_130), .O(gate155inter1));
  and2  gate1459(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1460(.a(s_130), .O(gate155inter3));
  inv1  gate1461(.a(s_131), .O(gate155inter4));
  nand2 gate1462(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1463(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1464(.a(G432), .O(gate155inter7));
  inv1  gate1465(.a(G525), .O(gate155inter8));
  nand2 gate1466(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1467(.a(s_131), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1468(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1469(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1470(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1345(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1346(.a(gate163inter0), .b(s_114), .O(gate163inter1));
  and2  gate1347(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1348(.a(s_114), .O(gate163inter3));
  inv1  gate1349(.a(s_115), .O(gate163inter4));
  nand2 gate1350(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1351(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1352(.a(G456), .O(gate163inter7));
  inv1  gate1353(.a(G537), .O(gate163inter8));
  nand2 gate1354(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1355(.a(s_115), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1356(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1357(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1358(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate953(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate954(.a(gate170inter0), .b(s_58), .O(gate170inter1));
  and2  gate955(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate956(.a(s_58), .O(gate170inter3));
  inv1  gate957(.a(s_59), .O(gate170inter4));
  nand2 gate958(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate959(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate960(.a(G477), .O(gate170inter7));
  inv1  gate961(.a(G546), .O(gate170inter8));
  nand2 gate962(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate963(.a(s_59), .b(gate170inter3), .O(gate170inter10));
  nor2  gate964(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate965(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate966(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1499(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1500(.a(gate174inter0), .b(s_136), .O(gate174inter1));
  and2  gate1501(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1502(.a(s_136), .O(gate174inter3));
  inv1  gate1503(.a(s_137), .O(gate174inter4));
  nand2 gate1504(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1505(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1506(.a(G489), .O(gate174inter7));
  inv1  gate1507(.a(G552), .O(gate174inter8));
  nand2 gate1508(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1509(.a(s_137), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1510(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1511(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1512(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate715(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate716(.a(gate179inter0), .b(s_24), .O(gate179inter1));
  and2  gate717(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate718(.a(s_24), .O(gate179inter3));
  inv1  gate719(.a(s_25), .O(gate179inter4));
  nand2 gate720(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate721(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate722(.a(G504), .O(gate179inter7));
  inv1  gate723(.a(G561), .O(gate179inter8));
  nand2 gate724(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate725(.a(s_25), .b(gate179inter3), .O(gate179inter10));
  nor2  gate726(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate727(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate728(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate743(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate744(.a(gate181inter0), .b(s_28), .O(gate181inter1));
  and2  gate745(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate746(.a(s_28), .O(gate181inter3));
  inv1  gate747(.a(s_29), .O(gate181inter4));
  nand2 gate748(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate749(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate750(.a(G510), .O(gate181inter7));
  inv1  gate751(.a(G564), .O(gate181inter8));
  nand2 gate752(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate753(.a(s_29), .b(gate181inter3), .O(gate181inter10));
  nor2  gate754(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate755(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate756(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1751(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1752(.a(gate199inter0), .b(s_172), .O(gate199inter1));
  and2  gate1753(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1754(.a(s_172), .O(gate199inter3));
  inv1  gate1755(.a(s_173), .O(gate199inter4));
  nand2 gate1756(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1757(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1758(.a(G598), .O(gate199inter7));
  inv1  gate1759(.a(G599), .O(gate199inter8));
  nand2 gate1760(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1761(.a(s_173), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1762(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1763(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1764(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1331(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1332(.a(gate205inter0), .b(s_112), .O(gate205inter1));
  and2  gate1333(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1334(.a(s_112), .O(gate205inter3));
  inv1  gate1335(.a(s_113), .O(gate205inter4));
  nand2 gate1336(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1337(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1338(.a(G622), .O(gate205inter7));
  inv1  gate1339(.a(G627), .O(gate205inter8));
  nand2 gate1340(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1341(.a(s_113), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1342(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1343(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1344(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate799(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate800(.a(gate207inter0), .b(s_36), .O(gate207inter1));
  and2  gate801(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate802(.a(s_36), .O(gate207inter3));
  inv1  gate803(.a(s_37), .O(gate207inter4));
  nand2 gate804(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate805(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate806(.a(G622), .O(gate207inter7));
  inv1  gate807(.a(G632), .O(gate207inter8));
  nand2 gate808(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate809(.a(s_37), .b(gate207inter3), .O(gate207inter10));
  nor2  gate810(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate811(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate812(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1695(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1696(.a(gate214inter0), .b(s_164), .O(gate214inter1));
  and2  gate1697(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1698(.a(s_164), .O(gate214inter3));
  inv1  gate1699(.a(s_165), .O(gate214inter4));
  nand2 gate1700(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1701(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1702(.a(G612), .O(gate214inter7));
  inv1  gate1703(.a(G672), .O(gate214inter8));
  nand2 gate1704(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1705(.a(s_165), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1706(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1707(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1708(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate603(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate604(.a(gate219inter0), .b(s_8), .O(gate219inter1));
  and2  gate605(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate606(.a(s_8), .O(gate219inter3));
  inv1  gate607(.a(s_9), .O(gate219inter4));
  nand2 gate608(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate609(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate610(.a(G632), .O(gate219inter7));
  inv1  gate611(.a(G681), .O(gate219inter8));
  nand2 gate612(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate613(.a(s_9), .b(gate219inter3), .O(gate219inter10));
  nor2  gate614(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate615(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate616(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1359(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1360(.a(gate222inter0), .b(s_116), .O(gate222inter1));
  and2  gate1361(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1362(.a(s_116), .O(gate222inter3));
  inv1  gate1363(.a(s_117), .O(gate222inter4));
  nand2 gate1364(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1365(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1366(.a(G632), .O(gate222inter7));
  inv1  gate1367(.a(G684), .O(gate222inter8));
  nand2 gate1368(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1369(.a(s_117), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1370(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1371(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1372(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1191(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1192(.a(gate224inter0), .b(s_92), .O(gate224inter1));
  and2  gate1193(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1194(.a(s_92), .O(gate224inter3));
  inv1  gate1195(.a(s_93), .O(gate224inter4));
  nand2 gate1196(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1197(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1198(.a(G637), .O(gate224inter7));
  inv1  gate1199(.a(G687), .O(gate224inter8));
  nand2 gate1200(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1201(.a(s_93), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1202(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1203(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1204(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate575(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate576(.a(gate230inter0), .b(s_4), .O(gate230inter1));
  and2  gate577(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate578(.a(s_4), .O(gate230inter3));
  inv1  gate579(.a(s_5), .O(gate230inter4));
  nand2 gate580(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate581(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate582(.a(G700), .O(gate230inter7));
  inv1  gate583(.a(G701), .O(gate230inter8));
  nand2 gate584(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate585(.a(s_5), .b(gate230inter3), .O(gate230inter10));
  nor2  gate586(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate587(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate588(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate897(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate898(.a(gate231inter0), .b(s_50), .O(gate231inter1));
  and2  gate899(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate900(.a(s_50), .O(gate231inter3));
  inv1  gate901(.a(s_51), .O(gate231inter4));
  nand2 gate902(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate903(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate904(.a(G702), .O(gate231inter7));
  inv1  gate905(.a(G703), .O(gate231inter8));
  nand2 gate906(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate907(.a(s_51), .b(gate231inter3), .O(gate231inter10));
  nor2  gate908(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate909(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate910(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate757(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate758(.a(gate237inter0), .b(s_30), .O(gate237inter1));
  and2  gate759(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate760(.a(s_30), .O(gate237inter3));
  inv1  gate761(.a(s_31), .O(gate237inter4));
  nand2 gate762(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate763(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate764(.a(G254), .O(gate237inter7));
  inv1  gate765(.a(G706), .O(gate237inter8));
  nand2 gate766(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate767(.a(s_31), .b(gate237inter3), .O(gate237inter10));
  nor2  gate768(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate769(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate770(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate701(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate702(.a(gate239inter0), .b(s_22), .O(gate239inter1));
  and2  gate703(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate704(.a(s_22), .O(gate239inter3));
  inv1  gate705(.a(s_23), .O(gate239inter4));
  nand2 gate706(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate707(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate708(.a(G260), .O(gate239inter7));
  inv1  gate709(.a(G712), .O(gate239inter8));
  nand2 gate710(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate711(.a(s_23), .b(gate239inter3), .O(gate239inter10));
  nor2  gate712(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate713(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate714(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate981(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate982(.a(gate240inter0), .b(s_62), .O(gate240inter1));
  and2  gate983(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate984(.a(s_62), .O(gate240inter3));
  inv1  gate985(.a(s_63), .O(gate240inter4));
  nand2 gate986(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate987(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate988(.a(G263), .O(gate240inter7));
  inv1  gate989(.a(G715), .O(gate240inter8));
  nand2 gate990(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate991(.a(s_63), .b(gate240inter3), .O(gate240inter10));
  nor2  gate992(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate993(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate994(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1415(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1416(.a(gate243inter0), .b(s_124), .O(gate243inter1));
  and2  gate1417(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1418(.a(s_124), .O(gate243inter3));
  inv1  gate1419(.a(s_125), .O(gate243inter4));
  nand2 gate1420(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1421(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1422(.a(G245), .O(gate243inter7));
  inv1  gate1423(.a(G733), .O(gate243inter8));
  nand2 gate1424(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1425(.a(s_125), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1426(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1427(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1428(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1443(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1444(.a(gate249inter0), .b(s_128), .O(gate249inter1));
  and2  gate1445(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1446(.a(s_128), .O(gate249inter3));
  inv1  gate1447(.a(s_129), .O(gate249inter4));
  nand2 gate1448(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1449(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1450(.a(G254), .O(gate249inter7));
  inv1  gate1451(.a(G742), .O(gate249inter8));
  nand2 gate1452(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1453(.a(s_129), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1454(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1455(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1456(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1597(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1598(.a(gate255inter0), .b(s_150), .O(gate255inter1));
  and2  gate1599(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1600(.a(s_150), .O(gate255inter3));
  inv1  gate1601(.a(s_151), .O(gate255inter4));
  nand2 gate1602(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1603(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1604(.a(G263), .O(gate255inter7));
  inv1  gate1605(.a(G751), .O(gate255inter8));
  nand2 gate1606(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1607(.a(s_151), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1608(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1609(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1610(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1821(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1822(.a(gate257inter0), .b(s_182), .O(gate257inter1));
  and2  gate1823(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1824(.a(s_182), .O(gate257inter3));
  inv1  gate1825(.a(s_183), .O(gate257inter4));
  nand2 gate1826(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1827(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1828(.a(G754), .O(gate257inter7));
  inv1  gate1829(.a(G755), .O(gate257inter8));
  nand2 gate1830(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1831(.a(s_183), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1832(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1833(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1834(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1107(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1108(.a(gate259inter0), .b(s_80), .O(gate259inter1));
  and2  gate1109(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1110(.a(s_80), .O(gate259inter3));
  inv1  gate1111(.a(s_81), .O(gate259inter4));
  nand2 gate1112(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1113(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1114(.a(G758), .O(gate259inter7));
  inv1  gate1115(.a(G759), .O(gate259inter8));
  nand2 gate1116(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1117(.a(s_81), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1118(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1119(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1120(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1653(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1654(.a(gate266inter0), .b(s_158), .O(gate266inter1));
  and2  gate1655(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1656(.a(s_158), .O(gate266inter3));
  inv1  gate1657(.a(s_159), .O(gate266inter4));
  nand2 gate1658(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1659(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1660(.a(G645), .O(gate266inter7));
  inv1  gate1661(.a(G773), .O(gate266inter8));
  nand2 gate1662(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1663(.a(s_159), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1664(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1665(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1666(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate687(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate688(.a(gate267inter0), .b(s_20), .O(gate267inter1));
  and2  gate689(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate690(.a(s_20), .O(gate267inter3));
  inv1  gate691(.a(s_21), .O(gate267inter4));
  nand2 gate692(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate693(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate694(.a(G648), .O(gate267inter7));
  inv1  gate695(.a(G776), .O(gate267inter8));
  nand2 gate696(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate697(.a(s_21), .b(gate267inter3), .O(gate267inter10));
  nor2  gate698(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate699(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate700(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1639(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1640(.a(gate272inter0), .b(s_156), .O(gate272inter1));
  and2  gate1641(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1642(.a(s_156), .O(gate272inter3));
  inv1  gate1643(.a(s_157), .O(gate272inter4));
  nand2 gate1644(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1645(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1646(.a(G663), .O(gate272inter7));
  inv1  gate1647(.a(G791), .O(gate272inter8));
  nand2 gate1648(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1649(.a(s_157), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1650(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1651(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1652(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1779(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1780(.a(gate279inter0), .b(s_176), .O(gate279inter1));
  and2  gate1781(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1782(.a(s_176), .O(gate279inter3));
  inv1  gate1783(.a(s_177), .O(gate279inter4));
  nand2 gate1784(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1785(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1786(.a(G651), .O(gate279inter7));
  inv1  gate1787(.a(G803), .O(gate279inter8));
  nand2 gate1788(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1789(.a(s_177), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1790(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1791(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1792(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate547(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate548(.a(gate282inter0), .b(s_0), .O(gate282inter1));
  and2  gate549(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate550(.a(s_0), .O(gate282inter3));
  inv1  gate551(.a(s_1), .O(gate282inter4));
  nand2 gate552(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate553(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate554(.a(G782), .O(gate282inter7));
  inv1  gate555(.a(G806), .O(gate282inter8));
  nand2 gate556(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate557(.a(s_1), .b(gate282inter3), .O(gate282inter10));
  nor2  gate558(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate559(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate560(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1121(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1122(.a(gate284inter0), .b(s_82), .O(gate284inter1));
  and2  gate1123(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1124(.a(s_82), .O(gate284inter3));
  inv1  gate1125(.a(s_83), .O(gate284inter4));
  nand2 gate1126(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1127(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1128(.a(G785), .O(gate284inter7));
  inv1  gate1129(.a(G809), .O(gate284inter8));
  nand2 gate1130(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1131(.a(s_83), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1132(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1133(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1134(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1527(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1528(.a(gate285inter0), .b(s_140), .O(gate285inter1));
  and2  gate1529(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1530(.a(s_140), .O(gate285inter3));
  inv1  gate1531(.a(s_141), .O(gate285inter4));
  nand2 gate1532(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1533(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1534(.a(G660), .O(gate285inter7));
  inv1  gate1535(.a(G812), .O(gate285inter8));
  nand2 gate1536(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1537(.a(s_141), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1538(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1539(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1540(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1471(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1472(.a(gate288inter0), .b(s_132), .O(gate288inter1));
  and2  gate1473(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1474(.a(s_132), .O(gate288inter3));
  inv1  gate1475(.a(s_133), .O(gate288inter4));
  nand2 gate1476(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1477(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1478(.a(G791), .O(gate288inter7));
  inv1  gate1479(.a(G815), .O(gate288inter8));
  nand2 gate1480(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1481(.a(s_133), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1482(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1483(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1484(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1541(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1542(.a(gate290inter0), .b(s_142), .O(gate290inter1));
  and2  gate1543(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1544(.a(s_142), .O(gate290inter3));
  inv1  gate1545(.a(s_143), .O(gate290inter4));
  nand2 gate1546(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1547(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1548(.a(G820), .O(gate290inter7));
  inv1  gate1549(.a(G821), .O(gate290inter8));
  nand2 gate1550(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1551(.a(s_143), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1552(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1553(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1554(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1205(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1206(.a(gate291inter0), .b(s_94), .O(gate291inter1));
  and2  gate1207(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1208(.a(s_94), .O(gate291inter3));
  inv1  gate1209(.a(s_95), .O(gate291inter4));
  nand2 gate1210(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1211(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1212(.a(G822), .O(gate291inter7));
  inv1  gate1213(.a(G823), .O(gate291inter8));
  nand2 gate1214(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1215(.a(s_95), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1216(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1217(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1218(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate911(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate912(.a(gate292inter0), .b(s_52), .O(gate292inter1));
  and2  gate913(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate914(.a(s_52), .O(gate292inter3));
  inv1  gate915(.a(s_53), .O(gate292inter4));
  nand2 gate916(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate917(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate918(.a(G824), .O(gate292inter7));
  inv1  gate919(.a(G825), .O(gate292inter8));
  nand2 gate920(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate921(.a(s_53), .b(gate292inter3), .O(gate292inter10));
  nor2  gate922(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate923(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate924(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1135(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1136(.a(gate294inter0), .b(s_84), .O(gate294inter1));
  and2  gate1137(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1138(.a(s_84), .O(gate294inter3));
  inv1  gate1139(.a(s_85), .O(gate294inter4));
  nand2 gate1140(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1141(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1142(.a(G832), .O(gate294inter7));
  inv1  gate1143(.a(G833), .O(gate294inter8));
  nand2 gate1144(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1145(.a(s_85), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1146(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1147(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1148(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1303(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1304(.a(gate388inter0), .b(s_108), .O(gate388inter1));
  and2  gate1305(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1306(.a(s_108), .O(gate388inter3));
  inv1  gate1307(.a(s_109), .O(gate388inter4));
  nand2 gate1308(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1309(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1310(.a(G2), .O(gate388inter7));
  inv1  gate1311(.a(G1039), .O(gate388inter8));
  nand2 gate1312(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1313(.a(s_109), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1314(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1315(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1316(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1163(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1164(.a(gate403inter0), .b(s_88), .O(gate403inter1));
  and2  gate1165(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1166(.a(s_88), .O(gate403inter3));
  inv1  gate1167(.a(s_89), .O(gate403inter4));
  nand2 gate1168(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1169(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1170(.a(G17), .O(gate403inter7));
  inv1  gate1171(.a(G1084), .O(gate403inter8));
  nand2 gate1172(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1173(.a(s_89), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1174(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1175(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1176(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1513(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1514(.a(gate406inter0), .b(s_138), .O(gate406inter1));
  and2  gate1515(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1516(.a(s_138), .O(gate406inter3));
  inv1  gate1517(.a(s_139), .O(gate406inter4));
  nand2 gate1518(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1519(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1520(.a(G20), .O(gate406inter7));
  inv1  gate1521(.a(G1093), .O(gate406inter8));
  nand2 gate1522(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1523(.a(s_139), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1524(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1525(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1526(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1093(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1094(.a(gate410inter0), .b(s_78), .O(gate410inter1));
  and2  gate1095(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1096(.a(s_78), .O(gate410inter3));
  inv1  gate1097(.a(s_79), .O(gate410inter4));
  nand2 gate1098(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1099(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1100(.a(G24), .O(gate410inter7));
  inv1  gate1101(.a(G1105), .O(gate410inter8));
  nand2 gate1102(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1103(.a(s_79), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1104(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1105(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1106(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate995(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate996(.a(gate416inter0), .b(s_64), .O(gate416inter1));
  and2  gate997(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate998(.a(s_64), .O(gate416inter3));
  inv1  gate999(.a(s_65), .O(gate416inter4));
  nand2 gate1000(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1001(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1002(.a(G30), .O(gate416inter7));
  inv1  gate1003(.a(G1123), .O(gate416inter8));
  nand2 gate1004(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1005(.a(s_65), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1006(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1007(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1008(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1765(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1766(.a(gate421inter0), .b(s_174), .O(gate421inter1));
  and2  gate1767(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1768(.a(s_174), .O(gate421inter3));
  inv1  gate1769(.a(s_175), .O(gate421inter4));
  nand2 gate1770(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1771(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1772(.a(G2), .O(gate421inter7));
  inv1  gate1773(.a(G1135), .O(gate421inter8));
  nand2 gate1774(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1775(.a(s_175), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1776(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1777(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1778(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1219(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1220(.a(gate424inter0), .b(s_96), .O(gate424inter1));
  and2  gate1221(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1222(.a(s_96), .O(gate424inter3));
  inv1  gate1223(.a(s_97), .O(gate424inter4));
  nand2 gate1224(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1225(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1226(.a(G1042), .O(gate424inter7));
  inv1  gate1227(.a(G1138), .O(gate424inter8));
  nand2 gate1228(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1229(.a(s_97), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1230(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1231(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1232(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1373(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1374(.a(gate427inter0), .b(s_118), .O(gate427inter1));
  and2  gate1375(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1376(.a(s_118), .O(gate427inter3));
  inv1  gate1377(.a(s_119), .O(gate427inter4));
  nand2 gate1378(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1379(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1380(.a(G5), .O(gate427inter7));
  inv1  gate1381(.a(G1144), .O(gate427inter8));
  nand2 gate1382(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1383(.a(s_119), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1384(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1385(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1386(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1555(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1556(.a(gate433inter0), .b(s_144), .O(gate433inter1));
  and2  gate1557(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1558(.a(s_144), .O(gate433inter3));
  inv1  gate1559(.a(s_145), .O(gate433inter4));
  nand2 gate1560(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1561(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1562(.a(G8), .O(gate433inter7));
  inv1  gate1563(.a(G1153), .O(gate433inter8));
  nand2 gate1564(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1565(.a(s_145), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1566(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1567(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1568(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1401(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1402(.a(gate436inter0), .b(s_122), .O(gate436inter1));
  and2  gate1403(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1404(.a(s_122), .O(gate436inter3));
  inv1  gate1405(.a(s_123), .O(gate436inter4));
  nand2 gate1406(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1407(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1408(.a(G1060), .O(gate436inter7));
  inv1  gate1409(.a(G1156), .O(gate436inter8));
  nand2 gate1410(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1411(.a(s_123), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1412(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1413(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1414(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate883(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate884(.a(gate437inter0), .b(s_48), .O(gate437inter1));
  and2  gate885(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate886(.a(s_48), .O(gate437inter3));
  inv1  gate887(.a(s_49), .O(gate437inter4));
  nand2 gate888(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate889(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate890(.a(G10), .O(gate437inter7));
  inv1  gate891(.a(G1159), .O(gate437inter8));
  nand2 gate892(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate893(.a(s_49), .b(gate437inter3), .O(gate437inter10));
  nor2  gate894(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate895(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate896(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1667(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1668(.a(gate442inter0), .b(s_160), .O(gate442inter1));
  and2  gate1669(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1670(.a(s_160), .O(gate442inter3));
  inv1  gate1671(.a(s_161), .O(gate442inter4));
  nand2 gate1672(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1673(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1674(.a(G1069), .O(gate442inter7));
  inv1  gate1675(.a(G1165), .O(gate442inter8));
  nand2 gate1676(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1677(.a(s_161), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1678(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1679(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1680(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1849(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1850(.a(gate443inter0), .b(s_186), .O(gate443inter1));
  and2  gate1851(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1852(.a(s_186), .O(gate443inter3));
  inv1  gate1853(.a(s_187), .O(gate443inter4));
  nand2 gate1854(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1855(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1856(.a(G13), .O(gate443inter7));
  inv1  gate1857(.a(G1168), .O(gate443inter8));
  nand2 gate1858(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1859(.a(s_187), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1860(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1861(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1862(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate869(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate870(.a(gate444inter0), .b(s_46), .O(gate444inter1));
  and2  gate871(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate872(.a(s_46), .O(gate444inter3));
  inv1  gate873(.a(s_47), .O(gate444inter4));
  nand2 gate874(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate875(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate876(.a(G1072), .O(gate444inter7));
  inv1  gate877(.a(G1168), .O(gate444inter8));
  nand2 gate878(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate879(.a(s_47), .b(gate444inter3), .O(gate444inter10));
  nor2  gate880(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate881(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate882(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1863(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1864(.a(gate451inter0), .b(s_188), .O(gate451inter1));
  and2  gate1865(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1866(.a(s_188), .O(gate451inter3));
  inv1  gate1867(.a(s_189), .O(gate451inter4));
  nand2 gate1868(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1869(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1870(.a(G17), .O(gate451inter7));
  inv1  gate1871(.a(G1180), .O(gate451inter8));
  nand2 gate1872(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1873(.a(s_189), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1874(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1875(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1876(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate841(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate842(.a(gate461inter0), .b(s_42), .O(gate461inter1));
  and2  gate843(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate844(.a(s_42), .O(gate461inter3));
  inv1  gate845(.a(s_43), .O(gate461inter4));
  nand2 gate846(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate847(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate848(.a(G22), .O(gate461inter7));
  inv1  gate849(.a(G1195), .O(gate461inter8));
  nand2 gate850(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate851(.a(s_43), .b(gate461inter3), .O(gate461inter10));
  nor2  gate852(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate853(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate854(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate967(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate968(.a(gate468inter0), .b(s_60), .O(gate468inter1));
  and2  gate969(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate970(.a(s_60), .O(gate468inter3));
  inv1  gate971(.a(s_61), .O(gate468inter4));
  nand2 gate972(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate973(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate974(.a(G1108), .O(gate468inter7));
  inv1  gate975(.a(G1204), .O(gate468inter8));
  nand2 gate976(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate977(.a(s_61), .b(gate468inter3), .O(gate468inter10));
  nor2  gate978(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate979(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate980(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate617(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate618(.a(gate478inter0), .b(s_10), .O(gate478inter1));
  and2  gate619(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate620(.a(s_10), .O(gate478inter3));
  inv1  gate621(.a(s_11), .O(gate478inter4));
  nand2 gate622(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate623(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate624(.a(G1123), .O(gate478inter7));
  inv1  gate625(.a(G1219), .O(gate478inter8));
  nand2 gate626(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate627(.a(s_11), .b(gate478inter3), .O(gate478inter10));
  nor2  gate628(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate629(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate630(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate729(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate730(.a(gate488inter0), .b(s_26), .O(gate488inter1));
  and2  gate731(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate732(.a(s_26), .O(gate488inter3));
  inv1  gate733(.a(s_27), .O(gate488inter4));
  nand2 gate734(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate735(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate736(.a(G1238), .O(gate488inter7));
  inv1  gate737(.a(G1239), .O(gate488inter8));
  nand2 gate738(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate739(.a(s_27), .b(gate488inter3), .O(gate488inter10));
  nor2  gate740(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate741(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate742(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1625(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1626(.a(gate495inter0), .b(s_154), .O(gate495inter1));
  and2  gate1627(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1628(.a(s_154), .O(gate495inter3));
  inv1  gate1629(.a(s_155), .O(gate495inter4));
  nand2 gate1630(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1631(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1632(.a(G1252), .O(gate495inter7));
  inv1  gate1633(.a(G1253), .O(gate495inter8));
  nand2 gate1634(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1635(.a(s_155), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1636(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1637(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1638(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1247(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1248(.a(gate503inter0), .b(s_100), .O(gate503inter1));
  and2  gate1249(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1250(.a(s_100), .O(gate503inter3));
  inv1  gate1251(.a(s_101), .O(gate503inter4));
  nand2 gate1252(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1253(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1254(.a(G1268), .O(gate503inter7));
  inv1  gate1255(.a(G1269), .O(gate503inter8));
  nand2 gate1256(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1257(.a(s_101), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1258(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1259(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1260(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1737(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1738(.a(gate504inter0), .b(s_170), .O(gate504inter1));
  and2  gate1739(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1740(.a(s_170), .O(gate504inter3));
  inv1  gate1741(.a(s_171), .O(gate504inter4));
  nand2 gate1742(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1743(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1744(.a(G1270), .O(gate504inter7));
  inv1  gate1745(.a(G1271), .O(gate504inter8));
  nand2 gate1746(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1747(.a(s_171), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1748(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1749(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1750(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1793(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1794(.a(gate506inter0), .b(s_178), .O(gate506inter1));
  and2  gate1795(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1796(.a(s_178), .O(gate506inter3));
  inv1  gate1797(.a(s_179), .O(gate506inter4));
  nand2 gate1798(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1799(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1800(.a(G1274), .O(gate506inter7));
  inv1  gate1801(.a(G1275), .O(gate506inter8));
  nand2 gate1802(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1803(.a(s_179), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1804(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1805(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1806(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1275(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1276(.a(gate510inter0), .b(s_104), .O(gate510inter1));
  and2  gate1277(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1278(.a(s_104), .O(gate510inter3));
  inv1  gate1279(.a(s_105), .O(gate510inter4));
  nand2 gate1280(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1281(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1282(.a(G1282), .O(gate510inter7));
  inv1  gate1283(.a(G1283), .O(gate510inter8));
  nand2 gate1284(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1285(.a(s_105), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1286(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1287(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1288(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate785(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate786(.a(gate513inter0), .b(s_34), .O(gate513inter1));
  and2  gate787(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate788(.a(s_34), .O(gate513inter3));
  inv1  gate789(.a(s_35), .O(gate513inter4));
  nand2 gate790(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate791(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate792(.a(G1288), .O(gate513inter7));
  inv1  gate793(.a(G1289), .O(gate513inter8));
  nand2 gate794(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate795(.a(s_35), .b(gate513inter3), .O(gate513inter10));
  nor2  gate796(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate797(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate798(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1569(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1570(.a(gate514inter0), .b(s_146), .O(gate514inter1));
  and2  gate1571(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1572(.a(s_146), .O(gate514inter3));
  inv1  gate1573(.a(s_147), .O(gate514inter4));
  nand2 gate1574(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1575(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1576(.a(G1290), .O(gate514inter7));
  inv1  gate1577(.a(G1291), .O(gate514inter8));
  nand2 gate1578(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1579(.a(s_147), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1580(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1581(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1582(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule