module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2493(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2494(.a(gate9inter0), .b(s_278), .O(gate9inter1));
  and2  gate2495(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2496(.a(s_278), .O(gate9inter3));
  inv1  gate2497(.a(s_279), .O(gate9inter4));
  nand2 gate2498(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2499(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2500(.a(G1), .O(gate9inter7));
  inv1  gate2501(.a(G2), .O(gate9inter8));
  nand2 gate2502(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2503(.a(s_279), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2504(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2505(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2506(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2283(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2284(.a(gate13inter0), .b(s_248), .O(gate13inter1));
  and2  gate2285(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2286(.a(s_248), .O(gate13inter3));
  inv1  gate2287(.a(s_249), .O(gate13inter4));
  nand2 gate2288(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2289(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2290(.a(G9), .O(gate13inter7));
  inv1  gate2291(.a(G10), .O(gate13inter8));
  nand2 gate2292(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2293(.a(s_249), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2294(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2295(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2296(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1863(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1864(.a(gate14inter0), .b(s_188), .O(gate14inter1));
  and2  gate1865(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1866(.a(s_188), .O(gate14inter3));
  inv1  gate1867(.a(s_189), .O(gate14inter4));
  nand2 gate1868(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1869(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1870(.a(G11), .O(gate14inter7));
  inv1  gate1871(.a(G12), .O(gate14inter8));
  nand2 gate1872(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1873(.a(s_189), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1874(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1875(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1876(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1485(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1486(.a(gate15inter0), .b(s_134), .O(gate15inter1));
  and2  gate1487(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1488(.a(s_134), .O(gate15inter3));
  inv1  gate1489(.a(s_135), .O(gate15inter4));
  nand2 gate1490(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1491(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1492(.a(G13), .O(gate15inter7));
  inv1  gate1493(.a(G14), .O(gate15inter8));
  nand2 gate1494(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1495(.a(s_135), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1496(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1497(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1498(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2185(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2186(.a(gate17inter0), .b(s_234), .O(gate17inter1));
  and2  gate2187(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2188(.a(s_234), .O(gate17inter3));
  inv1  gate2189(.a(s_235), .O(gate17inter4));
  nand2 gate2190(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2191(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2192(.a(G17), .O(gate17inter7));
  inv1  gate2193(.a(G18), .O(gate17inter8));
  nand2 gate2194(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2195(.a(s_235), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2196(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2197(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2198(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate995(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate996(.a(gate18inter0), .b(s_64), .O(gate18inter1));
  and2  gate997(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate998(.a(s_64), .O(gate18inter3));
  inv1  gate999(.a(s_65), .O(gate18inter4));
  nand2 gate1000(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1001(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1002(.a(G19), .O(gate18inter7));
  inv1  gate1003(.a(G20), .O(gate18inter8));
  nand2 gate1004(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1005(.a(s_65), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1006(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1007(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1008(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1023(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1024(.a(gate20inter0), .b(s_68), .O(gate20inter1));
  and2  gate1025(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1026(.a(s_68), .O(gate20inter3));
  inv1  gate1027(.a(s_69), .O(gate20inter4));
  nand2 gate1028(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1029(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1030(.a(G23), .O(gate20inter7));
  inv1  gate1031(.a(G24), .O(gate20inter8));
  nand2 gate1032(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1033(.a(s_69), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1034(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1035(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1036(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1821(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1822(.a(gate22inter0), .b(s_182), .O(gate22inter1));
  and2  gate1823(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1824(.a(s_182), .O(gate22inter3));
  inv1  gate1825(.a(s_183), .O(gate22inter4));
  nand2 gate1826(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1827(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1828(.a(G27), .O(gate22inter7));
  inv1  gate1829(.a(G28), .O(gate22inter8));
  nand2 gate1830(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1831(.a(s_183), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1832(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1833(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1834(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate743(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate744(.a(gate26inter0), .b(s_28), .O(gate26inter1));
  and2  gate745(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate746(.a(s_28), .O(gate26inter3));
  inv1  gate747(.a(s_29), .O(gate26inter4));
  nand2 gate748(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate749(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate750(.a(G9), .O(gate26inter7));
  inv1  gate751(.a(G13), .O(gate26inter8));
  nand2 gate752(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate753(.a(s_29), .b(gate26inter3), .O(gate26inter10));
  nor2  gate754(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate755(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate756(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1359(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1360(.a(gate35inter0), .b(s_116), .O(gate35inter1));
  and2  gate1361(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1362(.a(s_116), .O(gate35inter3));
  inv1  gate1363(.a(s_117), .O(gate35inter4));
  nand2 gate1364(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1365(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1366(.a(G18), .O(gate35inter7));
  inv1  gate1367(.a(G22), .O(gate35inter8));
  nand2 gate1368(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1369(.a(s_117), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1370(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1371(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1372(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1233(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1234(.a(gate36inter0), .b(s_98), .O(gate36inter1));
  and2  gate1235(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1236(.a(s_98), .O(gate36inter3));
  inv1  gate1237(.a(s_99), .O(gate36inter4));
  nand2 gate1238(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1239(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1240(.a(G26), .O(gate36inter7));
  inv1  gate1241(.a(G30), .O(gate36inter8));
  nand2 gate1242(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1243(.a(s_99), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1244(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1245(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1246(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate575(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate576(.a(gate38inter0), .b(s_4), .O(gate38inter1));
  and2  gate577(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate578(.a(s_4), .O(gate38inter3));
  inv1  gate579(.a(s_5), .O(gate38inter4));
  nand2 gate580(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate581(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate582(.a(G27), .O(gate38inter7));
  inv1  gate583(.a(G31), .O(gate38inter8));
  nand2 gate584(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate585(.a(s_5), .b(gate38inter3), .O(gate38inter10));
  nor2  gate586(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate587(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate588(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1163(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1164(.a(gate39inter0), .b(s_88), .O(gate39inter1));
  and2  gate1165(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1166(.a(s_88), .O(gate39inter3));
  inv1  gate1167(.a(s_89), .O(gate39inter4));
  nand2 gate1168(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1169(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1170(.a(G20), .O(gate39inter7));
  inv1  gate1171(.a(G24), .O(gate39inter8));
  nand2 gate1172(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1173(.a(s_89), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1174(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1175(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1176(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate2367(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2368(.a(gate40inter0), .b(s_260), .O(gate40inter1));
  and2  gate2369(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2370(.a(s_260), .O(gate40inter3));
  inv1  gate2371(.a(s_261), .O(gate40inter4));
  nand2 gate2372(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2373(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2374(.a(G28), .O(gate40inter7));
  inv1  gate2375(.a(G32), .O(gate40inter8));
  nand2 gate2376(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2377(.a(s_261), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2378(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2379(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2380(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate603(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate604(.a(gate41inter0), .b(s_8), .O(gate41inter1));
  and2  gate605(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate606(.a(s_8), .O(gate41inter3));
  inv1  gate607(.a(s_9), .O(gate41inter4));
  nand2 gate608(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate609(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate610(.a(G1), .O(gate41inter7));
  inv1  gate611(.a(G266), .O(gate41inter8));
  nand2 gate612(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate613(.a(s_9), .b(gate41inter3), .O(gate41inter10));
  nor2  gate614(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate615(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate616(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate813(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate814(.a(gate42inter0), .b(s_38), .O(gate42inter1));
  and2  gate815(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate816(.a(s_38), .O(gate42inter3));
  inv1  gate817(.a(s_39), .O(gate42inter4));
  nand2 gate818(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate819(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate820(.a(G2), .O(gate42inter7));
  inv1  gate821(.a(G266), .O(gate42inter8));
  nand2 gate822(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate823(.a(s_39), .b(gate42inter3), .O(gate42inter10));
  nor2  gate824(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate825(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate826(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1583(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1584(.a(gate47inter0), .b(s_148), .O(gate47inter1));
  and2  gate1585(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1586(.a(s_148), .O(gate47inter3));
  inv1  gate1587(.a(s_149), .O(gate47inter4));
  nand2 gate1588(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1589(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1590(.a(G7), .O(gate47inter7));
  inv1  gate1591(.a(G275), .O(gate47inter8));
  nand2 gate1592(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1593(.a(s_149), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1594(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1595(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1596(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1499(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1500(.a(gate51inter0), .b(s_136), .O(gate51inter1));
  and2  gate1501(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1502(.a(s_136), .O(gate51inter3));
  inv1  gate1503(.a(s_137), .O(gate51inter4));
  nand2 gate1504(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1505(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1506(.a(G11), .O(gate51inter7));
  inv1  gate1507(.a(G281), .O(gate51inter8));
  nand2 gate1508(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1509(.a(s_137), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1510(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1511(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1512(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1331(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1332(.a(gate53inter0), .b(s_112), .O(gate53inter1));
  and2  gate1333(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1334(.a(s_112), .O(gate53inter3));
  inv1  gate1335(.a(s_113), .O(gate53inter4));
  nand2 gate1336(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1337(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1338(.a(G13), .O(gate53inter7));
  inv1  gate1339(.a(G284), .O(gate53inter8));
  nand2 gate1340(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1341(.a(s_113), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1342(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1343(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1344(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1681(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1682(.a(gate56inter0), .b(s_162), .O(gate56inter1));
  and2  gate1683(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1684(.a(s_162), .O(gate56inter3));
  inv1  gate1685(.a(s_163), .O(gate56inter4));
  nand2 gate1686(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1687(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1688(.a(G16), .O(gate56inter7));
  inv1  gate1689(.a(G287), .O(gate56inter8));
  nand2 gate1690(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1691(.a(s_163), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1692(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1693(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1694(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1079(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1080(.a(gate61inter0), .b(s_76), .O(gate61inter1));
  and2  gate1081(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1082(.a(s_76), .O(gate61inter3));
  inv1  gate1083(.a(s_77), .O(gate61inter4));
  nand2 gate1084(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1085(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1086(.a(G21), .O(gate61inter7));
  inv1  gate1087(.a(G296), .O(gate61inter8));
  nand2 gate1088(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1089(.a(s_77), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1090(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1091(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1092(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2479(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2480(.a(gate62inter0), .b(s_276), .O(gate62inter1));
  and2  gate2481(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2482(.a(s_276), .O(gate62inter3));
  inv1  gate2483(.a(s_277), .O(gate62inter4));
  nand2 gate2484(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2485(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2486(.a(G22), .O(gate62inter7));
  inv1  gate2487(.a(G296), .O(gate62inter8));
  nand2 gate2488(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2489(.a(s_277), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2490(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2491(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2492(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2311(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2312(.a(gate63inter0), .b(s_252), .O(gate63inter1));
  and2  gate2313(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2314(.a(s_252), .O(gate63inter3));
  inv1  gate2315(.a(s_253), .O(gate63inter4));
  nand2 gate2316(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2317(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2318(.a(G23), .O(gate63inter7));
  inv1  gate2319(.a(G299), .O(gate63inter8));
  nand2 gate2320(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2321(.a(s_253), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2322(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2323(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2324(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2073(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2074(.a(gate67inter0), .b(s_218), .O(gate67inter1));
  and2  gate2075(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2076(.a(s_218), .O(gate67inter3));
  inv1  gate2077(.a(s_219), .O(gate67inter4));
  nand2 gate2078(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2079(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2080(.a(G27), .O(gate67inter7));
  inv1  gate2081(.a(G305), .O(gate67inter8));
  nand2 gate2082(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2083(.a(s_219), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2084(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2085(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2086(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1765(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1766(.a(gate72inter0), .b(s_174), .O(gate72inter1));
  and2  gate1767(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1768(.a(s_174), .O(gate72inter3));
  inv1  gate1769(.a(s_175), .O(gate72inter4));
  nand2 gate1770(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1771(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1772(.a(G32), .O(gate72inter7));
  inv1  gate1773(.a(G311), .O(gate72inter8));
  nand2 gate1774(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1775(.a(s_175), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1776(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1777(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1778(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1261(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1262(.a(gate75inter0), .b(s_102), .O(gate75inter1));
  and2  gate1263(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1264(.a(s_102), .O(gate75inter3));
  inv1  gate1265(.a(s_103), .O(gate75inter4));
  nand2 gate1266(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1267(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1268(.a(G9), .O(gate75inter7));
  inv1  gate1269(.a(G317), .O(gate75inter8));
  nand2 gate1270(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1271(.a(s_103), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1272(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1273(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1274(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate981(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate982(.a(gate76inter0), .b(s_62), .O(gate76inter1));
  and2  gate983(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate984(.a(s_62), .O(gate76inter3));
  inv1  gate985(.a(s_63), .O(gate76inter4));
  nand2 gate986(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate987(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate988(.a(G13), .O(gate76inter7));
  inv1  gate989(.a(G317), .O(gate76inter8));
  nand2 gate990(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate991(.a(s_63), .b(gate76inter3), .O(gate76inter10));
  nor2  gate992(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate993(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate994(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1065(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1066(.a(gate77inter0), .b(s_74), .O(gate77inter1));
  and2  gate1067(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1068(.a(s_74), .O(gate77inter3));
  inv1  gate1069(.a(s_75), .O(gate77inter4));
  nand2 gate1070(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1071(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1072(.a(G2), .O(gate77inter7));
  inv1  gate1073(.a(G320), .O(gate77inter8));
  nand2 gate1074(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1075(.a(s_75), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1076(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1077(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1078(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate2269(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2270(.a(gate78inter0), .b(s_246), .O(gate78inter1));
  and2  gate2271(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2272(.a(s_246), .O(gate78inter3));
  inv1  gate2273(.a(s_247), .O(gate78inter4));
  nand2 gate2274(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2275(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2276(.a(G6), .O(gate78inter7));
  inv1  gate2277(.a(G320), .O(gate78inter8));
  nand2 gate2278(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2279(.a(s_247), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2280(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2281(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2282(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1303(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1304(.a(gate85inter0), .b(s_108), .O(gate85inter1));
  and2  gate1305(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1306(.a(s_108), .O(gate85inter3));
  inv1  gate1307(.a(s_109), .O(gate85inter4));
  nand2 gate1308(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1309(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1310(.a(G4), .O(gate85inter7));
  inv1  gate1311(.a(G332), .O(gate85inter8));
  nand2 gate1312(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1313(.a(s_109), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1314(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1315(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1316(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate645(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate646(.a(gate91inter0), .b(s_14), .O(gate91inter1));
  and2  gate647(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate648(.a(s_14), .O(gate91inter3));
  inv1  gate649(.a(s_15), .O(gate91inter4));
  nand2 gate650(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate651(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate652(.a(G25), .O(gate91inter7));
  inv1  gate653(.a(G341), .O(gate91inter8));
  nand2 gate654(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate655(.a(s_15), .b(gate91inter3), .O(gate91inter10));
  nor2  gate656(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate657(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate658(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1569(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1570(.a(gate92inter0), .b(s_146), .O(gate92inter1));
  and2  gate1571(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1572(.a(s_146), .O(gate92inter3));
  inv1  gate1573(.a(s_147), .O(gate92inter4));
  nand2 gate1574(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1575(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1576(.a(G29), .O(gate92inter7));
  inv1  gate1577(.a(G341), .O(gate92inter8));
  nand2 gate1578(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1579(.a(s_147), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1580(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1581(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1582(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1905(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1906(.a(gate93inter0), .b(s_194), .O(gate93inter1));
  and2  gate1907(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1908(.a(s_194), .O(gate93inter3));
  inv1  gate1909(.a(s_195), .O(gate93inter4));
  nand2 gate1910(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1911(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1912(.a(G18), .O(gate93inter7));
  inv1  gate1913(.a(G344), .O(gate93inter8));
  nand2 gate1914(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1915(.a(s_195), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1916(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1917(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1918(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1037(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1038(.a(gate95inter0), .b(s_70), .O(gate95inter1));
  and2  gate1039(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1040(.a(s_70), .O(gate95inter3));
  inv1  gate1041(.a(s_71), .O(gate95inter4));
  nand2 gate1042(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1043(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1044(.a(G26), .O(gate95inter7));
  inv1  gate1045(.a(G347), .O(gate95inter8));
  nand2 gate1046(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1047(.a(s_71), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1048(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1049(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1050(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1205(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1206(.a(gate99inter0), .b(s_94), .O(gate99inter1));
  and2  gate1207(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1208(.a(s_94), .O(gate99inter3));
  inv1  gate1209(.a(s_95), .O(gate99inter4));
  nand2 gate1210(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1211(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1212(.a(G27), .O(gate99inter7));
  inv1  gate1213(.a(G353), .O(gate99inter8));
  nand2 gate1214(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1215(.a(s_95), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1216(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1217(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1218(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1555(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1556(.a(gate102inter0), .b(s_144), .O(gate102inter1));
  and2  gate1557(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1558(.a(s_144), .O(gate102inter3));
  inv1  gate1559(.a(s_145), .O(gate102inter4));
  nand2 gate1560(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1561(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1562(.a(G24), .O(gate102inter7));
  inv1  gate1563(.a(G356), .O(gate102inter8));
  nand2 gate1564(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1565(.a(s_145), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1566(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1567(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1568(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate799(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate800(.a(gate106inter0), .b(s_36), .O(gate106inter1));
  and2  gate801(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate802(.a(s_36), .O(gate106inter3));
  inv1  gate803(.a(s_37), .O(gate106inter4));
  nand2 gate804(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate805(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate806(.a(G364), .O(gate106inter7));
  inv1  gate807(.a(G365), .O(gate106inter8));
  nand2 gate808(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate809(.a(s_37), .b(gate106inter3), .O(gate106inter10));
  nor2  gate810(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate811(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate812(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate939(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate940(.a(gate109inter0), .b(s_56), .O(gate109inter1));
  and2  gate941(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate942(.a(s_56), .O(gate109inter3));
  inv1  gate943(.a(s_57), .O(gate109inter4));
  nand2 gate944(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate945(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate946(.a(G370), .O(gate109inter7));
  inv1  gate947(.a(G371), .O(gate109inter8));
  nand2 gate948(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate949(.a(s_57), .b(gate109inter3), .O(gate109inter10));
  nor2  gate950(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate951(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate952(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1471(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1472(.a(gate110inter0), .b(s_132), .O(gate110inter1));
  and2  gate1473(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1474(.a(s_132), .O(gate110inter3));
  inv1  gate1475(.a(s_133), .O(gate110inter4));
  nand2 gate1476(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1477(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1478(.a(G372), .O(gate110inter7));
  inv1  gate1479(.a(G373), .O(gate110inter8));
  nand2 gate1480(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1481(.a(s_133), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1482(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1483(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1484(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1947(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1948(.a(gate112inter0), .b(s_200), .O(gate112inter1));
  and2  gate1949(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1950(.a(s_200), .O(gate112inter3));
  inv1  gate1951(.a(s_201), .O(gate112inter4));
  nand2 gate1952(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1953(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1954(.a(G376), .O(gate112inter7));
  inv1  gate1955(.a(G377), .O(gate112inter8));
  nand2 gate1956(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1957(.a(s_201), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1958(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1959(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1960(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1737(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1738(.a(gate115inter0), .b(s_170), .O(gate115inter1));
  and2  gate1739(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1740(.a(s_170), .O(gate115inter3));
  inv1  gate1741(.a(s_171), .O(gate115inter4));
  nand2 gate1742(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1743(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1744(.a(G382), .O(gate115inter7));
  inv1  gate1745(.a(G383), .O(gate115inter8));
  nand2 gate1746(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1747(.a(s_171), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1748(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1749(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1750(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1415(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1416(.a(gate117inter0), .b(s_124), .O(gate117inter1));
  and2  gate1417(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1418(.a(s_124), .O(gate117inter3));
  inv1  gate1419(.a(s_125), .O(gate117inter4));
  nand2 gate1420(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1421(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1422(.a(G386), .O(gate117inter7));
  inv1  gate1423(.a(G387), .O(gate117inter8));
  nand2 gate1424(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1425(.a(s_125), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1426(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1427(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1428(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1107(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1108(.a(gate119inter0), .b(s_80), .O(gate119inter1));
  and2  gate1109(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1110(.a(s_80), .O(gate119inter3));
  inv1  gate1111(.a(s_81), .O(gate119inter4));
  nand2 gate1112(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1113(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1114(.a(G390), .O(gate119inter7));
  inv1  gate1115(.a(G391), .O(gate119inter8));
  nand2 gate1116(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1117(.a(s_81), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1118(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1119(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1120(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1877(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1878(.a(gate120inter0), .b(s_190), .O(gate120inter1));
  and2  gate1879(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1880(.a(s_190), .O(gate120inter3));
  inv1  gate1881(.a(s_191), .O(gate120inter4));
  nand2 gate1882(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1883(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1884(.a(G392), .O(gate120inter7));
  inv1  gate1885(.a(G393), .O(gate120inter8));
  nand2 gate1886(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1887(.a(s_191), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1888(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1889(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1890(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1513(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1514(.a(gate125inter0), .b(s_138), .O(gate125inter1));
  and2  gate1515(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1516(.a(s_138), .O(gate125inter3));
  inv1  gate1517(.a(s_139), .O(gate125inter4));
  nand2 gate1518(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1519(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1520(.a(G402), .O(gate125inter7));
  inv1  gate1521(.a(G403), .O(gate125inter8));
  nand2 gate1522(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1523(.a(s_139), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1524(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1525(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1526(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2339(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2340(.a(gate134inter0), .b(s_256), .O(gate134inter1));
  and2  gate2341(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2342(.a(s_256), .O(gate134inter3));
  inv1  gate2343(.a(s_257), .O(gate134inter4));
  nand2 gate2344(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2345(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2346(.a(G420), .O(gate134inter7));
  inv1  gate2347(.a(G421), .O(gate134inter8));
  nand2 gate2348(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2349(.a(s_257), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2350(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2351(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2352(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1961(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1962(.a(gate136inter0), .b(s_202), .O(gate136inter1));
  and2  gate1963(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1964(.a(s_202), .O(gate136inter3));
  inv1  gate1965(.a(s_203), .O(gate136inter4));
  nand2 gate1966(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1967(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1968(.a(G424), .O(gate136inter7));
  inv1  gate1969(.a(G425), .O(gate136inter8));
  nand2 gate1970(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1971(.a(s_203), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1972(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1973(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1974(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1597(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1598(.a(gate142inter0), .b(s_150), .O(gate142inter1));
  and2  gate1599(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1600(.a(s_150), .O(gate142inter3));
  inv1  gate1601(.a(s_151), .O(gate142inter4));
  nand2 gate1602(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1603(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1604(.a(G456), .O(gate142inter7));
  inv1  gate1605(.a(G459), .O(gate142inter8));
  nand2 gate1606(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1607(.a(s_151), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1608(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1609(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1610(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2059(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2060(.a(gate144inter0), .b(s_216), .O(gate144inter1));
  and2  gate2061(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2062(.a(s_216), .O(gate144inter3));
  inv1  gate2063(.a(s_217), .O(gate144inter4));
  nand2 gate2064(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2065(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2066(.a(G468), .O(gate144inter7));
  inv1  gate2067(.a(G471), .O(gate144inter8));
  nand2 gate2068(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2069(.a(s_217), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2070(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2071(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2072(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2101(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2102(.a(gate146inter0), .b(s_222), .O(gate146inter1));
  and2  gate2103(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2104(.a(s_222), .O(gate146inter3));
  inv1  gate2105(.a(s_223), .O(gate146inter4));
  nand2 gate2106(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2107(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2108(.a(G480), .O(gate146inter7));
  inv1  gate2109(.a(G483), .O(gate146inter8));
  nand2 gate2110(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2111(.a(s_223), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2112(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2113(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2114(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1009(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1010(.a(gate147inter0), .b(s_66), .O(gate147inter1));
  and2  gate1011(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1012(.a(s_66), .O(gate147inter3));
  inv1  gate1013(.a(s_67), .O(gate147inter4));
  nand2 gate1014(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1015(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1016(.a(G486), .O(gate147inter7));
  inv1  gate1017(.a(G489), .O(gate147inter8));
  nand2 gate1018(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1019(.a(s_67), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1020(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1021(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1022(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2003(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2004(.a(gate155inter0), .b(s_208), .O(gate155inter1));
  and2  gate2005(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2006(.a(s_208), .O(gate155inter3));
  inv1  gate2007(.a(s_209), .O(gate155inter4));
  nand2 gate2008(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2009(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2010(.a(G432), .O(gate155inter7));
  inv1  gate2011(.a(G525), .O(gate155inter8));
  nand2 gate2012(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2013(.a(s_209), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2014(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2015(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2016(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate673(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate674(.a(gate162inter0), .b(s_18), .O(gate162inter1));
  and2  gate675(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate676(.a(s_18), .O(gate162inter3));
  inv1  gate677(.a(s_19), .O(gate162inter4));
  nand2 gate678(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate679(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate680(.a(G453), .O(gate162inter7));
  inv1  gate681(.a(G534), .O(gate162inter8));
  nand2 gate682(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate683(.a(s_19), .b(gate162inter3), .O(gate162inter10));
  nor2  gate684(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate685(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate686(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2353(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2354(.a(gate164inter0), .b(s_258), .O(gate164inter1));
  and2  gate2355(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2356(.a(s_258), .O(gate164inter3));
  inv1  gate2357(.a(s_259), .O(gate164inter4));
  nand2 gate2358(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2359(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2360(.a(G459), .O(gate164inter7));
  inv1  gate2361(.a(G537), .O(gate164inter8));
  nand2 gate2362(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2363(.a(s_259), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2364(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2365(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2366(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1149(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1150(.a(gate168inter0), .b(s_86), .O(gate168inter1));
  and2  gate1151(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1152(.a(s_86), .O(gate168inter3));
  inv1  gate1153(.a(s_87), .O(gate168inter4));
  nand2 gate1154(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1155(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1156(.a(G471), .O(gate168inter7));
  inv1  gate1157(.a(G543), .O(gate168inter8));
  nand2 gate1158(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1159(.a(s_87), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1160(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1161(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1162(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2577(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2578(.a(gate172inter0), .b(s_290), .O(gate172inter1));
  and2  gate2579(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2580(.a(s_290), .O(gate172inter3));
  inv1  gate2581(.a(s_291), .O(gate172inter4));
  nand2 gate2582(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2583(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2584(.a(G483), .O(gate172inter7));
  inv1  gate2585(.a(G549), .O(gate172inter8));
  nand2 gate2586(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2587(.a(s_291), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2588(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2589(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2590(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1121(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1122(.a(gate174inter0), .b(s_82), .O(gate174inter1));
  and2  gate1123(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1124(.a(s_82), .O(gate174inter3));
  inv1  gate1125(.a(s_83), .O(gate174inter4));
  nand2 gate1126(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1127(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1128(.a(G489), .O(gate174inter7));
  inv1  gate1129(.a(G552), .O(gate174inter8));
  nand2 gate1130(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1131(.a(s_83), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1132(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1133(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1134(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1933(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1934(.a(gate180inter0), .b(s_198), .O(gate180inter1));
  and2  gate1935(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1936(.a(s_198), .O(gate180inter3));
  inv1  gate1937(.a(s_199), .O(gate180inter4));
  nand2 gate1938(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1939(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1940(.a(G507), .O(gate180inter7));
  inv1  gate1941(.a(G561), .O(gate180inter8));
  nand2 gate1942(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1943(.a(s_199), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1944(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1945(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1946(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate2297(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2298(.a(gate181inter0), .b(s_250), .O(gate181inter1));
  and2  gate2299(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2300(.a(s_250), .O(gate181inter3));
  inv1  gate2301(.a(s_251), .O(gate181inter4));
  nand2 gate2302(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2303(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2304(.a(G510), .O(gate181inter7));
  inv1  gate2305(.a(G564), .O(gate181inter8));
  nand2 gate2306(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2307(.a(s_251), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2308(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2309(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2310(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2157(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2158(.a(gate190inter0), .b(s_230), .O(gate190inter1));
  and2  gate2159(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2160(.a(s_230), .O(gate190inter3));
  inv1  gate2161(.a(s_231), .O(gate190inter4));
  nand2 gate2162(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2163(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2164(.a(G580), .O(gate190inter7));
  inv1  gate2165(.a(G581), .O(gate190inter8));
  nand2 gate2166(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2167(.a(s_231), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2168(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2169(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2170(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2325(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2326(.a(gate191inter0), .b(s_254), .O(gate191inter1));
  and2  gate2327(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2328(.a(s_254), .O(gate191inter3));
  inv1  gate2329(.a(s_255), .O(gate191inter4));
  nand2 gate2330(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2331(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2332(.a(G582), .O(gate191inter7));
  inv1  gate2333(.a(G583), .O(gate191inter8));
  nand2 gate2334(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2335(.a(s_255), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2336(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2337(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2338(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1611(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1612(.a(gate193inter0), .b(s_152), .O(gate193inter1));
  and2  gate1613(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1614(.a(s_152), .O(gate193inter3));
  inv1  gate1615(.a(s_153), .O(gate193inter4));
  nand2 gate1616(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1617(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1618(.a(G586), .O(gate193inter7));
  inv1  gate1619(.a(G587), .O(gate193inter8));
  nand2 gate1620(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1621(.a(s_153), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1622(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1623(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1624(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate771(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate772(.a(gate194inter0), .b(s_32), .O(gate194inter1));
  and2  gate773(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate774(.a(s_32), .O(gate194inter3));
  inv1  gate775(.a(s_33), .O(gate194inter4));
  nand2 gate776(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate777(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate778(.a(G588), .O(gate194inter7));
  inv1  gate779(.a(G589), .O(gate194inter8));
  nand2 gate780(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate781(.a(s_33), .b(gate194inter3), .O(gate194inter10));
  nor2  gate782(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate783(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate784(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1177(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1178(.a(gate197inter0), .b(s_90), .O(gate197inter1));
  and2  gate1179(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1180(.a(s_90), .O(gate197inter3));
  inv1  gate1181(.a(s_91), .O(gate197inter4));
  nand2 gate1182(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1183(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1184(.a(G594), .O(gate197inter7));
  inv1  gate1185(.a(G595), .O(gate197inter8));
  nand2 gate1186(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1187(.a(s_91), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1188(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1189(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1190(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1653(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1654(.a(gate199inter0), .b(s_158), .O(gate199inter1));
  and2  gate1655(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1656(.a(s_158), .O(gate199inter3));
  inv1  gate1657(.a(s_159), .O(gate199inter4));
  nand2 gate1658(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1659(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1660(.a(G598), .O(gate199inter7));
  inv1  gate1661(.a(G599), .O(gate199inter8));
  nand2 gate1662(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1663(.a(s_159), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1664(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1665(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1666(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate883(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate884(.a(gate201inter0), .b(s_48), .O(gate201inter1));
  and2  gate885(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate886(.a(s_48), .O(gate201inter3));
  inv1  gate887(.a(s_49), .O(gate201inter4));
  nand2 gate888(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate889(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate890(.a(G602), .O(gate201inter7));
  inv1  gate891(.a(G607), .O(gate201inter8));
  nand2 gate892(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate893(.a(s_49), .b(gate201inter3), .O(gate201inter10));
  nor2  gate894(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate895(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate896(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1835(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1836(.a(gate202inter0), .b(s_184), .O(gate202inter1));
  and2  gate1837(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1838(.a(s_184), .O(gate202inter3));
  inv1  gate1839(.a(s_185), .O(gate202inter4));
  nand2 gate1840(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1841(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1842(.a(G612), .O(gate202inter7));
  inv1  gate1843(.a(G617), .O(gate202inter8));
  nand2 gate1844(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1845(.a(s_185), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1846(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1847(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1848(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate2465(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2466(.a(gate203inter0), .b(s_274), .O(gate203inter1));
  and2  gate2467(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2468(.a(s_274), .O(gate203inter3));
  inv1  gate2469(.a(s_275), .O(gate203inter4));
  nand2 gate2470(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2471(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2472(.a(G602), .O(gate203inter7));
  inv1  gate2473(.a(G612), .O(gate203inter8));
  nand2 gate2474(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2475(.a(s_275), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2476(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2477(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2478(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1527(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1528(.a(gate206inter0), .b(s_140), .O(gate206inter1));
  and2  gate1529(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1530(.a(s_140), .O(gate206inter3));
  inv1  gate1531(.a(s_141), .O(gate206inter4));
  nand2 gate1532(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1533(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1534(.a(G632), .O(gate206inter7));
  inv1  gate1535(.a(G637), .O(gate206inter8));
  nand2 gate1536(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1537(.a(s_141), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1538(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1539(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1540(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2451(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2452(.a(gate207inter0), .b(s_272), .O(gate207inter1));
  and2  gate2453(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2454(.a(s_272), .O(gate207inter3));
  inv1  gate2455(.a(s_273), .O(gate207inter4));
  nand2 gate2456(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2457(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2458(.a(G622), .O(gate207inter7));
  inv1  gate2459(.a(G632), .O(gate207inter8));
  nand2 gate2460(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2461(.a(s_273), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2462(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2463(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2464(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate967(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate968(.a(gate209inter0), .b(s_60), .O(gate209inter1));
  and2  gate969(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate970(.a(s_60), .O(gate209inter3));
  inv1  gate971(.a(s_61), .O(gate209inter4));
  nand2 gate972(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate973(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate974(.a(G602), .O(gate209inter7));
  inv1  gate975(.a(G666), .O(gate209inter8));
  nand2 gate976(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate977(.a(s_61), .b(gate209inter3), .O(gate209inter10));
  nor2  gate978(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate979(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate980(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1695(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1696(.a(gate210inter0), .b(s_164), .O(gate210inter1));
  and2  gate1697(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1698(.a(s_164), .O(gate210inter3));
  inv1  gate1699(.a(s_165), .O(gate210inter4));
  nand2 gate1700(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1701(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1702(.a(G607), .O(gate210inter7));
  inv1  gate1703(.a(G666), .O(gate210inter8));
  nand2 gate1704(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1705(.a(s_165), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1706(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1707(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1708(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1345(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1346(.a(gate213inter0), .b(s_114), .O(gate213inter1));
  and2  gate1347(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1348(.a(s_114), .O(gate213inter3));
  inv1  gate1349(.a(s_115), .O(gate213inter4));
  nand2 gate1350(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1351(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1352(.a(G602), .O(gate213inter7));
  inv1  gate1353(.a(G672), .O(gate213inter8));
  nand2 gate1354(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1355(.a(s_115), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1356(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1357(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1358(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1219(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1220(.a(gate215inter0), .b(s_96), .O(gate215inter1));
  and2  gate1221(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1222(.a(s_96), .O(gate215inter3));
  inv1  gate1223(.a(s_97), .O(gate215inter4));
  nand2 gate1224(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1225(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1226(.a(G607), .O(gate215inter7));
  inv1  gate1227(.a(G675), .O(gate215inter8));
  nand2 gate1228(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1229(.a(s_97), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1230(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1231(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1232(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1289(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1290(.a(gate216inter0), .b(s_106), .O(gate216inter1));
  and2  gate1291(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1292(.a(s_106), .O(gate216inter3));
  inv1  gate1293(.a(s_107), .O(gate216inter4));
  nand2 gate1294(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1295(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1296(.a(G617), .O(gate216inter7));
  inv1  gate1297(.a(G675), .O(gate216inter8));
  nand2 gate1298(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1299(.a(s_107), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1300(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1301(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1302(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2535(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2536(.a(gate225inter0), .b(s_284), .O(gate225inter1));
  and2  gate2537(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2538(.a(s_284), .O(gate225inter3));
  inv1  gate2539(.a(s_285), .O(gate225inter4));
  nand2 gate2540(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2541(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2542(.a(G690), .O(gate225inter7));
  inv1  gate2543(.a(G691), .O(gate225inter8));
  nand2 gate2544(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2545(.a(s_285), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2546(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2547(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2548(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1247(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1248(.a(gate229inter0), .b(s_100), .O(gate229inter1));
  and2  gate1249(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1250(.a(s_100), .O(gate229inter3));
  inv1  gate1251(.a(s_101), .O(gate229inter4));
  nand2 gate1252(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1253(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1254(.a(G698), .O(gate229inter7));
  inv1  gate1255(.a(G699), .O(gate229inter8));
  nand2 gate1256(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1257(.a(s_101), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1258(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1259(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1260(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1373(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1374(.a(gate230inter0), .b(s_118), .O(gate230inter1));
  and2  gate1375(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1376(.a(s_118), .O(gate230inter3));
  inv1  gate1377(.a(s_119), .O(gate230inter4));
  nand2 gate1378(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1379(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1380(.a(G700), .O(gate230inter7));
  inv1  gate1381(.a(G701), .O(gate230inter8));
  nand2 gate1382(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1383(.a(s_119), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1384(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1385(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1386(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1975(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1976(.a(gate231inter0), .b(s_204), .O(gate231inter1));
  and2  gate1977(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1978(.a(s_204), .O(gate231inter3));
  inv1  gate1979(.a(s_205), .O(gate231inter4));
  nand2 gate1980(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1981(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1982(.a(G702), .O(gate231inter7));
  inv1  gate1983(.a(G703), .O(gate231inter8));
  nand2 gate1984(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1985(.a(s_205), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1986(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1987(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1988(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2549(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2550(.a(gate232inter0), .b(s_286), .O(gate232inter1));
  and2  gate2551(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2552(.a(s_286), .O(gate232inter3));
  inv1  gate2553(.a(s_287), .O(gate232inter4));
  nand2 gate2554(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2555(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2556(.a(G704), .O(gate232inter7));
  inv1  gate2557(.a(G705), .O(gate232inter8));
  nand2 gate2558(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2559(.a(s_287), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2560(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2561(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2562(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1891(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1892(.a(gate234inter0), .b(s_192), .O(gate234inter1));
  and2  gate1893(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1894(.a(s_192), .O(gate234inter3));
  inv1  gate1895(.a(s_193), .O(gate234inter4));
  nand2 gate1896(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1897(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1898(.a(G245), .O(gate234inter7));
  inv1  gate1899(.a(G721), .O(gate234inter8));
  nand2 gate1900(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1901(.a(s_193), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1902(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1903(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1904(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1779(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1780(.a(gate235inter0), .b(s_176), .O(gate235inter1));
  and2  gate1781(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1782(.a(s_176), .O(gate235inter3));
  inv1  gate1783(.a(s_177), .O(gate235inter4));
  nand2 gate1784(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1785(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1786(.a(G248), .O(gate235inter7));
  inv1  gate1787(.a(G724), .O(gate235inter8));
  nand2 gate1788(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1789(.a(s_177), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1790(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1791(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1792(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate953(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate954(.a(gate237inter0), .b(s_58), .O(gate237inter1));
  and2  gate955(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate956(.a(s_58), .O(gate237inter3));
  inv1  gate957(.a(s_59), .O(gate237inter4));
  nand2 gate958(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate959(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate960(.a(G254), .O(gate237inter7));
  inv1  gate961(.a(G706), .O(gate237inter8));
  nand2 gate962(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate963(.a(s_59), .b(gate237inter3), .O(gate237inter10));
  nor2  gate964(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate965(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate966(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1849(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1850(.a(gate238inter0), .b(s_186), .O(gate238inter1));
  and2  gate1851(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1852(.a(s_186), .O(gate238inter3));
  inv1  gate1853(.a(s_187), .O(gate238inter4));
  nand2 gate1854(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1855(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1856(.a(G257), .O(gate238inter7));
  inv1  gate1857(.a(G709), .O(gate238inter8));
  nand2 gate1858(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1859(.a(s_187), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1860(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1861(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1862(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2031(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2032(.a(gate241inter0), .b(s_212), .O(gate241inter1));
  and2  gate2033(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2034(.a(s_212), .O(gate241inter3));
  inv1  gate2035(.a(s_213), .O(gate241inter4));
  nand2 gate2036(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2037(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2038(.a(G242), .O(gate241inter7));
  inv1  gate2039(.a(G730), .O(gate241inter8));
  nand2 gate2040(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2041(.a(s_213), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2042(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2043(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2044(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2423(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2424(.a(gate244inter0), .b(s_268), .O(gate244inter1));
  and2  gate2425(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2426(.a(s_268), .O(gate244inter3));
  inv1  gate2427(.a(s_269), .O(gate244inter4));
  nand2 gate2428(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2429(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2430(.a(G721), .O(gate244inter7));
  inv1  gate2431(.a(G733), .O(gate244inter8));
  nand2 gate2432(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2433(.a(s_269), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2434(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2435(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2436(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate897(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate898(.a(gate247inter0), .b(s_50), .O(gate247inter1));
  and2  gate899(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate900(.a(s_50), .O(gate247inter3));
  inv1  gate901(.a(s_51), .O(gate247inter4));
  nand2 gate902(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate903(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate904(.a(G251), .O(gate247inter7));
  inv1  gate905(.a(G739), .O(gate247inter8));
  nand2 gate906(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate907(.a(s_51), .b(gate247inter3), .O(gate247inter10));
  nor2  gate908(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate909(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate910(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2521(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2522(.a(gate248inter0), .b(s_282), .O(gate248inter1));
  and2  gate2523(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2524(.a(s_282), .O(gate248inter3));
  inv1  gate2525(.a(s_283), .O(gate248inter4));
  nand2 gate2526(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2527(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2528(.a(G727), .O(gate248inter7));
  inv1  gate2529(.a(G739), .O(gate248inter8));
  nand2 gate2530(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2531(.a(s_283), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2532(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2533(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2534(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1429(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1430(.a(gate249inter0), .b(s_126), .O(gate249inter1));
  and2  gate1431(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1432(.a(s_126), .O(gate249inter3));
  inv1  gate1433(.a(s_127), .O(gate249inter4));
  nand2 gate1434(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1435(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1436(.a(G254), .O(gate249inter7));
  inv1  gate1437(.a(G742), .O(gate249inter8));
  nand2 gate1438(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1439(.a(s_127), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1440(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1441(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1442(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2507(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2508(.a(gate253inter0), .b(s_280), .O(gate253inter1));
  and2  gate2509(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2510(.a(s_280), .O(gate253inter3));
  inv1  gate2511(.a(s_281), .O(gate253inter4));
  nand2 gate2512(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2513(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2514(.a(G260), .O(gate253inter7));
  inv1  gate2515(.a(G748), .O(gate253inter8));
  nand2 gate2516(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2517(.a(s_281), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2518(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2519(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2520(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1457(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1458(.a(gate259inter0), .b(s_130), .O(gate259inter1));
  and2  gate1459(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1460(.a(s_130), .O(gate259inter3));
  inv1  gate1461(.a(s_131), .O(gate259inter4));
  nand2 gate1462(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1463(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1464(.a(G758), .O(gate259inter7));
  inv1  gate1465(.a(G759), .O(gate259inter8));
  nand2 gate1466(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1467(.a(s_131), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1468(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1469(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1470(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2199(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2200(.a(gate263inter0), .b(s_236), .O(gate263inter1));
  and2  gate2201(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2202(.a(s_236), .O(gate263inter3));
  inv1  gate2203(.a(s_237), .O(gate263inter4));
  nand2 gate2204(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2205(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2206(.a(G766), .O(gate263inter7));
  inv1  gate2207(.a(G767), .O(gate263inter8));
  nand2 gate2208(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2209(.a(s_237), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2210(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2211(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2212(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2115(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2116(.a(gate267inter0), .b(s_224), .O(gate267inter1));
  and2  gate2117(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2118(.a(s_224), .O(gate267inter3));
  inv1  gate2119(.a(s_225), .O(gate267inter4));
  nand2 gate2120(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2121(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2122(.a(G648), .O(gate267inter7));
  inv1  gate2123(.a(G776), .O(gate267inter8));
  nand2 gate2124(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2125(.a(s_225), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2126(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2127(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2128(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2563(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2564(.a(gate268inter0), .b(s_288), .O(gate268inter1));
  and2  gate2565(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2566(.a(s_288), .O(gate268inter3));
  inv1  gate2567(.a(s_289), .O(gate268inter4));
  nand2 gate2568(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2569(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2570(.a(G651), .O(gate268inter7));
  inv1  gate2571(.a(G779), .O(gate268inter8));
  nand2 gate2572(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2573(.a(s_289), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2574(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2575(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2576(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate827(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate828(.a(gate271inter0), .b(s_40), .O(gate271inter1));
  and2  gate829(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate830(.a(s_40), .O(gate271inter3));
  inv1  gate831(.a(s_41), .O(gate271inter4));
  nand2 gate832(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate833(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate834(.a(G660), .O(gate271inter7));
  inv1  gate835(.a(G788), .O(gate271inter8));
  nand2 gate836(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate837(.a(s_41), .b(gate271inter3), .O(gate271inter10));
  nor2  gate838(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate839(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate840(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate715(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate716(.a(gate276inter0), .b(s_24), .O(gate276inter1));
  and2  gate717(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate718(.a(s_24), .O(gate276inter3));
  inv1  gate719(.a(s_25), .O(gate276inter4));
  nand2 gate720(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate721(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate722(.a(G773), .O(gate276inter7));
  inv1  gate723(.a(G797), .O(gate276inter8));
  nand2 gate724(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate725(.a(s_25), .b(gate276inter3), .O(gate276inter10));
  nor2  gate726(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate727(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate728(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2017(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2018(.a(gate280inter0), .b(s_210), .O(gate280inter1));
  and2  gate2019(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2020(.a(s_210), .O(gate280inter3));
  inv1  gate2021(.a(s_211), .O(gate280inter4));
  nand2 gate2022(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2023(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2024(.a(G779), .O(gate280inter7));
  inv1  gate2025(.a(G803), .O(gate280inter8));
  nand2 gate2026(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2027(.a(s_211), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2028(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2029(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2030(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1625(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1626(.a(gate284inter0), .b(s_154), .O(gate284inter1));
  and2  gate1627(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1628(.a(s_154), .O(gate284inter3));
  inv1  gate1629(.a(s_155), .O(gate284inter4));
  nand2 gate1630(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1631(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1632(.a(G785), .O(gate284inter7));
  inv1  gate1633(.a(G809), .O(gate284inter8));
  nand2 gate1634(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1635(.a(s_155), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1636(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1637(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1638(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1275(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1276(.a(gate288inter0), .b(s_104), .O(gate288inter1));
  and2  gate1277(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1278(.a(s_104), .O(gate288inter3));
  inv1  gate1279(.a(s_105), .O(gate288inter4));
  nand2 gate1280(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1281(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1282(.a(G791), .O(gate288inter7));
  inv1  gate1283(.a(G815), .O(gate288inter8));
  nand2 gate1284(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1285(.a(s_105), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1286(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1287(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1288(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate617(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate618(.a(gate292inter0), .b(s_10), .O(gate292inter1));
  and2  gate619(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate620(.a(s_10), .O(gate292inter3));
  inv1  gate621(.a(s_11), .O(gate292inter4));
  nand2 gate622(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate623(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate624(.a(G824), .O(gate292inter7));
  inv1  gate625(.a(G825), .O(gate292inter8));
  nand2 gate626(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate627(.a(s_11), .b(gate292inter3), .O(gate292inter10));
  nor2  gate628(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate629(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate630(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1093(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1094(.a(gate293inter0), .b(s_78), .O(gate293inter1));
  and2  gate1095(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1096(.a(s_78), .O(gate293inter3));
  inv1  gate1097(.a(s_79), .O(gate293inter4));
  nand2 gate1098(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1099(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1100(.a(G828), .O(gate293inter7));
  inv1  gate1101(.a(G829), .O(gate293inter8));
  nand2 gate1102(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1103(.a(s_79), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1104(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1105(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1106(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate2045(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2046(.a(gate390inter0), .b(s_214), .O(gate390inter1));
  and2  gate2047(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2048(.a(s_214), .O(gate390inter3));
  inv1  gate2049(.a(s_215), .O(gate390inter4));
  nand2 gate2050(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2051(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2052(.a(G4), .O(gate390inter7));
  inv1  gate2053(.a(G1045), .O(gate390inter8));
  nand2 gate2054(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2055(.a(s_215), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2056(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2057(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2058(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1793(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1794(.a(gate391inter0), .b(s_178), .O(gate391inter1));
  and2  gate1795(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1796(.a(s_178), .O(gate391inter3));
  inv1  gate1797(.a(s_179), .O(gate391inter4));
  nand2 gate1798(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1799(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1800(.a(G5), .O(gate391inter7));
  inv1  gate1801(.a(G1048), .O(gate391inter8));
  nand2 gate1802(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1803(.a(s_179), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1804(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1805(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1806(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate785(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate786(.a(gate394inter0), .b(s_34), .O(gate394inter1));
  and2  gate787(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate788(.a(s_34), .O(gate394inter3));
  inv1  gate789(.a(s_35), .O(gate394inter4));
  nand2 gate790(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate791(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate792(.a(G8), .O(gate394inter7));
  inv1  gate793(.a(G1057), .O(gate394inter8));
  nand2 gate794(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate795(.a(s_35), .b(gate394inter3), .O(gate394inter10));
  nor2  gate796(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate797(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate798(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate869(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate870(.a(gate395inter0), .b(s_46), .O(gate395inter1));
  and2  gate871(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate872(.a(s_46), .O(gate395inter3));
  inv1  gate873(.a(s_47), .O(gate395inter4));
  nand2 gate874(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate875(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate876(.a(G9), .O(gate395inter7));
  inv1  gate877(.a(G1060), .O(gate395inter8));
  nand2 gate878(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate879(.a(s_47), .b(gate395inter3), .O(gate395inter10));
  nor2  gate880(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate881(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate882(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1709(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1710(.a(gate400inter0), .b(s_166), .O(gate400inter1));
  and2  gate1711(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1712(.a(s_166), .O(gate400inter3));
  inv1  gate1713(.a(s_167), .O(gate400inter4));
  nand2 gate1714(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1715(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1716(.a(G14), .O(gate400inter7));
  inv1  gate1717(.a(G1075), .O(gate400inter8));
  nand2 gate1718(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1719(.a(s_167), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1720(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1721(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1722(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1723(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1724(.a(gate402inter0), .b(s_168), .O(gate402inter1));
  and2  gate1725(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1726(.a(s_168), .O(gate402inter3));
  inv1  gate1727(.a(s_169), .O(gate402inter4));
  nand2 gate1728(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1729(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1730(.a(G16), .O(gate402inter7));
  inv1  gate1731(.a(G1081), .O(gate402inter8));
  nand2 gate1732(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1733(.a(s_169), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1734(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1735(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1736(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate659(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate660(.a(gate403inter0), .b(s_16), .O(gate403inter1));
  and2  gate661(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate662(.a(s_16), .O(gate403inter3));
  inv1  gate663(.a(s_17), .O(gate403inter4));
  nand2 gate664(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate665(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate666(.a(G17), .O(gate403inter7));
  inv1  gate667(.a(G1084), .O(gate403inter8));
  nand2 gate668(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate669(.a(s_17), .b(gate403inter3), .O(gate403inter10));
  nor2  gate670(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate671(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate672(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1541(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1542(.a(gate409inter0), .b(s_142), .O(gate409inter1));
  and2  gate1543(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1544(.a(s_142), .O(gate409inter3));
  inv1  gate1545(.a(s_143), .O(gate409inter4));
  nand2 gate1546(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1547(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1548(.a(G23), .O(gate409inter7));
  inv1  gate1549(.a(G1102), .O(gate409inter8));
  nand2 gate1550(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1551(.a(s_143), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1552(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1553(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1554(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate589(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate590(.a(gate411inter0), .b(s_6), .O(gate411inter1));
  and2  gate591(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate592(.a(s_6), .O(gate411inter3));
  inv1  gate593(.a(s_7), .O(gate411inter4));
  nand2 gate594(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate595(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate596(.a(G25), .O(gate411inter7));
  inv1  gate597(.a(G1108), .O(gate411inter8));
  nand2 gate598(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate599(.a(s_7), .b(gate411inter3), .O(gate411inter10));
  nor2  gate600(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate601(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate602(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1919(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1920(.a(gate412inter0), .b(s_196), .O(gate412inter1));
  and2  gate1921(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1922(.a(s_196), .O(gate412inter3));
  inv1  gate1923(.a(s_197), .O(gate412inter4));
  nand2 gate1924(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1925(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1926(.a(G26), .O(gate412inter7));
  inv1  gate1927(.a(G1111), .O(gate412inter8));
  nand2 gate1928(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1929(.a(s_197), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1930(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1931(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1932(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate2395(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2396(.a(gate413inter0), .b(s_264), .O(gate413inter1));
  and2  gate2397(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2398(.a(s_264), .O(gate413inter3));
  inv1  gate2399(.a(s_265), .O(gate413inter4));
  nand2 gate2400(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2401(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2402(.a(G27), .O(gate413inter7));
  inv1  gate2403(.a(G1114), .O(gate413inter8));
  nand2 gate2404(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2405(.a(s_265), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2406(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2407(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2408(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2255(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2256(.a(gate417inter0), .b(s_244), .O(gate417inter1));
  and2  gate2257(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2258(.a(s_244), .O(gate417inter3));
  inv1  gate2259(.a(s_245), .O(gate417inter4));
  nand2 gate2260(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2261(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2262(.a(G31), .O(gate417inter7));
  inv1  gate2263(.a(G1126), .O(gate417inter8));
  nand2 gate2264(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2265(.a(s_245), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2266(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2267(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2268(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1387(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1388(.a(gate418inter0), .b(s_120), .O(gate418inter1));
  and2  gate1389(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1390(.a(s_120), .O(gate418inter3));
  inv1  gate1391(.a(s_121), .O(gate418inter4));
  nand2 gate1392(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1393(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1394(.a(G32), .O(gate418inter7));
  inv1  gate1395(.a(G1129), .O(gate418inter8));
  nand2 gate1396(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1397(.a(s_121), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1398(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1399(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1400(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2409(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2410(.a(gate421inter0), .b(s_266), .O(gate421inter1));
  and2  gate2411(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2412(.a(s_266), .O(gate421inter3));
  inv1  gate2413(.a(s_267), .O(gate421inter4));
  nand2 gate2414(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2415(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2416(.a(G2), .O(gate421inter7));
  inv1  gate2417(.a(G1135), .O(gate421inter8));
  nand2 gate2418(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2419(.a(s_267), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2420(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2421(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2422(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1051(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1052(.a(gate422inter0), .b(s_72), .O(gate422inter1));
  and2  gate1053(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1054(.a(s_72), .O(gate422inter3));
  inv1  gate1055(.a(s_73), .O(gate422inter4));
  nand2 gate1056(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1057(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1058(.a(G1039), .O(gate422inter7));
  inv1  gate1059(.a(G1135), .O(gate422inter8));
  nand2 gate1060(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1061(.a(s_73), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1062(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1063(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1064(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2213(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2214(.a(gate424inter0), .b(s_238), .O(gate424inter1));
  and2  gate2215(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2216(.a(s_238), .O(gate424inter3));
  inv1  gate2217(.a(s_239), .O(gate424inter4));
  nand2 gate2218(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2219(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2220(.a(G1042), .O(gate424inter7));
  inv1  gate2221(.a(G1138), .O(gate424inter8));
  nand2 gate2222(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2223(.a(s_239), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2224(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2225(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2226(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1751(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1752(.a(gate425inter0), .b(s_172), .O(gate425inter1));
  and2  gate1753(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1754(.a(s_172), .O(gate425inter3));
  inv1  gate1755(.a(s_173), .O(gate425inter4));
  nand2 gate1756(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1757(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1758(.a(G4), .O(gate425inter7));
  inv1  gate1759(.a(G1141), .O(gate425inter8));
  nand2 gate1760(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1761(.a(s_173), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1762(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1763(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1764(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2129(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2130(.a(gate427inter0), .b(s_226), .O(gate427inter1));
  and2  gate2131(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2132(.a(s_226), .O(gate427inter3));
  inv1  gate2133(.a(s_227), .O(gate427inter4));
  nand2 gate2134(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2135(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2136(.a(G5), .O(gate427inter7));
  inv1  gate2137(.a(G1144), .O(gate427inter8));
  nand2 gate2138(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2139(.a(s_227), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2140(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2141(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2142(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1443(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1444(.a(gate430inter0), .b(s_128), .O(gate430inter1));
  and2  gate1445(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1446(.a(s_128), .O(gate430inter3));
  inv1  gate1447(.a(s_129), .O(gate430inter4));
  nand2 gate1448(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1449(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1450(.a(G1051), .O(gate430inter7));
  inv1  gate1451(.a(G1147), .O(gate430inter8));
  nand2 gate1452(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1453(.a(s_129), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1454(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1455(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1456(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2437(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2438(.a(gate432inter0), .b(s_270), .O(gate432inter1));
  and2  gate2439(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2440(.a(s_270), .O(gate432inter3));
  inv1  gate2441(.a(s_271), .O(gate432inter4));
  nand2 gate2442(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2443(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2444(.a(G1054), .O(gate432inter7));
  inv1  gate2445(.a(G1150), .O(gate432inter8));
  nand2 gate2446(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2447(.a(s_271), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2448(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2449(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2450(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1989(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1990(.a(gate433inter0), .b(s_206), .O(gate433inter1));
  and2  gate1991(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1992(.a(s_206), .O(gate433inter3));
  inv1  gate1993(.a(s_207), .O(gate433inter4));
  nand2 gate1994(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1995(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1996(.a(G8), .O(gate433inter7));
  inv1  gate1997(.a(G1153), .O(gate433inter8));
  nand2 gate1998(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1999(.a(s_207), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2000(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2001(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2002(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate2171(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2172(.a(gate437inter0), .b(s_232), .O(gate437inter1));
  and2  gate2173(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2174(.a(s_232), .O(gate437inter3));
  inv1  gate2175(.a(s_233), .O(gate437inter4));
  nand2 gate2176(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2177(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2178(.a(G10), .O(gate437inter7));
  inv1  gate2179(.a(G1159), .O(gate437inter8));
  nand2 gate2180(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2181(.a(s_233), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2182(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2183(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2184(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1807(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1808(.a(gate442inter0), .b(s_180), .O(gate442inter1));
  and2  gate1809(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1810(.a(s_180), .O(gate442inter3));
  inv1  gate1811(.a(s_181), .O(gate442inter4));
  nand2 gate1812(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1813(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1814(.a(G1069), .O(gate442inter7));
  inv1  gate1815(.a(G1165), .O(gate442inter8));
  nand2 gate1816(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1817(.a(s_181), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1818(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1819(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1820(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1191(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1192(.a(gate443inter0), .b(s_92), .O(gate443inter1));
  and2  gate1193(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1194(.a(s_92), .O(gate443inter3));
  inv1  gate1195(.a(s_93), .O(gate443inter4));
  nand2 gate1196(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1197(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1198(.a(G13), .O(gate443inter7));
  inv1  gate1199(.a(G1168), .O(gate443inter8));
  nand2 gate1200(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1201(.a(s_93), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1202(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1203(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1204(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1317(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1318(.a(gate445inter0), .b(s_110), .O(gate445inter1));
  and2  gate1319(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1320(.a(s_110), .O(gate445inter3));
  inv1  gate1321(.a(s_111), .O(gate445inter4));
  nand2 gate1322(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1323(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1324(.a(G14), .O(gate445inter7));
  inv1  gate1325(.a(G1171), .O(gate445inter8));
  nand2 gate1326(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1327(.a(s_111), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1328(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1329(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1330(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1401(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1402(.a(gate450inter0), .b(s_122), .O(gate450inter1));
  and2  gate1403(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1404(.a(s_122), .O(gate450inter3));
  inv1  gate1405(.a(s_123), .O(gate450inter4));
  nand2 gate1406(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1407(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1408(.a(G1081), .O(gate450inter7));
  inv1  gate1409(.a(G1177), .O(gate450inter8));
  nand2 gate1410(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1411(.a(s_123), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1412(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1413(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1414(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate729(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate730(.a(gate451inter0), .b(s_26), .O(gate451inter1));
  and2  gate731(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate732(.a(s_26), .O(gate451inter3));
  inv1  gate733(.a(s_27), .O(gate451inter4));
  nand2 gate734(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate735(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate736(.a(G17), .O(gate451inter7));
  inv1  gate737(.a(G1180), .O(gate451inter8));
  nand2 gate738(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate739(.a(s_27), .b(gate451inter3), .O(gate451inter10));
  nor2  gate740(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate741(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate742(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1135(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1136(.a(gate463inter0), .b(s_84), .O(gate463inter1));
  and2  gate1137(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1138(.a(s_84), .O(gate463inter3));
  inv1  gate1139(.a(s_85), .O(gate463inter4));
  nand2 gate1140(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1141(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1142(.a(G23), .O(gate463inter7));
  inv1  gate1143(.a(G1198), .O(gate463inter8));
  nand2 gate1144(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1145(.a(s_85), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1146(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1147(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1148(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate701(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate702(.a(gate464inter0), .b(s_22), .O(gate464inter1));
  and2  gate703(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate704(.a(s_22), .O(gate464inter3));
  inv1  gate705(.a(s_23), .O(gate464inter4));
  nand2 gate706(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate707(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate708(.a(G1102), .O(gate464inter7));
  inv1  gate709(.a(G1198), .O(gate464inter8));
  nand2 gate710(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate711(.a(s_23), .b(gate464inter3), .O(gate464inter10));
  nor2  gate712(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate713(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate714(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2381(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2382(.a(gate465inter0), .b(s_262), .O(gate465inter1));
  and2  gate2383(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2384(.a(s_262), .O(gate465inter3));
  inv1  gate2385(.a(s_263), .O(gate465inter4));
  nand2 gate2386(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2387(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2388(.a(G24), .O(gate465inter7));
  inv1  gate2389(.a(G1201), .O(gate465inter8));
  nand2 gate2390(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2391(.a(s_263), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2392(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2393(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2394(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate547(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate548(.a(gate466inter0), .b(s_0), .O(gate466inter1));
  and2  gate549(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate550(.a(s_0), .O(gate466inter3));
  inv1  gate551(.a(s_1), .O(gate466inter4));
  nand2 gate552(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate553(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate554(.a(G1105), .O(gate466inter7));
  inv1  gate555(.a(G1201), .O(gate466inter8));
  nand2 gate556(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate557(.a(s_1), .b(gate466inter3), .O(gate466inter10));
  nor2  gate558(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate559(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate560(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate757(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate758(.a(gate467inter0), .b(s_30), .O(gate467inter1));
  and2  gate759(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate760(.a(s_30), .O(gate467inter3));
  inv1  gate761(.a(s_31), .O(gate467inter4));
  nand2 gate762(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate763(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate764(.a(G25), .O(gate467inter7));
  inv1  gate765(.a(G1204), .O(gate467inter8));
  nand2 gate766(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate767(.a(s_31), .b(gate467inter3), .O(gate467inter10));
  nor2  gate768(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate769(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate770(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate561(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate562(.a(gate472inter0), .b(s_2), .O(gate472inter1));
  and2  gate563(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate564(.a(s_2), .O(gate472inter3));
  inv1  gate565(.a(s_3), .O(gate472inter4));
  nand2 gate566(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate567(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate568(.a(G1114), .O(gate472inter7));
  inv1  gate569(.a(G1210), .O(gate472inter8));
  nand2 gate570(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate571(.a(s_3), .b(gate472inter3), .O(gate472inter10));
  nor2  gate572(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate573(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate574(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate631(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate632(.a(gate474inter0), .b(s_12), .O(gate474inter1));
  and2  gate633(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate634(.a(s_12), .O(gate474inter3));
  inv1  gate635(.a(s_13), .O(gate474inter4));
  nand2 gate636(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate637(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate638(.a(G1117), .O(gate474inter7));
  inv1  gate639(.a(G1213), .O(gate474inter8));
  nand2 gate640(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate641(.a(s_13), .b(gate474inter3), .O(gate474inter10));
  nor2  gate642(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate643(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate644(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1639(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1640(.a(gate475inter0), .b(s_156), .O(gate475inter1));
  and2  gate1641(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1642(.a(s_156), .O(gate475inter3));
  inv1  gate1643(.a(s_157), .O(gate475inter4));
  nand2 gate1644(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1645(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1646(.a(G29), .O(gate475inter7));
  inv1  gate1647(.a(G1216), .O(gate475inter8));
  nand2 gate1648(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1649(.a(s_157), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1650(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1651(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1652(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate925(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate926(.a(gate485inter0), .b(s_54), .O(gate485inter1));
  and2  gate927(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate928(.a(s_54), .O(gate485inter3));
  inv1  gate929(.a(s_55), .O(gate485inter4));
  nand2 gate930(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate931(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate932(.a(G1232), .O(gate485inter7));
  inv1  gate933(.a(G1233), .O(gate485inter8));
  nand2 gate934(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate935(.a(s_55), .b(gate485inter3), .O(gate485inter10));
  nor2  gate936(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate937(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate938(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate855(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate856(.a(gate486inter0), .b(s_44), .O(gate486inter1));
  and2  gate857(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate858(.a(s_44), .O(gate486inter3));
  inv1  gate859(.a(s_45), .O(gate486inter4));
  nand2 gate860(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate861(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate862(.a(G1234), .O(gate486inter7));
  inv1  gate863(.a(G1235), .O(gate486inter8));
  nand2 gate864(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate865(.a(s_45), .b(gate486inter3), .O(gate486inter10));
  nor2  gate866(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate867(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate868(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2143(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2144(.a(gate489inter0), .b(s_228), .O(gate489inter1));
  and2  gate2145(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2146(.a(s_228), .O(gate489inter3));
  inv1  gate2147(.a(s_229), .O(gate489inter4));
  nand2 gate2148(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2149(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2150(.a(G1240), .O(gate489inter7));
  inv1  gate2151(.a(G1241), .O(gate489inter8));
  nand2 gate2152(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2153(.a(s_229), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2154(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2155(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2156(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate687(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate688(.a(gate497inter0), .b(s_20), .O(gate497inter1));
  and2  gate689(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate690(.a(s_20), .O(gate497inter3));
  inv1  gate691(.a(s_21), .O(gate497inter4));
  nand2 gate692(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate693(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate694(.a(G1256), .O(gate497inter7));
  inv1  gate695(.a(G1257), .O(gate497inter8));
  nand2 gate696(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate697(.a(s_21), .b(gate497inter3), .O(gate497inter10));
  nor2  gate698(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate699(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate700(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate2241(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2242(.a(gate498inter0), .b(s_242), .O(gate498inter1));
  and2  gate2243(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2244(.a(s_242), .O(gate498inter3));
  inv1  gate2245(.a(s_243), .O(gate498inter4));
  nand2 gate2246(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2247(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2248(.a(G1258), .O(gate498inter7));
  inv1  gate2249(.a(G1259), .O(gate498inter8));
  nand2 gate2250(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2251(.a(s_243), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2252(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2253(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2254(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate841(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate842(.a(gate499inter0), .b(s_42), .O(gate499inter1));
  and2  gate843(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate844(.a(s_42), .O(gate499inter3));
  inv1  gate845(.a(s_43), .O(gate499inter4));
  nand2 gate846(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate847(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate848(.a(G1260), .O(gate499inter7));
  inv1  gate849(.a(G1261), .O(gate499inter8));
  nand2 gate850(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate851(.a(s_43), .b(gate499inter3), .O(gate499inter10));
  nor2  gate852(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate853(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate854(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2087(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2088(.a(gate506inter0), .b(s_220), .O(gate506inter1));
  and2  gate2089(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2090(.a(s_220), .O(gate506inter3));
  inv1  gate2091(.a(s_221), .O(gate506inter4));
  nand2 gate2092(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2093(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2094(.a(G1274), .O(gate506inter7));
  inv1  gate2095(.a(G1275), .O(gate506inter8));
  nand2 gate2096(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2097(.a(s_221), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2098(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2099(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2100(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1667(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1668(.a(gate508inter0), .b(s_160), .O(gate508inter1));
  and2  gate1669(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1670(.a(s_160), .O(gate508inter3));
  inv1  gate1671(.a(s_161), .O(gate508inter4));
  nand2 gate1672(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1673(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1674(.a(G1278), .O(gate508inter7));
  inv1  gate1675(.a(G1279), .O(gate508inter8));
  nand2 gate1676(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1677(.a(s_161), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1678(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1679(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1680(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate911(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate912(.a(gate513inter0), .b(s_52), .O(gate513inter1));
  and2  gate913(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate914(.a(s_52), .O(gate513inter3));
  inv1  gate915(.a(s_53), .O(gate513inter4));
  nand2 gate916(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate917(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate918(.a(G1288), .O(gate513inter7));
  inv1  gate919(.a(G1289), .O(gate513inter8));
  nand2 gate920(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate921(.a(s_53), .b(gate513inter3), .O(gate513inter10));
  nor2  gate922(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate923(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate924(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate2227(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2228(.a(gate514inter0), .b(s_240), .O(gate514inter1));
  and2  gate2229(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2230(.a(s_240), .O(gate514inter3));
  inv1  gate2231(.a(s_241), .O(gate514inter4));
  nand2 gate2232(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2233(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2234(.a(G1290), .O(gate514inter7));
  inv1  gate2235(.a(G1291), .O(gate514inter8));
  nand2 gate2236(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2237(.a(s_241), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2238(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2239(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2240(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule