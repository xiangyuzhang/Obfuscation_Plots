module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1765(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1766(.a(gate9inter0), .b(s_174), .O(gate9inter1));
  and2  gate1767(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1768(.a(s_174), .O(gate9inter3));
  inv1  gate1769(.a(s_175), .O(gate9inter4));
  nand2 gate1770(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1771(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1772(.a(G1), .O(gate9inter7));
  inv1  gate1773(.a(G2), .O(gate9inter8));
  nand2 gate1774(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1775(.a(s_175), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1776(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1777(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1778(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate869(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate870(.a(gate15inter0), .b(s_46), .O(gate15inter1));
  and2  gate871(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate872(.a(s_46), .O(gate15inter3));
  inv1  gate873(.a(s_47), .O(gate15inter4));
  nand2 gate874(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate875(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate876(.a(G13), .O(gate15inter7));
  inv1  gate877(.a(G14), .O(gate15inter8));
  nand2 gate878(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate879(.a(s_47), .b(gate15inter3), .O(gate15inter10));
  nor2  gate880(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate881(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate882(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1569(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1570(.a(gate16inter0), .b(s_146), .O(gate16inter1));
  and2  gate1571(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1572(.a(s_146), .O(gate16inter3));
  inv1  gate1573(.a(s_147), .O(gate16inter4));
  nand2 gate1574(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1575(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1576(.a(G15), .O(gate16inter7));
  inv1  gate1577(.a(G16), .O(gate16inter8));
  nand2 gate1578(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1579(.a(s_147), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1580(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1581(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1582(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate631(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate632(.a(gate18inter0), .b(s_12), .O(gate18inter1));
  and2  gate633(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate634(.a(s_12), .O(gate18inter3));
  inv1  gate635(.a(s_13), .O(gate18inter4));
  nand2 gate636(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate637(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate638(.a(G19), .O(gate18inter7));
  inv1  gate639(.a(G20), .O(gate18inter8));
  nand2 gate640(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate641(.a(s_13), .b(gate18inter3), .O(gate18inter10));
  nor2  gate642(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate643(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate644(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1597(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1598(.a(gate20inter0), .b(s_150), .O(gate20inter1));
  and2  gate1599(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1600(.a(s_150), .O(gate20inter3));
  inv1  gate1601(.a(s_151), .O(gate20inter4));
  nand2 gate1602(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1603(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1604(.a(G23), .O(gate20inter7));
  inv1  gate1605(.a(G24), .O(gate20inter8));
  nand2 gate1606(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1607(.a(s_151), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1608(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1609(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1610(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1093(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1094(.a(gate26inter0), .b(s_78), .O(gate26inter1));
  and2  gate1095(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1096(.a(s_78), .O(gate26inter3));
  inv1  gate1097(.a(s_79), .O(gate26inter4));
  nand2 gate1098(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1099(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1100(.a(G9), .O(gate26inter7));
  inv1  gate1101(.a(G13), .O(gate26inter8));
  nand2 gate1102(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1103(.a(s_79), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1104(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1105(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1106(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate813(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate814(.a(gate28inter0), .b(s_38), .O(gate28inter1));
  and2  gate815(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate816(.a(s_38), .O(gate28inter3));
  inv1  gate817(.a(s_39), .O(gate28inter4));
  nand2 gate818(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate819(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate820(.a(G10), .O(gate28inter7));
  inv1  gate821(.a(G14), .O(gate28inter8));
  nand2 gate822(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate823(.a(s_39), .b(gate28inter3), .O(gate28inter10));
  nor2  gate824(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate825(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate826(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate729(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate730(.a(gate29inter0), .b(s_26), .O(gate29inter1));
  and2  gate731(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate732(.a(s_26), .O(gate29inter3));
  inv1  gate733(.a(s_27), .O(gate29inter4));
  nand2 gate734(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate735(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate736(.a(G3), .O(gate29inter7));
  inv1  gate737(.a(G7), .O(gate29inter8));
  nand2 gate738(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate739(.a(s_27), .b(gate29inter3), .O(gate29inter10));
  nor2  gate740(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate741(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate742(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1527(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1528(.a(gate33inter0), .b(s_140), .O(gate33inter1));
  and2  gate1529(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1530(.a(s_140), .O(gate33inter3));
  inv1  gate1531(.a(s_141), .O(gate33inter4));
  nand2 gate1532(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1533(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1534(.a(G17), .O(gate33inter7));
  inv1  gate1535(.a(G21), .O(gate33inter8));
  nand2 gate1536(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1537(.a(s_141), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1538(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1539(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1540(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1471(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1472(.a(gate38inter0), .b(s_132), .O(gate38inter1));
  and2  gate1473(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1474(.a(s_132), .O(gate38inter3));
  inv1  gate1475(.a(s_133), .O(gate38inter4));
  nand2 gate1476(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1477(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1478(.a(G27), .O(gate38inter7));
  inv1  gate1479(.a(G31), .O(gate38inter8));
  nand2 gate1480(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1481(.a(s_133), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1482(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1483(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1484(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate547(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate548(.a(gate45inter0), .b(s_0), .O(gate45inter1));
  and2  gate549(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate550(.a(s_0), .O(gate45inter3));
  inv1  gate551(.a(s_1), .O(gate45inter4));
  nand2 gate552(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate553(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate554(.a(G5), .O(gate45inter7));
  inv1  gate555(.a(G272), .O(gate45inter8));
  nand2 gate556(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate557(.a(s_1), .b(gate45inter3), .O(gate45inter10));
  nor2  gate558(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate559(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate560(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1513(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1514(.a(gate48inter0), .b(s_138), .O(gate48inter1));
  and2  gate1515(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1516(.a(s_138), .O(gate48inter3));
  inv1  gate1517(.a(s_139), .O(gate48inter4));
  nand2 gate1518(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1519(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1520(.a(G8), .O(gate48inter7));
  inv1  gate1521(.a(G275), .O(gate48inter8));
  nand2 gate1522(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1523(.a(s_139), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1524(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1525(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1526(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate575(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate576(.a(gate52inter0), .b(s_4), .O(gate52inter1));
  and2  gate577(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate578(.a(s_4), .O(gate52inter3));
  inv1  gate579(.a(s_5), .O(gate52inter4));
  nand2 gate580(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate581(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate582(.a(G12), .O(gate52inter7));
  inv1  gate583(.a(G281), .O(gate52inter8));
  nand2 gate584(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate585(.a(s_5), .b(gate52inter3), .O(gate52inter10));
  nor2  gate586(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate587(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate588(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate687(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate688(.a(gate55inter0), .b(s_20), .O(gate55inter1));
  and2  gate689(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate690(.a(s_20), .O(gate55inter3));
  inv1  gate691(.a(s_21), .O(gate55inter4));
  nand2 gate692(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate693(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate694(.a(G15), .O(gate55inter7));
  inv1  gate695(.a(G287), .O(gate55inter8));
  nand2 gate696(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate697(.a(s_21), .b(gate55inter3), .O(gate55inter10));
  nor2  gate698(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate699(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate700(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1051(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1052(.a(gate56inter0), .b(s_72), .O(gate56inter1));
  and2  gate1053(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1054(.a(s_72), .O(gate56inter3));
  inv1  gate1055(.a(s_73), .O(gate56inter4));
  nand2 gate1056(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1057(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1058(.a(G16), .O(gate56inter7));
  inv1  gate1059(.a(G287), .O(gate56inter8));
  nand2 gate1060(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1061(.a(s_73), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1062(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1063(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1064(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1023(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1024(.a(gate59inter0), .b(s_68), .O(gate59inter1));
  and2  gate1025(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1026(.a(s_68), .O(gate59inter3));
  inv1  gate1027(.a(s_69), .O(gate59inter4));
  nand2 gate1028(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1029(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1030(.a(G19), .O(gate59inter7));
  inv1  gate1031(.a(G293), .O(gate59inter8));
  nand2 gate1032(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1033(.a(s_69), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1034(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1035(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1036(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1205(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1206(.a(gate63inter0), .b(s_94), .O(gate63inter1));
  and2  gate1207(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1208(.a(s_94), .O(gate63inter3));
  inv1  gate1209(.a(s_95), .O(gate63inter4));
  nand2 gate1210(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1211(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1212(.a(G23), .O(gate63inter7));
  inv1  gate1213(.a(G299), .O(gate63inter8));
  nand2 gate1214(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1215(.a(s_95), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1216(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1217(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1218(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1331(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1332(.a(gate65inter0), .b(s_112), .O(gate65inter1));
  and2  gate1333(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1334(.a(s_112), .O(gate65inter3));
  inv1  gate1335(.a(s_113), .O(gate65inter4));
  nand2 gate1336(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1337(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1338(.a(G25), .O(gate65inter7));
  inv1  gate1339(.a(G302), .O(gate65inter8));
  nand2 gate1340(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1341(.a(s_113), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1342(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1343(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1344(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate785(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate786(.a(gate67inter0), .b(s_34), .O(gate67inter1));
  and2  gate787(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate788(.a(s_34), .O(gate67inter3));
  inv1  gate789(.a(s_35), .O(gate67inter4));
  nand2 gate790(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate791(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate792(.a(G27), .O(gate67inter7));
  inv1  gate793(.a(G305), .O(gate67inter8));
  nand2 gate794(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate795(.a(s_35), .b(gate67inter3), .O(gate67inter10));
  nor2  gate796(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate797(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate798(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1373(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1374(.a(gate72inter0), .b(s_118), .O(gate72inter1));
  and2  gate1375(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1376(.a(s_118), .O(gate72inter3));
  inv1  gate1377(.a(s_119), .O(gate72inter4));
  nand2 gate1378(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1379(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1380(.a(G32), .O(gate72inter7));
  inv1  gate1381(.a(G311), .O(gate72inter8));
  nand2 gate1382(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1383(.a(s_119), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1384(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1385(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1386(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1779(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1780(.a(gate78inter0), .b(s_176), .O(gate78inter1));
  and2  gate1781(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1782(.a(s_176), .O(gate78inter3));
  inv1  gate1783(.a(s_177), .O(gate78inter4));
  nand2 gate1784(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1785(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1786(.a(G6), .O(gate78inter7));
  inv1  gate1787(.a(G320), .O(gate78inter8));
  nand2 gate1788(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1789(.a(s_177), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1790(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1791(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1792(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate827(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate828(.a(gate80inter0), .b(s_40), .O(gate80inter1));
  and2  gate829(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate830(.a(s_40), .O(gate80inter3));
  inv1  gate831(.a(s_41), .O(gate80inter4));
  nand2 gate832(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate833(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate834(.a(G14), .O(gate80inter7));
  inv1  gate835(.a(G323), .O(gate80inter8));
  nand2 gate836(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate837(.a(s_41), .b(gate80inter3), .O(gate80inter10));
  nor2  gate838(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate839(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate840(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1611(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1612(.a(gate85inter0), .b(s_152), .O(gate85inter1));
  and2  gate1613(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1614(.a(s_152), .O(gate85inter3));
  inv1  gate1615(.a(s_153), .O(gate85inter4));
  nand2 gate1616(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1617(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1618(.a(G4), .O(gate85inter7));
  inv1  gate1619(.a(G332), .O(gate85inter8));
  nand2 gate1620(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1621(.a(s_153), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1622(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1623(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1624(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1709(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1710(.a(gate91inter0), .b(s_166), .O(gate91inter1));
  and2  gate1711(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1712(.a(s_166), .O(gate91inter3));
  inv1  gate1713(.a(s_167), .O(gate91inter4));
  nand2 gate1714(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1715(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1716(.a(G25), .O(gate91inter7));
  inv1  gate1717(.a(G341), .O(gate91inter8));
  nand2 gate1718(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1719(.a(s_167), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1720(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1721(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1722(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate589(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate590(.a(gate93inter0), .b(s_6), .O(gate93inter1));
  and2  gate591(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate592(.a(s_6), .O(gate93inter3));
  inv1  gate593(.a(s_7), .O(gate93inter4));
  nand2 gate594(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate595(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate596(.a(G18), .O(gate93inter7));
  inv1  gate597(.a(G344), .O(gate93inter8));
  nand2 gate598(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate599(.a(s_7), .b(gate93inter3), .O(gate93inter10));
  nor2  gate600(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate601(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate602(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1261(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1262(.a(gate97inter0), .b(s_102), .O(gate97inter1));
  and2  gate1263(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1264(.a(s_102), .O(gate97inter3));
  inv1  gate1265(.a(s_103), .O(gate97inter4));
  nand2 gate1266(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1267(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1268(.a(G19), .O(gate97inter7));
  inv1  gate1269(.a(G350), .O(gate97inter8));
  nand2 gate1270(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1271(.a(s_103), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1272(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1273(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1274(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1681(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1682(.a(gate98inter0), .b(s_162), .O(gate98inter1));
  and2  gate1683(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1684(.a(s_162), .O(gate98inter3));
  inv1  gate1685(.a(s_163), .O(gate98inter4));
  nand2 gate1686(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1687(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1688(.a(G23), .O(gate98inter7));
  inv1  gate1689(.a(G350), .O(gate98inter8));
  nand2 gate1690(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1691(.a(s_163), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1692(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1693(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1694(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1359(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1360(.a(gate109inter0), .b(s_116), .O(gate109inter1));
  and2  gate1361(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1362(.a(s_116), .O(gate109inter3));
  inv1  gate1363(.a(s_117), .O(gate109inter4));
  nand2 gate1364(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1365(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1366(.a(G370), .O(gate109inter7));
  inv1  gate1367(.a(G371), .O(gate109inter8));
  nand2 gate1368(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1369(.a(s_117), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1370(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1371(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1372(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1163(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1164(.a(gate110inter0), .b(s_88), .O(gate110inter1));
  and2  gate1165(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1166(.a(s_88), .O(gate110inter3));
  inv1  gate1167(.a(s_89), .O(gate110inter4));
  nand2 gate1168(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1169(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1170(.a(G372), .O(gate110inter7));
  inv1  gate1171(.a(G373), .O(gate110inter8));
  nand2 gate1172(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1173(.a(s_89), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1174(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1175(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1176(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1667(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1668(.a(gate119inter0), .b(s_160), .O(gate119inter1));
  and2  gate1669(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1670(.a(s_160), .O(gate119inter3));
  inv1  gate1671(.a(s_161), .O(gate119inter4));
  nand2 gate1672(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1673(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1674(.a(G390), .O(gate119inter7));
  inv1  gate1675(.a(G391), .O(gate119inter8));
  nand2 gate1676(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1677(.a(s_161), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1678(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1679(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1680(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate981(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate982(.a(gate122inter0), .b(s_62), .O(gate122inter1));
  and2  gate983(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate984(.a(s_62), .O(gate122inter3));
  inv1  gate985(.a(s_63), .O(gate122inter4));
  nand2 gate986(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate987(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate988(.a(G396), .O(gate122inter7));
  inv1  gate989(.a(G397), .O(gate122inter8));
  nand2 gate990(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate991(.a(s_63), .b(gate122inter3), .O(gate122inter10));
  nor2  gate992(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate993(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate994(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1555(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1556(.a(gate125inter0), .b(s_144), .O(gate125inter1));
  and2  gate1557(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1558(.a(s_144), .O(gate125inter3));
  inv1  gate1559(.a(s_145), .O(gate125inter4));
  nand2 gate1560(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1561(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1562(.a(G402), .O(gate125inter7));
  inv1  gate1563(.a(G403), .O(gate125inter8));
  nand2 gate1564(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1565(.a(s_145), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1566(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1567(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1568(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1149(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1150(.a(gate137inter0), .b(s_86), .O(gate137inter1));
  and2  gate1151(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1152(.a(s_86), .O(gate137inter3));
  inv1  gate1153(.a(s_87), .O(gate137inter4));
  nand2 gate1154(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1155(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1156(.a(G426), .O(gate137inter7));
  inv1  gate1157(.a(G429), .O(gate137inter8));
  nand2 gate1158(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1159(.a(s_87), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1160(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1161(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1162(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1079(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1080(.a(gate139inter0), .b(s_76), .O(gate139inter1));
  and2  gate1081(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1082(.a(s_76), .O(gate139inter3));
  inv1  gate1083(.a(s_77), .O(gate139inter4));
  nand2 gate1084(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1085(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1086(.a(G438), .O(gate139inter7));
  inv1  gate1087(.a(G441), .O(gate139inter8));
  nand2 gate1088(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1089(.a(s_77), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1090(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1091(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1092(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1653(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1654(.a(gate142inter0), .b(s_158), .O(gate142inter1));
  and2  gate1655(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1656(.a(s_158), .O(gate142inter3));
  inv1  gate1657(.a(s_159), .O(gate142inter4));
  nand2 gate1658(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1659(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1660(.a(G456), .O(gate142inter7));
  inv1  gate1661(.a(G459), .O(gate142inter8));
  nand2 gate1662(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1663(.a(s_159), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1664(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1665(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1666(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1457(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1458(.a(gate145inter0), .b(s_130), .O(gate145inter1));
  and2  gate1459(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1460(.a(s_130), .O(gate145inter3));
  inv1  gate1461(.a(s_131), .O(gate145inter4));
  nand2 gate1462(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1463(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1464(.a(G474), .O(gate145inter7));
  inv1  gate1465(.a(G477), .O(gate145inter8));
  nand2 gate1466(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1467(.a(s_131), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1468(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1469(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1470(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1065(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1066(.a(gate158inter0), .b(s_74), .O(gate158inter1));
  and2  gate1067(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1068(.a(s_74), .O(gate158inter3));
  inv1  gate1069(.a(s_75), .O(gate158inter4));
  nand2 gate1070(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1071(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1072(.a(G441), .O(gate158inter7));
  inv1  gate1073(.a(G528), .O(gate158inter8));
  nand2 gate1074(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1075(.a(s_75), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1076(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1077(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1078(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate561(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate562(.a(gate160inter0), .b(s_2), .O(gate160inter1));
  and2  gate563(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate564(.a(s_2), .O(gate160inter3));
  inv1  gate565(.a(s_3), .O(gate160inter4));
  nand2 gate566(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate567(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate568(.a(G447), .O(gate160inter7));
  inv1  gate569(.a(G531), .O(gate160inter8));
  nand2 gate570(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate571(.a(s_3), .b(gate160inter3), .O(gate160inter10));
  nor2  gate572(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate573(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate574(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate673(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate674(.a(gate162inter0), .b(s_18), .O(gate162inter1));
  and2  gate675(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate676(.a(s_18), .O(gate162inter3));
  inv1  gate677(.a(s_19), .O(gate162inter4));
  nand2 gate678(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate679(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate680(.a(G453), .O(gate162inter7));
  inv1  gate681(.a(G534), .O(gate162inter8));
  nand2 gate682(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate683(.a(s_19), .b(gate162inter3), .O(gate162inter10));
  nor2  gate684(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate685(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate686(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1037(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1038(.a(gate164inter0), .b(s_70), .O(gate164inter1));
  and2  gate1039(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1040(.a(s_70), .O(gate164inter3));
  inv1  gate1041(.a(s_71), .O(gate164inter4));
  nand2 gate1042(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1043(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1044(.a(G459), .O(gate164inter7));
  inv1  gate1045(.a(G537), .O(gate164inter8));
  nand2 gate1046(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1047(.a(s_71), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1048(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1049(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1050(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1415(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1416(.a(gate174inter0), .b(s_124), .O(gate174inter1));
  and2  gate1417(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1418(.a(s_124), .O(gate174inter3));
  inv1  gate1419(.a(s_125), .O(gate174inter4));
  nand2 gate1420(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1421(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1422(.a(G489), .O(gate174inter7));
  inv1  gate1423(.a(G552), .O(gate174inter8));
  nand2 gate1424(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1425(.a(s_125), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1426(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1427(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1428(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1219(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1220(.a(gate177inter0), .b(s_96), .O(gate177inter1));
  and2  gate1221(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1222(.a(s_96), .O(gate177inter3));
  inv1  gate1223(.a(s_97), .O(gate177inter4));
  nand2 gate1224(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1225(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1226(.a(G498), .O(gate177inter7));
  inv1  gate1227(.a(G558), .O(gate177inter8));
  nand2 gate1228(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1229(.a(s_97), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1230(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1231(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1232(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate757(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate758(.a(gate178inter0), .b(s_30), .O(gate178inter1));
  and2  gate759(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate760(.a(s_30), .O(gate178inter3));
  inv1  gate761(.a(s_31), .O(gate178inter4));
  nand2 gate762(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate763(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate764(.a(G501), .O(gate178inter7));
  inv1  gate765(.a(G558), .O(gate178inter8));
  nand2 gate766(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate767(.a(s_31), .b(gate178inter3), .O(gate178inter10));
  nor2  gate768(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate769(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate770(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1723(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1724(.a(gate181inter0), .b(s_168), .O(gate181inter1));
  and2  gate1725(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1726(.a(s_168), .O(gate181inter3));
  inv1  gate1727(.a(s_169), .O(gate181inter4));
  nand2 gate1728(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1729(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1730(.a(G510), .O(gate181inter7));
  inv1  gate1731(.a(G564), .O(gate181inter8));
  nand2 gate1732(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1733(.a(s_169), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1734(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1735(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1736(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1737(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1738(.a(gate182inter0), .b(s_170), .O(gate182inter1));
  and2  gate1739(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1740(.a(s_170), .O(gate182inter3));
  inv1  gate1741(.a(s_171), .O(gate182inter4));
  nand2 gate1742(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1743(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1744(.a(G513), .O(gate182inter7));
  inv1  gate1745(.a(G564), .O(gate182inter8));
  nand2 gate1746(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1747(.a(s_171), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1748(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1749(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1750(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate883(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate884(.a(gate191inter0), .b(s_48), .O(gate191inter1));
  and2  gate885(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate886(.a(s_48), .O(gate191inter3));
  inv1  gate887(.a(s_49), .O(gate191inter4));
  nand2 gate888(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate889(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate890(.a(G582), .O(gate191inter7));
  inv1  gate891(.a(G583), .O(gate191inter8));
  nand2 gate892(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate893(.a(s_49), .b(gate191inter3), .O(gate191inter10));
  nor2  gate894(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate895(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate896(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1289(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1290(.a(gate192inter0), .b(s_106), .O(gate192inter1));
  and2  gate1291(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1292(.a(s_106), .O(gate192inter3));
  inv1  gate1293(.a(s_107), .O(gate192inter4));
  nand2 gate1294(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1295(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1296(.a(G584), .O(gate192inter7));
  inv1  gate1297(.a(G585), .O(gate192inter8));
  nand2 gate1298(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1299(.a(s_107), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1300(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1301(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1302(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate939(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate940(.a(gate209inter0), .b(s_56), .O(gate209inter1));
  and2  gate941(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate942(.a(s_56), .O(gate209inter3));
  inv1  gate943(.a(s_57), .O(gate209inter4));
  nand2 gate944(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate945(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate946(.a(G602), .O(gate209inter7));
  inv1  gate947(.a(G666), .O(gate209inter8));
  nand2 gate948(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate949(.a(s_57), .b(gate209inter3), .O(gate209inter10));
  nor2  gate950(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate951(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate952(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate967(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate968(.a(gate211inter0), .b(s_60), .O(gate211inter1));
  and2  gate969(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate970(.a(s_60), .O(gate211inter3));
  inv1  gate971(.a(s_61), .O(gate211inter4));
  nand2 gate972(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate973(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate974(.a(G612), .O(gate211inter7));
  inv1  gate975(.a(G669), .O(gate211inter8));
  nand2 gate976(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate977(.a(s_61), .b(gate211inter3), .O(gate211inter10));
  nor2  gate978(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate979(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate980(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate743(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate744(.a(gate236inter0), .b(s_28), .O(gate236inter1));
  and2  gate745(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate746(.a(s_28), .O(gate236inter3));
  inv1  gate747(.a(s_29), .O(gate236inter4));
  nand2 gate748(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate749(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate750(.a(G251), .O(gate236inter7));
  inv1  gate751(.a(G727), .O(gate236inter8));
  nand2 gate752(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate753(.a(s_29), .b(gate236inter3), .O(gate236inter10));
  nor2  gate754(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate755(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate756(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1625(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1626(.a(gate237inter0), .b(s_154), .O(gate237inter1));
  and2  gate1627(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1628(.a(s_154), .O(gate237inter3));
  inv1  gate1629(.a(s_155), .O(gate237inter4));
  nand2 gate1630(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1631(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1632(.a(G254), .O(gate237inter7));
  inv1  gate1633(.a(G706), .O(gate237inter8));
  nand2 gate1634(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1635(.a(s_155), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1636(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1637(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1638(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1135(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1136(.a(gate253inter0), .b(s_84), .O(gate253inter1));
  and2  gate1137(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1138(.a(s_84), .O(gate253inter3));
  inv1  gate1139(.a(s_85), .O(gate253inter4));
  nand2 gate1140(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1141(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1142(.a(G260), .O(gate253inter7));
  inv1  gate1143(.a(G748), .O(gate253inter8));
  nand2 gate1144(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1145(.a(s_85), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1146(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1147(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1148(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate953(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate954(.a(gate257inter0), .b(s_58), .O(gate257inter1));
  and2  gate955(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate956(.a(s_58), .O(gate257inter3));
  inv1  gate957(.a(s_59), .O(gate257inter4));
  nand2 gate958(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate959(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate960(.a(G754), .O(gate257inter7));
  inv1  gate961(.a(G755), .O(gate257inter8));
  nand2 gate962(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate963(.a(s_59), .b(gate257inter3), .O(gate257inter10));
  nor2  gate964(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate965(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate966(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1695(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1696(.a(gate258inter0), .b(s_164), .O(gate258inter1));
  and2  gate1697(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1698(.a(s_164), .O(gate258inter3));
  inv1  gate1699(.a(s_165), .O(gate258inter4));
  nand2 gate1700(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1701(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1702(.a(G756), .O(gate258inter7));
  inv1  gate1703(.a(G757), .O(gate258inter8));
  nand2 gate1704(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1705(.a(s_165), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1706(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1707(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1708(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1107(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1108(.a(gate267inter0), .b(s_80), .O(gate267inter1));
  and2  gate1109(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1110(.a(s_80), .O(gate267inter3));
  inv1  gate1111(.a(s_81), .O(gate267inter4));
  nand2 gate1112(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1113(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1114(.a(G648), .O(gate267inter7));
  inv1  gate1115(.a(G776), .O(gate267inter8));
  nand2 gate1116(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1117(.a(s_81), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1118(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1119(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1120(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1345(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1346(.a(gate270inter0), .b(s_114), .O(gate270inter1));
  and2  gate1347(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1348(.a(s_114), .O(gate270inter3));
  inv1  gate1349(.a(s_115), .O(gate270inter4));
  nand2 gate1350(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1351(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1352(.a(G657), .O(gate270inter7));
  inv1  gate1353(.a(G785), .O(gate270inter8));
  nand2 gate1354(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1355(.a(s_115), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1356(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1357(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1358(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1499(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1500(.a(gate276inter0), .b(s_136), .O(gate276inter1));
  and2  gate1501(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1502(.a(s_136), .O(gate276inter3));
  inv1  gate1503(.a(s_137), .O(gate276inter4));
  nand2 gate1504(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1505(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1506(.a(G773), .O(gate276inter7));
  inv1  gate1507(.a(G797), .O(gate276inter8));
  nand2 gate1508(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1509(.a(s_137), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1510(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1511(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1512(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate715(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate716(.a(gate277inter0), .b(s_24), .O(gate277inter1));
  and2  gate717(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate718(.a(s_24), .O(gate277inter3));
  inv1  gate719(.a(s_25), .O(gate277inter4));
  nand2 gate720(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate721(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate722(.a(G648), .O(gate277inter7));
  inv1  gate723(.a(G800), .O(gate277inter8));
  nand2 gate724(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate725(.a(s_25), .b(gate277inter3), .O(gate277inter10));
  nor2  gate726(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate727(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate728(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate659(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate660(.a(gate283inter0), .b(s_16), .O(gate283inter1));
  and2  gate661(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate662(.a(s_16), .O(gate283inter3));
  inv1  gate663(.a(s_17), .O(gate283inter4));
  nand2 gate664(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate665(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate666(.a(G657), .O(gate283inter7));
  inv1  gate667(.a(G809), .O(gate283inter8));
  nand2 gate668(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate669(.a(s_17), .b(gate283inter3), .O(gate283inter10));
  nor2  gate670(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate671(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate672(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1639(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1640(.a(gate284inter0), .b(s_156), .O(gate284inter1));
  and2  gate1641(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1642(.a(s_156), .O(gate284inter3));
  inv1  gate1643(.a(s_157), .O(gate284inter4));
  nand2 gate1644(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1645(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1646(.a(G785), .O(gate284inter7));
  inv1  gate1647(.a(G809), .O(gate284inter8));
  nand2 gate1648(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1649(.a(s_157), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1650(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1651(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1652(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate771(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate772(.a(gate286inter0), .b(s_32), .O(gate286inter1));
  and2  gate773(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate774(.a(s_32), .O(gate286inter3));
  inv1  gate775(.a(s_33), .O(gate286inter4));
  nand2 gate776(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate777(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate778(.a(G788), .O(gate286inter7));
  inv1  gate779(.a(G812), .O(gate286inter8));
  nand2 gate780(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate781(.a(s_33), .b(gate286inter3), .O(gate286inter10));
  nor2  gate782(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate783(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate784(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate995(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate996(.a(gate291inter0), .b(s_64), .O(gate291inter1));
  and2  gate997(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate998(.a(s_64), .O(gate291inter3));
  inv1  gate999(.a(s_65), .O(gate291inter4));
  nand2 gate1000(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1001(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1002(.a(G822), .O(gate291inter7));
  inv1  gate1003(.a(G823), .O(gate291inter8));
  nand2 gate1004(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1005(.a(s_65), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1006(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1007(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1008(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate617(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate618(.a(gate294inter0), .b(s_10), .O(gate294inter1));
  and2  gate619(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate620(.a(s_10), .O(gate294inter3));
  inv1  gate621(.a(s_11), .O(gate294inter4));
  nand2 gate622(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate623(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate624(.a(G832), .O(gate294inter7));
  inv1  gate625(.a(G833), .O(gate294inter8));
  nand2 gate626(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate627(.a(s_11), .b(gate294inter3), .O(gate294inter10));
  nor2  gate628(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate629(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate630(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate841(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate842(.a(gate389inter0), .b(s_42), .O(gate389inter1));
  and2  gate843(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate844(.a(s_42), .O(gate389inter3));
  inv1  gate845(.a(s_43), .O(gate389inter4));
  nand2 gate846(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate847(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate848(.a(G3), .O(gate389inter7));
  inv1  gate849(.a(G1042), .O(gate389inter8));
  nand2 gate850(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate851(.a(s_43), .b(gate389inter3), .O(gate389inter10));
  nor2  gate852(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate853(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate854(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1807(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1808(.a(gate394inter0), .b(s_180), .O(gate394inter1));
  and2  gate1809(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1810(.a(s_180), .O(gate394inter3));
  inv1  gate1811(.a(s_181), .O(gate394inter4));
  nand2 gate1812(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1813(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1814(.a(G8), .O(gate394inter7));
  inv1  gate1815(.a(G1057), .O(gate394inter8));
  nand2 gate1816(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1817(.a(s_181), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1818(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1819(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1820(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1429(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1430(.a(gate395inter0), .b(s_126), .O(gate395inter1));
  and2  gate1431(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1432(.a(s_126), .O(gate395inter3));
  inv1  gate1433(.a(s_127), .O(gate395inter4));
  nand2 gate1434(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1435(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1436(.a(G9), .O(gate395inter7));
  inv1  gate1437(.a(G1060), .O(gate395inter8));
  nand2 gate1438(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1439(.a(s_127), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1440(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1441(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1442(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1177(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1178(.a(gate398inter0), .b(s_90), .O(gate398inter1));
  and2  gate1179(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1180(.a(s_90), .O(gate398inter3));
  inv1  gate1181(.a(s_91), .O(gate398inter4));
  nand2 gate1182(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1183(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1184(.a(G12), .O(gate398inter7));
  inv1  gate1185(.a(G1069), .O(gate398inter8));
  nand2 gate1186(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1187(.a(s_91), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1188(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1189(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1190(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate701(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate702(.a(gate399inter0), .b(s_22), .O(gate399inter1));
  and2  gate703(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate704(.a(s_22), .O(gate399inter3));
  inv1  gate705(.a(s_23), .O(gate399inter4));
  nand2 gate706(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate707(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate708(.a(G13), .O(gate399inter7));
  inv1  gate709(.a(G1072), .O(gate399inter8));
  nand2 gate710(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate711(.a(s_23), .b(gate399inter3), .O(gate399inter10));
  nor2  gate712(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate713(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate714(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1541(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1542(.a(gate411inter0), .b(s_142), .O(gate411inter1));
  and2  gate1543(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1544(.a(s_142), .O(gate411inter3));
  inv1  gate1545(.a(s_143), .O(gate411inter4));
  nand2 gate1546(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1547(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1548(.a(G25), .O(gate411inter7));
  inv1  gate1549(.a(G1108), .O(gate411inter8));
  nand2 gate1550(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1551(.a(s_143), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1552(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1553(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1554(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1793(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1794(.a(gate413inter0), .b(s_178), .O(gate413inter1));
  and2  gate1795(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1796(.a(s_178), .O(gate413inter3));
  inv1  gate1797(.a(s_179), .O(gate413inter4));
  nand2 gate1798(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1799(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1800(.a(G27), .O(gate413inter7));
  inv1  gate1801(.a(G1114), .O(gate413inter8));
  nand2 gate1802(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1803(.a(s_179), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1804(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1805(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1806(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate925(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate926(.a(gate418inter0), .b(s_54), .O(gate418inter1));
  and2  gate927(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate928(.a(s_54), .O(gate418inter3));
  inv1  gate929(.a(s_55), .O(gate418inter4));
  nand2 gate930(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate931(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate932(.a(G32), .O(gate418inter7));
  inv1  gate933(.a(G1129), .O(gate418inter8));
  nand2 gate934(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate935(.a(s_55), .b(gate418inter3), .O(gate418inter10));
  nor2  gate936(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate937(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate938(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1009(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1010(.a(gate420inter0), .b(s_66), .O(gate420inter1));
  and2  gate1011(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1012(.a(s_66), .O(gate420inter3));
  inv1  gate1013(.a(s_67), .O(gate420inter4));
  nand2 gate1014(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1015(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1016(.a(G1036), .O(gate420inter7));
  inv1  gate1017(.a(G1132), .O(gate420inter8));
  nand2 gate1018(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1019(.a(s_67), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1020(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1021(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1022(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1387(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1388(.a(gate424inter0), .b(s_120), .O(gate424inter1));
  and2  gate1389(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1390(.a(s_120), .O(gate424inter3));
  inv1  gate1391(.a(s_121), .O(gate424inter4));
  nand2 gate1392(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1393(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1394(.a(G1042), .O(gate424inter7));
  inv1  gate1395(.a(G1138), .O(gate424inter8));
  nand2 gate1396(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1397(.a(s_121), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1398(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1399(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1400(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1247(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1248(.a(gate427inter0), .b(s_100), .O(gate427inter1));
  and2  gate1249(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1250(.a(s_100), .O(gate427inter3));
  inv1  gate1251(.a(s_101), .O(gate427inter4));
  nand2 gate1252(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1253(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1254(.a(G5), .O(gate427inter7));
  inv1  gate1255(.a(G1144), .O(gate427inter8));
  nand2 gate1256(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1257(.a(s_101), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1258(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1259(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1260(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1317(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1318(.a(gate428inter0), .b(s_110), .O(gate428inter1));
  and2  gate1319(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1320(.a(s_110), .O(gate428inter3));
  inv1  gate1321(.a(s_111), .O(gate428inter4));
  nand2 gate1322(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1323(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1324(.a(G1048), .O(gate428inter7));
  inv1  gate1325(.a(G1144), .O(gate428inter8));
  nand2 gate1326(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1327(.a(s_111), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1328(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1329(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1330(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate897(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate898(.a(gate433inter0), .b(s_50), .O(gate433inter1));
  and2  gate899(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate900(.a(s_50), .O(gate433inter3));
  inv1  gate901(.a(s_51), .O(gate433inter4));
  nand2 gate902(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate903(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate904(.a(G8), .O(gate433inter7));
  inv1  gate905(.a(G1153), .O(gate433inter8));
  nand2 gate906(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate907(.a(s_51), .b(gate433inter3), .O(gate433inter10));
  nor2  gate908(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate909(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate910(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1275(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1276(.a(gate440inter0), .b(s_104), .O(gate440inter1));
  and2  gate1277(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1278(.a(s_104), .O(gate440inter3));
  inv1  gate1279(.a(s_105), .O(gate440inter4));
  nand2 gate1280(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1281(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1282(.a(G1066), .O(gate440inter7));
  inv1  gate1283(.a(G1162), .O(gate440inter8));
  nand2 gate1284(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1285(.a(s_105), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1286(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1287(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1288(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate855(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate856(.a(gate446inter0), .b(s_44), .O(gate446inter1));
  and2  gate857(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate858(.a(s_44), .O(gate446inter3));
  inv1  gate859(.a(s_45), .O(gate446inter4));
  nand2 gate860(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate861(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate862(.a(G1075), .O(gate446inter7));
  inv1  gate863(.a(G1171), .O(gate446inter8));
  nand2 gate864(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate865(.a(s_45), .b(gate446inter3), .O(gate446inter10));
  nor2  gate866(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate867(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate868(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1485(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1486(.a(gate447inter0), .b(s_134), .O(gate447inter1));
  and2  gate1487(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1488(.a(s_134), .O(gate447inter3));
  inv1  gate1489(.a(s_135), .O(gate447inter4));
  nand2 gate1490(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1491(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1492(.a(G15), .O(gate447inter7));
  inv1  gate1493(.a(G1174), .O(gate447inter8));
  nand2 gate1494(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1495(.a(s_135), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1496(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1497(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1498(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate911(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate912(.a(gate452inter0), .b(s_52), .O(gate452inter1));
  and2  gate913(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate914(.a(s_52), .O(gate452inter3));
  inv1  gate915(.a(s_53), .O(gate452inter4));
  nand2 gate916(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate917(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate918(.a(G1084), .O(gate452inter7));
  inv1  gate919(.a(G1180), .O(gate452inter8));
  nand2 gate920(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate921(.a(s_53), .b(gate452inter3), .O(gate452inter10));
  nor2  gate922(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate923(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate924(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1233(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1234(.a(gate455inter0), .b(s_98), .O(gate455inter1));
  and2  gate1235(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1236(.a(s_98), .O(gate455inter3));
  inv1  gate1237(.a(s_99), .O(gate455inter4));
  nand2 gate1238(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1239(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1240(.a(G19), .O(gate455inter7));
  inv1  gate1241(.a(G1186), .O(gate455inter8));
  nand2 gate1242(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1243(.a(s_99), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1244(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1245(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1246(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1121(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1122(.a(gate457inter0), .b(s_82), .O(gate457inter1));
  and2  gate1123(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1124(.a(s_82), .O(gate457inter3));
  inv1  gate1125(.a(s_83), .O(gate457inter4));
  nand2 gate1126(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1127(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1128(.a(G20), .O(gate457inter7));
  inv1  gate1129(.a(G1189), .O(gate457inter8));
  nand2 gate1130(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1131(.a(s_83), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1132(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1133(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1134(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1583(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1584(.a(gate458inter0), .b(s_148), .O(gate458inter1));
  and2  gate1585(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1586(.a(s_148), .O(gate458inter3));
  inv1  gate1587(.a(s_149), .O(gate458inter4));
  nand2 gate1588(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1589(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1590(.a(G1093), .O(gate458inter7));
  inv1  gate1591(.a(G1189), .O(gate458inter8));
  nand2 gate1592(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1593(.a(s_149), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1594(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1595(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1596(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1401(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1402(.a(gate465inter0), .b(s_122), .O(gate465inter1));
  and2  gate1403(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1404(.a(s_122), .O(gate465inter3));
  inv1  gate1405(.a(s_123), .O(gate465inter4));
  nand2 gate1406(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1407(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1408(.a(G24), .O(gate465inter7));
  inv1  gate1409(.a(G1201), .O(gate465inter8));
  nand2 gate1410(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1411(.a(s_123), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1412(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1413(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1414(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1303(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1304(.a(gate470inter0), .b(s_108), .O(gate470inter1));
  and2  gate1305(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1306(.a(s_108), .O(gate470inter3));
  inv1  gate1307(.a(s_109), .O(gate470inter4));
  nand2 gate1308(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1309(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1310(.a(G1111), .O(gate470inter7));
  inv1  gate1311(.a(G1207), .O(gate470inter8));
  nand2 gate1312(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1313(.a(s_109), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1314(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1315(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1316(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate603(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate604(.a(gate472inter0), .b(s_8), .O(gate472inter1));
  and2  gate605(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate606(.a(s_8), .O(gate472inter3));
  inv1  gate607(.a(s_9), .O(gate472inter4));
  nand2 gate608(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate609(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate610(.a(G1114), .O(gate472inter7));
  inv1  gate611(.a(G1210), .O(gate472inter8));
  nand2 gate612(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate613(.a(s_9), .b(gate472inter3), .O(gate472inter10));
  nor2  gate614(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate615(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate616(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1191(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1192(.a(gate481inter0), .b(s_92), .O(gate481inter1));
  and2  gate1193(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1194(.a(s_92), .O(gate481inter3));
  inv1  gate1195(.a(s_93), .O(gate481inter4));
  nand2 gate1196(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1197(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1198(.a(G32), .O(gate481inter7));
  inv1  gate1199(.a(G1225), .O(gate481inter8));
  nand2 gate1200(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1201(.a(s_93), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1202(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1203(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1204(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1751(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1752(.a(gate498inter0), .b(s_172), .O(gate498inter1));
  and2  gate1753(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1754(.a(s_172), .O(gate498inter3));
  inv1  gate1755(.a(s_173), .O(gate498inter4));
  nand2 gate1756(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1757(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1758(.a(G1258), .O(gate498inter7));
  inv1  gate1759(.a(G1259), .O(gate498inter8));
  nand2 gate1760(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1761(.a(s_173), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1762(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1763(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1764(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate799(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate800(.a(gate501inter0), .b(s_36), .O(gate501inter1));
  and2  gate801(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate802(.a(s_36), .O(gate501inter3));
  inv1  gate803(.a(s_37), .O(gate501inter4));
  nand2 gate804(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate805(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate806(.a(G1264), .O(gate501inter7));
  inv1  gate807(.a(G1265), .O(gate501inter8));
  nand2 gate808(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate809(.a(s_37), .b(gate501inter3), .O(gate501inter10));
  nor2  gate810(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate811(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate812(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1443(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1444(.a(gate506inter0), .b(s_128), .O(gate506inter1));
  and2  gate1445(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1446(.a(s_128), .O(gate506inter3));
  inv1  gate1447(.a(s_129), .O(gate506inter4));
  nand2 gate1448(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1449(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1450(.a(G1274), .O(gate506inter7));
  inv1  gate1451(.a(G1275), .O(gate506inter8));
  nand2 gate1452(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1453(.a(s_129), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1454(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1455(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1456(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate645(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate646(.a(gate514inter0), .b(s_14), .O(gate514inter1));
  and2  gate647(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate648(.a(s_14), .O(gate514inter3));
  inv1  gate649(.a(s_15), .O(gate514inter4));
  nand2 gate650(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate651(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate652(.a(G1290), .O(gate514inter7));
  inv1  gate653(.a(G1291), .O(gate514inter8));
  nand2 gate654(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate655(.a(s_15), .b(gate514inter3), .O(gate514inter10));
  nor2  gate656(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate657(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate658(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule