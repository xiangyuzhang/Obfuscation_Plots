module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate575(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate576(.a(gate9inter0), .b(s_4), .O(gate9inter1));
  and2  gate577(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate578(.a(s_4), .O(gate9inter3));
  inv1  gate579(.a(s_5), .O(gate9inter4));
  nand2 gate580(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate581(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate582(.a(G1), .O(gate9inter7));
  inv1  gate583(.a(G2), .O(gate9inter8));
  nand2 gate584(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate585(.a(s_5), .b(gate9inter3), .O(gate9inter10));
  nor2  gate586(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate587(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate588(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1373(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1374(.a(gate21inter0), .b(s_118), .O(gate21inter1));
  and2  gate1375(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1376(.a(s_118), .O(gate21inter3));
  inv1  gate1377(.a(s_119), .O(gate21inter4));
  nand2 gate1378(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1379(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1380(.a(G25), .O(gate21inter7));
  inv1  gate1381(.a(G26), .O(gate21inter8));
  nand2 gate1382(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1383(.a(s_119), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1384(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1385(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1386(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1205(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1206(.a(gate26inter0), .b(s_94), .O(gate26inter1));
  and2  gate1207(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1208(.a(s_94), .O(gate26inter3));
  inv1  gate1209(.a(s_95), .O(gate26inter4));
  nand2 gate1210(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1211(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1212(.a(G9), .O(gate26inter7));
  inv1  gate1213(.a(G13), .O(gate26inter8));
  nand2 gate1214(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1215(.a(s_95), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1216(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1217(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1218(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate827(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate828(.a(gate30inter0), .b(s_40), .O(gate30inter1));
  and2  gate829(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate830(.a(s_40), .O(gate30inter3));
  inv1  gate831(.a(s_41), .O(gate30inter4));
  nand2 gate832(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate833(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate834(.a(G11), .O(gate30inter7));
  inv1  gate835(.a(G15), .O(gate30inter8));
  nand2 gate836(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate837(.a(s_41), .b(gate30inter3), .O(gate30inter10));
  nor2  gate838(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate839(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate840(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate771(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate772(.a(gate31inter0), .b(s_32), .O(gate31inter1));
  and2  gate773(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate774(.a(s_32), .O(gate31inter3));
  inv1  gate775(.a(s_33), .O(gate31inter4));
  nand2 gate776(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate777(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate778(.a(G4), .O(gate31inter7));
  inv1  gate779(.a(G8), .O(gate31inter8));
  nand2 gate780(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate781(.a(s_33), .b(gate31inter3), .O(gate31inter10));
  nor2  gate782(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate783(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate784(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate911(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate912(.a(gate38inter0), .b(s_52), .O(gate38inter1));
  and2  gate913(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate914(.a(s_52), .O(gate38inter3));
  inv1  gate915(.a(s_53), .O(gate38inter4));
  nand2 gate916(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate917(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate918(.a(G27), .O(gate38inter7));
  inv1  gate919(.a(G31), .O(gate38inter8));
  nand2 gate920(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate921(.a(s_53), .b(gate38inter3), .O(gate38inter10));
  nor2  gate922(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate923(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate924(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1107(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1108(.a(gate41inter0), .b(s_80), .O(gate41inter1));
  and2  gate1109(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1110(.a(s_80), .O(gate41inter3));
  inv1  gate1111(.a(s_81), .O(gate41inter4));
  nand2 gate1112(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1113(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1114(.a(G1), .O(gate41inter7));
  inv1  gate1115(.a(G266), .O(gate41inter8));
  nand2 gate1116(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1117(.a(s_81), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1118(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1119(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1120(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate547(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate548(.a(gate43inter0), .b(s_0), .O(gate43inter1));
  and2  gate549(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate550(.a(s_0), .O(gate43inter3));
  inv1  gate551(.a(s_1), .O(gate43inter4));
  nand2 gate552(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate553(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate554(.a(G3), .O(gate43inter7));
  inv1  gate555(.a(G269), .O(gate43inter8));
  nand2 gate556(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate557(.a(s_1), .b(gate43inter3), .O(gate43inter10));
  nor2  gate558(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate559(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate560(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate855(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate856(.a(gate44inter0), .b(s_44), .O(gate44inter1));
  and2  gate857(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate858(.a(s_44), .O(gate44inter3));
  inv1  gate859(.a(s_45), .O(gate44inter4));
  nand2 gate860(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate861(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate862(.a(G4), .O(gate44inter7));
  inv1  gate863(.a(G269), .O(gate44inter8));
  nand2 gate864(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate865(.a(s_45), .b(gate44inter3), .O(gate44inter10));
  nor2  gate866(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate867(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate868(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate701(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate702(.a(gate57inter0), .b(s_22), .O(gate57inter1));
  and2  gate703(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate704(.a(s_22), .O(gate57inter3));
  inv1  gate705(.a(s_23), .O(gate57inter4));
  nand2 gate706(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate707(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate708(.a(G17), .O(gate57inter7));
  inv1  gate709(.a(G290), .O(gate57inter8));
  nand2 gate710(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate711(.a(s_23), .b(gate57inter3), .O(gate57inter10));
  nor2  gate712(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate713(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate714(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1121(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1122(.a(gate58inter0), .b(s_82), .O(gate58inter1));
  and2  gate1123(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1124(.a(s_82), .O(gate58inter3));
  inv1  gate1125(.a(s_83), .O(gate58inter4));
  nand2 gate1126(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1127(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1128(.a(G18), .O(gate58inter7));
  inv1  gate1129(.a(G290), .O(gate58inter8));
  nand2 gate1130(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1131(.a(s_83), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1132(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1133(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1134(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1415(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1416(.a(gate80inter0), .b(s_124), .O(gate80inter1));
  and2  gate1417(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1418(.a(s_124), .O(gate80inter3));
  inv1  gate1419(.a(s_125), .O(gate80inter4));
  nand2 gate1420(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1421(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1422(.a(G14), .O(gate80inter7));
  inv1  gate1423(.a(G323), .O(gate80inter8));
  nand2 gate1424(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1425(.a(s_125), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1426(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1427(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1428(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1163(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1164(.a(gate81inter0), .b(s_88), .O(gate81inter1));
  and2  gate1165(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1166(.a(s_88), .O(gate81inter3));
  inv1  gate1167(.a(s_89), .O(gate81inter4));
  nand2 gate1168(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1169(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1170(.a(G3), .O(gate81inter7));
  inv1  gate1171(.a(G326), .O(gate81inter8));
  nand2 gate1172(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1173(.a(s_89), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1174(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1175(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1176(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1303(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1304(.a(gate94inter0), .b(s_108), .O(gate94inter1));
  and2  gate1305(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1306(.a(s_108), .O(gate94inter3));
  inv1  gate1307(.a(s_109), .O(gate94inter4));
  nand2 gate1308(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1309(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1310(.a(G22), .O(gate94inter7));
  inv1  gate1311(.a(G344), .O(gate94inter8));
  nand2 gate1312(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1313(.a(s_109), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1314(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1315(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1316(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1065(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1066(.a(gate104inter0), .b(s_74), .O(gate104inter1));
  and2  gate1067(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1068(.a(s_74), .O(gate104inter3));
  inv1  gate1069(.a(s_75), .O(gate104inter4));
  nand2 gate1070(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1071(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1072(.a(G32), .O(gate104inter7));
  inv1  gate1073(.a(G359), .O(gate104inter8));
  nand2 gate1074(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1075(.a(s_75), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1076(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1077(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1078(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate813(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate814(.a(gate107inter0), .b(s_38), .O(gate107inter1));
  and2  gate815(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate816(.a(s_38), .O(gate107inter3));
  inv1  gate817(.a(s_39), .O(gate107inter4));
  nand2 gate818(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate819(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate820(.a(G366), .O(gate107inter7));
  inv1  gate821(.a(G367), .O(gate107inter8));
  nand2 gate822(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate823(.a(s_39), .b(gate107inter3), .O(gate107inter10));
  nor2  gate824(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate825(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate826(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1037(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1038(.a(gate108inter0), .b(s_70), .O(gate108inter1));
  and2  gate1039(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1040(.a(s_70), .O(gate108inter3));
  inv1  gate1041(.a(s_71), .O(gate108inter4));
  nand2 gate1042(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1043(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1044(.a(G368), .O(gate108inter7));
  inv1  gate1045(.a(G369), .O(gate108inter8));
  nand2 gate1046(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1047(.a(s_71), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1048(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1049(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1050(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1499(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1500(.a(gate116inter0), .b(s_136), .O(gate116inter1));
  and2  gate1501(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1502(.a(s_136), .O(gate116inter3));
  inv1  gate1503(.a(s_137), .O(gate116inter4));
  nand2 gate1504(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1505(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1506(.a(G384), .O(gate116inter7));
  inv1  gate1507(.a(G385), .O(gate116inter8));
  nand2 gate1508(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1509(.a(s_137), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1510(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1511(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1512(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate785(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate786(.a(gate117inter0), .b(s_34), .O(gate117inter1));
  and2  gate787(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate788(.a(s_34), .O(gate117inter3));
  inv1  gate789(.a(s_35), .O(gate117inter4));
  nand2 gate790(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate791(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate792(.a(G386), .O(gate117inter7));
  inv1  gate793(.a(G387), .O(gate117inter8));
  nand2 gate794(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate795(.a(s_35), .b(gate117inter3), .O(gate117inter10));
  nor2  gate796(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate797(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate798(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1471(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1472(.a(gate124inter0), .b(s_132), .O(gate124inter1));
  and2  gate1473(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1474(.a(s_132), .O(gate124inter3));
  inv1  gate1475(.a(s_133), .O(gate124inter4));
  nand2 gate1476(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1477(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1478(.a(G400), .O(gate124inter7));
  inv1  gate1479(.a(G401), .O(gate124inter8));
  nand2 gate1480(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1481(.a(s_133), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1482(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1483(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1484(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1233(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1234(.a(gate135inter0), .b(s_98), .O(gate135inter1));
  and2  gate1235(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1236(.a(s_98), .O(gate135inter3));
  inv1  gate1237(.a(s_99), .O(gate135inter4));
  nand2 gate1238(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1239(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1240(.a(G422), .O(gate135inter7));
  inv1  gate1241(.a(G423), .O(gate135inter8));
  nand2 gate1242(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1243(.a(s_99), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1244(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1245(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1246(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate757(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate758(.a(gate149inter0), .b(s_30), .O(gate149inter1));
  and2  gate759(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate760(.a(s_30), .O(gate149inter3));
  inv1  gate761(.a(s_31), .O(gate149inter4));
  nand2 gate762(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate763(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate764(.a(G498), .O(gate149inter7));
  inv1  gate765(.a(G501), .O(gate149inter8));
  nand2 gate766(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate767(.a(s_31), .b(gate149inter3), .O(gate149inter10));
  nor2  gate768(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate769(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate770(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1359(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1360(.a(gate154inter0), .b(s_116), .O(gate154inter1));
  and2  gate1361(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1362(.a(s_116), .O(gate154inter3));
  inv1  gate1363(.a(s_117), .O(gate154inter4));
  nand2 gate1364(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1365(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1366(.a(G429), .O(gate154inter7));
  inv1  gate1367(.a(G522), .O(gate154inter8));
  nand2 gate1368(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1369(.a(s_117), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1370(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1371(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1372(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate729(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate730(.a(gate155inter0), .b(s_26), .O(gate155inter1));
  and2  gate731(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate732(.a(s_26), .O(gate155inter3));
  inv1  gate733(.a(s_27), .O(gate155inter4));
  nand2 gate734(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate735(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate736(.a(G432), .O(gate155inter7));
  inv1  gate737(.a(G525), .O(gate155inter8));
  nand2 gate738(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate739(.a(s_27), .b(gate155inter3), .O(gate155inter10));
  nor2  gate740(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate741(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate742(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate631(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate632(.a(gate161inter0), .b(s_12), .O(gate161inter1));
  and2  gate633(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate634(.a(s_12), .O(gate161inter3));
  inv1  gate635(.a(s_13), .O(gate161inter4));
  nand2 gate636(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate637(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate638(.a(G450), .O(gate161inter7));
  inv1  gate639(.a(G534), .O(gate161inter8));
  nand2 gate640(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate641(.a(s_13), .b(gate161inter3), .O(gate161inter10));
  nor2  gate642(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate643(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate644(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate841(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate842(.a(gate166inter0), .b(s_42), .O(gate166inter1));
  and2  gate843(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate844(.a(s_42), .O(gate166inter3));
  inv1  gate845(.a(s_43), .O(gate166inter4));
  nand2 gate846(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate847(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate848(.a(G465), .O(gate166inter7));
  inv1  gate849(.a(G540), .O(gate166inter8));
  nand2 gate850(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate851(.a(s_43), .b(gate166inter3), .O(gate166inter10));
  nor2  gate852(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate853(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate854(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate939(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate940(.a(gate171inter0), .b(s_56), .O(gate171inter1));
  and2  gate941(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate942(.a(s_56), .O(gate171inter3));
  inv1  gate943(.a(s_57), .O(gate171inter4));
  nand2 gate944(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate945(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate946(.a(G480), .O(gate171inter7));
  inv1  gate947(.a(G549), .O(gate171inter8));
  nand2 gate948(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate949(.a(s_57), .b(gate171inter3), .O(gate171inter10));
  nor2  gate950(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate951(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate952(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1135(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1136(.a(gate182inter0), .b(s_84), .O(gate182inter1));
  and2  gate1137(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1138(.a(s_84), .O(gate182inter3));
  inv1  gate1139(.a(s_85), .O(gate182inter4));
  nand2 gate1140(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1141(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1142(.a(G513), .O(gate182inter7));
  inv1  gate1143(.a(G564), .O(gate182inter8));
  nand2 gate1144(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1145(.a(s_85), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1146(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1147(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1148(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate799(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate800(.a(gate185inter0), .b(s_36), .O(gate185inter1));
  and2  gate801(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate802(.a(s_36), .O(gate185inter3));
  inv1  gate803(.a(s_37), .O(gate185inter4));
  nand2 gate804(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate805(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate806(.a(G570), .O(gate185inter7));
  inv1  gate807(.a(G571), .O(gate185inter8));
  nand2 gate808(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate809(.a(s_37), .b(gate185inter3), .O(gate185inter10));
  nor2  gate810(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate811(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate812(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1289(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1290(.a(gate186inter0), .b(s_106), .O(gate186inter1));
  and2  gate1291(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1292(.a(s_106), .O(gate186inter3));
  inv1  gate1293(.a(s_107), .O(gate186inter4));
  nand2 gate1294(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1295(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1296(.a(G572), .O(gate186inter7));
  inv1  gate1297(.a(G573), .O(gate186inter8));
  nand2 gate1298(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1299(.a(s_107), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1300(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1301(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1302(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1191(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1192(.a(gate190inter0), .b(s_92), .O(gate190inter1));
  and2  gate1193(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1194(.a(s_92), .O(gate190inter3));
  inv1  gate1195(.a(s_93), .O(gate190inter4));
  nand2 gate1196(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1197(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1198(.a(G580), .O(gate190inter7));
  inv1  gate1199(.a(G581), .O(gate190inter8));
  nand2 gate1200(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1201(.a(s_93), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1202(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1203(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1204(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate883(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate884(.a(gate192inter0), .b(s_48), .O(gate192inter1));
  and2  gate885(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate886(.a(s_48), .O(gate192inter3));
  inv1  gate887(.a(s_49), .O(gate192inter4));
  nand2 gate888(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate889(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate890(.a(G584), .O(gate192inter7));
  inv1  gate891(.a(G585), .O(gate192inter8));
  nand2 gate892(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate893(.a(s_49), .b(gate192inter3), .O(gate192inter10));
  nor2  gate894(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate895(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate896(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate617(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate618(.a(gate200inter0), .b(s_10), .O(gate200inter1));
  and2  gate619(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate620(.a(s_10), .O(gate200inter3));
  inv1  gate621(.a(s_11), .O(gate200inter4));
  nand2 gate622(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate623(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate624(.a(G600), .O(gate200inter7));
  inv1  gate625(.a(G601), .O(gate200inter8));
  nand2 gate626(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate627(.a(s_11), .b(gate200inter3), .O(gate200inter10));
  nor2  gate628(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate629(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate630(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1009(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1010(.a(gate203inter0), .b(s_66), .O(gate203inter1));
  and2  gate1011(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1012(.a(s_66), .O(gate203inter3));
  inv1  gate1013(.a(s_67), .O(gate203inter4));
  nand2 gate1014(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1015(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1016(.a(G602), .O(gate203inter7));
  inv1  gate1017(.a(G612), .O(gate203inter8));
  nand2 gate1018(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1019(.a(s_67), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1020(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1021(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1022(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1219(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1220(.a(gate205inter0), .b(s_96), .O(gate205inter1));
  and2  gate1221(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1222(.a(s_96), .O(gate205inter3));
  inv1  gate1223(.a(s_97), .O(gate205inter4));
  nand2 gate1224(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1225(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1226(.a(G622), .O(gate205inter7));
  inv1  gate1227(.a(G627), .O(gate205inter8));
  nand2 gate1228(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1229(.a(s_97), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1230(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1231(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1232(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate659(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate660(.a(gate210inter0), .b(s_16), .O(gate210inter1));
  and2  gate661(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate662(.a(s_16), .O(gate210inter3));
  inv1  gate663(.a(s_17), .O(gate210inter4));
  nand2 gate664(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate665(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate666(.a(G607), .O(gate210inter7));
  inv1  gate667(.a(G666), .O(gate210inter8));
  nand2 gate668(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate669(.a(s_17), .b(gate210inter3), .O(gate210inter10));
  nor2  gate670(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate671(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate672(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate967(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate968(.a(gate221inter0), .b(s_60), .O(gate221inter1));
  and2  gate969(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate970(.a(s_60), .O(gate221inter3));
  inv1  gate971(.a(s_61), .O(gate221inter4));
  nand2 gate972(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate973(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate974(.a(G622), .O(gate221inter7));
  inv1  gate975(.a(G684), .O(gate221inter8));
  nand2 gate976(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate977(.a(s_61), .b(gate221inter3), .O(gate221inter10));
  nor2  gate978(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate979(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate980(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate995(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate996(.a(gate233inter0), .b(s_64), .O(gate233inter1));
  and2  gate997(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate998(.a(s_64), .O(gate233inter3));
  inv1  gate999(.a(s_65), .O(gate233inter4));
  nand2 gate1000(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1001(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1002(.a(G242), .O(gate233inter7));
  inv1  gate1003(.a(G718), .O(gate233inter8));
  nand2 gate1004(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1005(.a(s_65), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1006(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1007(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1008(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate687(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate688(.a(gate236inter0), .b(s_20), .O(gate236inter1));
  and2  gate689(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate690(.a(s_20), .O(gate236inter3));
  inv1  gate691(.a(s_21), .O(gate236inter4));
  nand2 gate692(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate693(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate694(.a(G251), .O(gate236inter7));
  inv1  gate695(.a(G727), .O(gate236inter8));
  nand2 gate696(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate697(.a(s_21), .b(gate236inter3), .O(gate236inter10));
  nor2  gate698(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate699(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate700(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1345(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1346(.a(gate240inter0), .b(s_114), .O(gate240inter1));
  and2  gate1347(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1348(.a(s_114), .O(gate240inter3));
  inv1  gate1349(.a(s_115), .O(gate240inter4));
  nand2 gate1350(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1351(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1352(.a(G263), .O(gate240inter7));
  inv1  gate1353(.a(G715), .O(gate240inter8));
  nand2 gate1354(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1355(.a(s_115), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1356(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1357(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1358(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate589(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate590(.a(gate244inter0), .b(s_6), .O(gate244inter1));
  and2  gate591(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate592(.a(s_6), .O(gate244inter3));
  inv1  gate593(.a(s_7), .O(gate244inter4));
  nand2 gate594(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate595(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate596(.a(G721), .O(gate244inter7));
  inv1  gate597(.a(G733), .O(gate244inter8));
  nand2 gate598(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate599(.a(s_7), .b(gate244inter3), .O(gate244inter10));
  nor2  gate600(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate601(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate602(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate897(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate898(.a(gate253inter0), .b(s_50), .O(gate253inter1));
  and2  gate899(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate900(.a(s_50), .O(gate253inter3));
  inv1  gate901(.a(s_51), .O(gate253inter4));
  nand2 gate902(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate903(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate904(.a(G260), .O(gate253inter7));
  inv1  gate905(.a(G748), .O(gate253inter8));
  nand2 gate906(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate907(.a(s_51), .b(gate253inter3), .O(gate253inter10));
  nor2  gate908(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate909(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate910(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate981(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate982(.a(gate258inter0), .b(s_62), .O(gate258inter1));
  and2  gate983(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate984(.a(s_62), .O(gate258inter3));
  inv1  gate985(.a(s_63), .O(gate258inter4));
  nand2 gate986(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate987(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate988(.a(G756), .O(gate258inter7));
  inv1  gate989(.a(G757), .O(gate258inter8));
  nand2 gate990(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate991(.a(s_63), .b(gate258inter3), .O(gate258inter10));
  nor2  gate992(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate993(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate994(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate603(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate604(.a(gate263inter0), .b(s_8), .O(gate263inter1));
  and2  gate605(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate606(.a(s_8), .O(gate263inter3));
  inv1  gate607(.a(s_9), .O(gate263inter4));
  nand2 gate608(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate609(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate610(.a(G766), .O(gate263inter7));
  inv1  gate611(.a(G767), .O(gate263inter8));
  nand2 gate612(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate613(.a(s_9), .b(gate263inter3), .O(gate263inter10));
  nor2  gate614(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate615(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate616(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate673(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate674(.a(gate272inter0), .b(s_18), .O(gate272inter1));
  and2  gate675(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate676(.a(s_18), .O(gate272inter3));
  inv1  gate677(.a(s_19), .O(gate272inter4));
  nand2 gate678(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate679(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate680(.a(G663), .O(gate272inter7));
  inv1  gate681(.a(G791), .O(gate272inter8));
  nand2 gate682(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate683(.a(s_19), .b(gate272inter3), .O(gate272inter10));
  nor2  gate684(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate685(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate686(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1079(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1080(.a(gate282inter0), .b(s_76), .O(gate282inter1));
  and2  gate1081(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1082(.a(s_76), .O(gate282inter3));
  inv1  gate1083(.a(s_77), .O(gate282inter4));
  nand2 gate1084(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1085(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1086(.a(G782), .O(gate282inter7));
  inv1  gate1087(.a(G806), .O(gate282inter8));
  nand2 gate1088(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1089(.a(s_77), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1090(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1091(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1092(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1485(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1486(.a(gate291inter0), .b(s_134), .O(gate291inter1));
  and2  gate1487(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1488(.a(s_134), .O(gate291inter3));
  inv1  gate1489(.a(s_135), .O(gate291inter4));
  nand2 gate1490(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1491(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1492(.a(G822), .O(gate291inter7));
  inv1  gate1493(.a(G823), .O(gate291inter8));
  nand2 gate1494(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1495(.a(s_135), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1496(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1497(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1498(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1149(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1150(.a(gate296inter0), .b(s_86), .O(gate296inter1));
  and2  gate1151(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1152(.a(s_86), .O(gate296inter3));
  inv1  gate1153(.a(s_87), .O(gate296inter4));
  nand2 gate1154(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1155(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1156(.a(G826), .O(gate296inter7));
  inv1  gate1157(.a(G827), .O(gate296inter8));
  nand2 gate1158(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1159(.a(s_87), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1160(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1161(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1162(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1023(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1024(.a(gate387inter0), .b(s_68), .O(gate387inter1));
  and2  gate1025(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1026(.a(s_68), .O(gate387inter3));
  inv1  gate1027(.a(s_69), .O(gate387inter4));
  nand2 gate1028(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1029(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1030(.a(G1), .O(gate387inter7));
  inv1  gate1031(.a(G1036), .O(gate387inter8));
  nand2 gate1032(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1033(.a(s_69), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1034(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1035(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1036(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1331(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1332(.a(gate392inter0), .b(s_112), .O(gate392inter1));
  and2  gate1333(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1334(.a(s_112), .O(gate392inter3));
  inv1  gate1335(.a(s_113), .O(gate392inter4));
  nand2 gate1336(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1337(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1338(.a(G6), .O(gate392inter7));
  inv1  gate1339(.a(G1051), .O(gate392inter8));
  nand2 gate1340(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1341(.a(s_113), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1342(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1343(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1344(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1051(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1052(.a(gate397inter0), .b(s_72), .O(gate397inter1));
  and2  gate1053(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1054(.a(s_72), .O(gate397inter3));
  inv1  gate1055(.a(s_73), .O(gate397inter4));
  nand2 gate1056(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1057(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1058(.a(G11), .O(gate397inter7));
  inv1  gate1059(.a(G1066), .O(gate397inter8));
  nand2 gate1060(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1061(.a(s_73), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1062(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1063(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1064(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate743(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate744(.a(gate400inter0), .b(s_28), .O(gate400inter1));
  and2  gate745(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate746(.a(s_28), .O(gate400inter3));
  inv1  gate747(.a(s_29), .O(gate400inter4));
  nand2 gate748(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate749(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate750(.a(G14), .O(gate400inter7));
  inv1  gate751(.a(G1075), .O(gate400inter8));
  nand2 gate752(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate753(.a(s_29), .b(gate400inter3), .O(gate400inter10));
  nor2  gate754(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate755(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate756(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1261(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1262(.a(gate404inter0), .b(s_102), .O(gate404inter1));
  and2  gate1263(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1264(.a(s_102), .O(gate404inter3));
  inv1  gate1265(.a(s_103), .O(gate404inter4));
  nand2 gate1266(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1267(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1268(.a(G18), .O(gate404inter7));
  inv1  gate1269(.a(G1087), .O(gate404inter8));
  nand2 gate1270(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1271(.a(s_103), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1272(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1273(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1274(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate869(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate870(.a(gate405inter0), .b(s_46), .O(gate405inter1));
  and2  gate871(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate872(.a(s_46), .O(gate405inter3));
  inv1  gate873(.a(s_47), .O(gate405inter4));
  nand2 gate874(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate875(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate876(.a(G19), .O(gate405inter7));
  inv1  gate877(.a(G1090), .O(gate405inter8));
  nand2 gate878(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate879(.a(s_47), .b(gate405inter3), .O(gate405inter10));
  nor2  gate880(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate881(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate882(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate953(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate954(.a(gate417inter0), .b(s_58), .O(gate417inter1));
  and2  gate955(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate956(.a(s_58), .O(gate417inter3));
  inv1  gate957(.a(s_59), .O(gate417inter4));
  nand2 gate958(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate959(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate960(.a(G31), .O(gate417inter7));
  inv1  gate961(.a(G1126), .O(gate417inter8));
  nand2 gate962(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate963(.a(s_59), .b(gate417inter3), .O(gate417inter10));
  nor2  gate964(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate965(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate966(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1093(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1094(.a(gate420inter0), .b(s_78), .O(gate420inter1));
  and2  gate1095(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1096(.a(s_78), .O(gate420inter3));
  inv1  gate1097(.a(s_79), .O(gate420inter4));
  nand2 gate1098(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1099(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1100(.a(G1036), .O(gate420inter7));
  inv1  gate1101(.a(G1132), .O(gate420inter8));
  nand2 gate1102(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1103(.a(s_79), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1104(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1105(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1106(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate561(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate562(.a(gate422inter0), .b(s_2), .O(gate422inter1));
  and2  gate563(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate564(.a(s_2), .O(gate422inter3));
  inv1  gate565(.a(s_3), .O(gate422inter4));
  nand2 gate566(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate567(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate568(.a(G1039), .O(gate422inter7));
  inv1  gate569(.a(G1135), .O(gate422inter8));
  nand2 gate570(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate571(.a(s_3), .b(gate422inter3), .O(gate422inter10));
  nor2  gate572(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate573(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate574(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1429(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1430(.a(gate423inter0), .b(s_126), .O(gate423inter1));
  and2  gate1431(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1432(.a(s_126), .O(gate423inter3));
  inv1  gate1433(.a(s_127), .O(gate423inter4));
  nand2 gate1434(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1435(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1436(.a(G3), .O(gate423inter7));
  inv1  gate1437(.a(G1138), .O(gate423inter8));
  nand2 gate1438(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1439(.a(s_127), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1440(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1441(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1442(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1457(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1458(.a(gate425inter0), .b(s_130), .O(gate425inter1));
  and2  gate1459(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1460(.a(s_130), .O(gate425inter3));
  inv1  gate1461(.a(s_131), .O(gate425inter4));
  nand2 gate1462(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1463(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1464(.a(G4), .O(gate425inter7));
  inv1  gate1465(.a(G1141), .O(gate425inter8));
  nand2 gate1466(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1467(.a(s_131), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1468(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1469(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1470(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate645(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate646(.a(gate441inter0), .b(s_14), .O(gate441inter1));
  and2  gate647(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate648(.a(s_14), .O(gate441inter3));
  inv1  gate649(.a(s_15), .O(gate441inter4));
  nand2 gate650(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate651(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate652(.a(G12), .O(gate441inter7));
  inv1  gate653(.a(G1165), .O(gate441inter8));
  nand2 gate654(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate655(.a(s_15), .b(gate441inter3), .O(gate441inter10));
  nor2  gate656(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate657(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate658(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1401(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1402(.a(gate445inter0), .b(s_122), .O(gate445inter1));
  and2  gate1403(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1404(.a(s_122), .O(gate445inter3));
  inv1  gate1405(.a(s_123), .O(gate445inter4));
  nand2 gate1406(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1407(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1408(.a(G14), .O(gate445inter7));
  inv1  gate1409(.a(G1171), .O(gate445inter8));
  nand2 gate1410(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1411(.a(s_123), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1412(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1413(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1414(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1387(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1388(.a(gate446inter0), .b(s_120), .O(gate446inter1));
  and2  gate1389(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1390(.a(s_120), .O(gate446inter3));
  inv1  gate1391(.a(s_121), .O(gate446inter4));
  nand2 gate1392(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1393(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1394(.a(G1075), .O(gate446inter7));
  inv1  gate1395(.a(G1171), .O(gate446inter8));
  nand2 gate1396(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1397(.a(s_121), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1398(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1399(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1400(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1247(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1248(.a(gate456inter0), .b(s_100), .O(gate456inter1));
  and2  gate1249(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1250(.a(s_100), .O(gate456inter3));
  inv1  gate1251(.a(s_101), .O(gate456inter4));
  nand2 gate1252(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1253(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1254(.a(G1090), .O(gate456inter7));
  inv1  gate1255(.a(G1186), .O(gate456inter8));
  nand2 gate1256(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1257(.a(s_101), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1258(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1259(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1260(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate715(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate716(.a(gate457inter0), .b(s_24), .O(gate457inter1));
  and2  gate717(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate718(.a(s_24), .O(gate457inter3));
  inv1  gate719(.a(s_25), .O(gate457inter4));
  nand2 gate720(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate721(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate722(.a(G20), .O(gate457inter7));
  inv1  gate723(.a(G1189), .O(gate457inter8));
  nand2 gate724(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate725(.a(s_25), .b(gate457inter3), .O(gate457inter10));
  nor2  gate726(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate727(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate728(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1317(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1318(.a(gate489inter0), .b(s_110), .O(gate489inter1));
  and2  gate1319(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1320(.a(s_110), .O(gate489inter3));
  inv1  gate1321(.a(s_111), .O(gate489inter4));
  nand2 gate1322(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1323(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1324(.a(G1240), .O(gate489inter7));
  inv1  gate1325(.a(G1241), .O(gate489inter8));
  nand2 gate1326(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1327(.a(s_111), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1328(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1329(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1330(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1177(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1178(.a(gate492inter0), .b(s_90), .O(gate492inter1));
  and2  gate1179(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1180(.a(s_90), .O(gate492inter3));
  inv1  gate1181(.a(s_91), .O(gate492inter4));
  nand2 gate1182(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1183(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1184(.a(G1246), .O(gate492inter7));
  inv1  gate1185(.a(G1247), .O(gate492inter8));
  nand2 gate1186(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1187(.a(s_91), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1188(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1189(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1190(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1527(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1528(.a(gate496inter0), .b(s_140), .O(gate496inter1));
  and2  gate1529(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1530(.a(s_140), .O(gate496inter3));
  inv1  gate1531(.a(s_141), .O(gate496inter4));
  nand2 gate1532(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1533(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1534(.a(G1254), .O(gate496inter7));
  inv1  gate1535(.a(G1255), .O(gate496inter8));
  nand2 gate1536(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1537(.a(s_141), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1538(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1539(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1540(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1275(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1276(.a(gate497inter0), .b(s_104), .O(gate497inter1));
  and2  gate1277(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1278(.a(s_104), .O(gate497inter3));
  inv1  gate1279(.a(s_105), .O(gate497inter4));
  nand2 gate1280(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1281(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1282(.a(G1256), .O(gate497inter7));
  inv1  gate1283(.a(G1257), .O(gate497inter8));
  nand2 gate1284(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1285(.a(s_105), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1286(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1287(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1288(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1443(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1444(.a(gate498inter0), .b(s_128), .O(gate498inter1));
  and2  gate1445(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1446(.a(s_128), .O(gate498inter3));
  inv1  gate1447(.a(s_129), .O(gate498inter4));
  nand2 gate1448(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1449(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1450(.a(G1258), .O(gate498inter7));
  inv1  gate1451(.a(G1259), .O(gate498inter8));
  nand2 gate1452(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1453(.a(s_129), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1454(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1455(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1456(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate925(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate926(.a(gate501inter0), .b(s_54), .O(gate501inter1));
  and2  gate927(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate928(.a(s_54), .O(gate501inter3));
  inv1  gate929(.a(s_55), .O(gate501inter4));
  nand2 gate930(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate931(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate932(.a(G1264), .O(gate501inter7));
  inv1  gate933(.a(G1265), .O(gate501inter8));
  nand2 gate934(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate935(.a(s_55), .b(gate501inter3), .O(gate501inter10));
  nor2  gate936(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate937(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate938(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1513(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1514(.a(gate508inter0), .b(s_138), .O(gate508inter1));
  and2  gate1515(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1516(.a(s_138), .O(gate508inter3));
  inv1  gate1517(.a(s_139), .O(gate508inter4));
  nand2 gate1518(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1519(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1520(.a(G1278), .O(gate508inter7));
  inv1  gate1521(.a(G1279), .O(gate508inter8));
  nand2 gate1522(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1523(.a(s_139), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1524(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1525(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1526(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule