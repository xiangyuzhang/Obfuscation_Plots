module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );

  xor2  gate749(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate750(.a(gate21inter0), .b(s_84), .O(gate21inter1));
  and2  gate751(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate752(.a(s_84), .O(gate21inter3));
  inv1  gate753(.a(s_85), .O(gate21inter4));
  nand2 gate754(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate755(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate756(.a(N14), .O(gate21inter7));
  inv1  gate757(.a(N119), .O(gate21inter8));
  nand2 gate758(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate759(.a(s_85), .b(gate21inter3), .O(gate21inter10));
  nor2  gate760(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate761(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate762(.a(gate21inter12), .b(gate21inter1), .O(N158));

  xor2  gate483(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate484(.a(gate22inter0), .b(s_46), .O(gate22inter1));
  and2  gate485(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate486(.a(s_46), .O(gate22inter3));
  inv1  gate487(.a(s_47), .O(gate22inter4));
  nand2 gate488(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate489(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate490(.a(N122), .O(gate22inter7));
  inv1  gate491(.a(N17), .O(gate22inter8));
  nand2 gate492(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate493(.a(s_47), .b(gate22inter3), .O(gate22inter10));
  nor2  gate494(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate495(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate496(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate217(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate218(.a(gate24inter0), .b(s_8), .O(gate24inter1));
  and2  gate219(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate220(.a(s_8), .O(gate24inter3));
  inv1  gate221(.a(s_9), .O(gate24inter4));
  nand2 gate222(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate223(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate224(.a(N130), .O(gate24inter7));
  inv1  gate225(.a(N43), .O(gate24inter8));
  nand2 gate226(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate227(.a(s_9), .b(gate24inter3), .O(gate24inter10));
  nor2  gate228(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate229(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate230(.a(gate24inter12), .b(gate24inter1), .O(N165));

  xor2  gate203(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate204(.a(gate25inter0), .b(s_6), .O(gate25inter1));
  and2  gate205(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate206(.a(s_6), .O(gate25inter3));
  inv1  gate207(.a(s_7), .O(gate25inter4));
  nand2 gate208(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate209(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate210(.a(N134), .O(gate25inter7));
  inv1  gate211(.a(N56), .O(gate25inter8));
  nand2 gate212(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate213(.a(s_7), .b(gate25inter3), .O(gate25inter10));
  nor2  gate214(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate215(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate216(.a(gate25inter12), .b(gate25inter1), .O(N168));

  xor2  gate665(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate666(.a(gate26inter0), .b(s_72), .O(gate26inter1));
  and2  gate667(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate668(.a(s_72), .O(gate26inter3));
  inv1  gate669(.a(s_73), .O(gate26inter4));
  nand2 gate670(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate671(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate672(.a(N138), .O(gate26inter7));
  inv1  gate673(.a(N69), .O(gate26inter8));
  nand2 gate674(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate675(.a(s_73), .b(gate26inter3), .O(gate26inter10));
  nor2  gate676(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate677(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate678(.a(gate26inter12), .b(gate26inter1), .O(N171));
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate525(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate526(.a(gate30inter0), .b(s_52), .O(gate30inter1));
  and2  gate527(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate528(.a(s_52), .O(gate30inter3));
  inv1  gate529(.a(s_53), .O(gate30inter4));
  nand2 gate530(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate531(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate532(.a(N21), .O(gate30inter7));
  inv1  gate533(.a(N123), .O(gate30inter8));
  nand2 gate534(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate535(.a(s_53), .b(gate30inter3), .O(gate30inter10));
  nor2  gate536(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate537(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate538(.a(gate30inter12), .b(gate30inter1), .O(N183));
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate595(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate596(.a(gate32inter0), .b(s_62), .O(gate32inter1));
  and2  gate597(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate598(.a(s_62), .O(gate32inter3));
  inv1  gate599(.a(s_63), .O(gate32inter4));
  nand2 gate600(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate601(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate602(.a(N34), .O(gate32inter7));
  inv1  gate603(.a(N127), .O(gate32inter8));
  nand2 gate604(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate605(.a(s_63), .b(gate32inter3), .O(gate32inter10));
  nor2  gate606(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate607(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate608(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate427(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate428(.a(gate36inter0), .b(s_38), .O(gate36inter1));
  and2  gate429(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate430(.a(s_38), .O(gate36inter3));
  inv1  gate431(.a(s_39), .O(gate36inter4));
  nand2 gate432(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate433(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate434(.a(N60), .O(gate36inter7));
  inv1  gate435(.a(N135), .O(gate36inter8));
  nand2 gate436(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate437(.a(s_39), .b(gate36inter3), .O(gate36inter10));
  nor2  gate438(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate439(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate440(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate175(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate176(.a(gate38inter0), .b(s_2), .O(gate38inter1));
  and2  gate177(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate178(.a(s_2), .O(gate38inter3));
  inv1  gate179(.a(s_3), .O(gate38inter4));
  nand2 gate180(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate181(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate182(.a(N73), .O(gate38inter7));
  inv1  gate183(.a(N139), .O(gate38inter8));
  nand2 gate184(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate185(.a(s_3), .b(gate38inter3), .O(gate38inter10));
  nor2  gate186(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate187(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate188(.a(gate38inter12), .b(gate38inter1), .O(N191));

  xor2  gate679(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate680(.a(gate39inter0), .b(s_74), .O(gate39inter1));
  and2  gate681(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate682(.a(s_74), .O(gate39inter3));
  inv1  gate683(.a(s_75), .O(gate39inter4));
  nand2 gate684(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate685(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate686(.a(N79), .O(gate39inter7));
  inv1  gate687(.a(N139), .O(gate39inter8));
  nand2 gate688(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate689(.a(s_75), .b(gate39inter3), .O(gate39inter10));
  nor2  gate690(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate691(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate692(.a(gate39inter12), .b(gate39inter1), .O(N192));

  xor2  gate399(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate400(.a(gate40inter0), .b(s_34), .O(gate40inter1));
  and2  gate401(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate402(.a(s_34), .O(gate40inter3));
  inv1  gate403(.a(s_35), .O(gate40inter4));
  nand2 gate404(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate405(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate406(.a(N86), .O(gate40inter7));
  inv1  gate407(.a(N143), .O(gate40inter8));
  nand2 gate408(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate409(.a(s_35), .b(gate40inter3), .O(gate40inter10));
  nor2  gate410(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate411(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate412(.a(gate40inter12), .b(gate40inter1), .O(N193));

  xor2  gate735(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate736(.a(gate41inter0), .b(s_82), .O(gate41inter1));
  and2  gate737(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate738(.a(s_82), .O(gate41inter3));
  inv1  gate739(.a(s_83), .O(gate41inter4));
  nand2 gate740(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate741(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate742(.a(N92), .O(gate41inter7));
  inv1  gate743(.a(N143), .O(gate41inter8));
  nand2 gate744(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate745(.a(s_83), .b(gate41inter3), .O(gate41inter10));
  nor2  gate746(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate747(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate748(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate329(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate330(.a(gate43inter0), .b(s_24), .O(gate43inter1));
  and2  gate331(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate332(.a(s_24), .O(gate43inter3));
  inv1  gate333(.a(s_25), .O(gate43inter4));
  nand2 gate334(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate335(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate336(.a(N105), .O(gate43inter7));
  inv1  gate337(.a(N147), .O(gate43inter8));
  nand2 gate338(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate339(.a(s_25), .b(gate43inter3), .O(gate43inter10));
  nor2  gate340(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate341(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate342(.a(gate43inter12), .b(gate43inter1), .O(N196));

  xor2  gate567(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate568(.a(gate44inter0), .b(s_58), .O(gate44inter1));
  and2  gate569(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate570(.a(s_58), .O(gate44inter3));
  inv1  gate571(.a(s_59), .O(gate44inter4));
  nand2 gate572(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate573(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate574(.a(N112), .O(gate44inter7));
  inv1  gate575(.a(N151), .O(gate44inter8));
  nand2 gate576(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate577(.a(s_59), .b(gate44inter3), .O(gate44inter10));
  nor2  gate578(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate579(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate580(.a(gate44inter12), .b(gate44inter1), .O(N197));

  xor2  gate609(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate610(.a(gate45inter0), .b(s_64), .O(gate45inter1));
  and2  gate611(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate612(.a(s_64), .O(gate45inter3));
  inv1  gate613(.a(s_65), .O(gate45inter4));
  nand2 gate614(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate615(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate616(.a(N115), .O(gate45inter7));
  inv1  gate617(.a(N151), .O(gate45inter8));
  nand2 gate618(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate619(.a(s_65), .b(gate45inter3), .O(gate45inter10));
  nor2  gate620(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate621(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate622(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate245(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate246(.a(gate52inter0), .b(s_12), .O(gate52inter1));
  and2  gate247(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate248(.a(s_12), .O(gate52inter3));
  inv1  gate249(.a(s_13), .O(gate52inter4));
  nand2 gate250(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate251(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate252(.a(N203), .O(gate52inter7));
  inv1  gate253(.a(N162), .O(gate52inter8));
  nand2 gate254(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate255(.a(s_13), .b(gate52inter3), .O(gate52inter10));
  nor2  gate256(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate257(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate258(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );

  xor2  gate763(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate764(.a(gate55inter0), .b(s_86), .O(gate55inter1));
  and2  gate765(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate766(.a(s_86), .O(gate55inter3));
  inv1  gate767(.a(s_87), .O(gate55inter4));
  nand2 gate768(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate769(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate770(.a(N203), .O(gate55inter7));
  inv1  gate771(.a(N171), .O(gate55inter8));
  nand2 gate772(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate773(.a(s_87), .b(gate55inter3), .O(gate55inter10));
  nor2  gate774(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate775(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate776(.a(gate55inter12), .b(gate55inter1), .O(N239));

  xor2  gate231(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate232(.a(gate56inter0), .b(s_10), .O(gate56inter1));
  and2  gate233(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate234(.a(s_10), .O(gate56inter3));
  inv1  gate235(.a(s_11), .O(gate56inter4));
  nand2 gate236(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate237(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate238(.a(N1), .O(gate56inter7));
  inv1  gate239(.a(N213), .O(gate56inter8));
  nand2 gate240(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate241(.a(s_11), .b(gate56inter3), .O(gate56inter10));
  nor2  gate242(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate243(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate244(.a(gate56inter12), .b(gate56inter1), .O(N242));

  xor2  gate511(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate512(.a(gate57inter0), .b(s_50), .O(gate57inter1));
  and2  gate513(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate514(.a(s_50), .O(gate57inter3));
  inv1  gate515(.a(s_51), .O(gate57inter4));
  nand2 gate516(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate517(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate518(.a(N203), .O(gate57inter7));
  inv1  gate519(.a(N174), .O(gate57inter8));
  nand2 gate520(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate521(.a(s_51), .b(gate57inter3), .O(gate57inter10));
  nor2  gate522(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate523(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate524(.a(gate57inter12), .b(gate57inter1), .O(N243));

  xor2  gate791(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate792(.a(gate58inter0), .b(s_90), .O(gate58inter1));
  and2  gate793(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate794(.a(s_90), .O(gate58inter3));
  inv1  gate795(.a(s_91), .O(gate58inter4));
  nand2 gate796(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate797(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate798(.a(N213), .O(gate58inter7));
  inv1  gate799(.a(N11), .O(gate58inter8));
  nand2 gate800(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate801(.a(s_91), .b(gate58inter3), .O(gate58inter10));
  nor2  gate802(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate803(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate804(.a(gate58inter12), .b(gate58inter1), .O(N246));

  xor2  gate301(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate302(.a(gate59inter0), .b(s_20), .O(gate59inter1));
  and2  gate303(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate304(.a(s_20), .O(gate59inter3));
  inv1  gate305(.a(s_21), .O(gate59inter4));
  nand2 gate306(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate307(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate308(.a(N203), .O(gate59inter7));
  inv1  gate309(.a(N177), .O(gate59inter8));
  nand2 gate310(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate311(.a(s_21), .b(gate59inter3), .O(gate59inter10));
  nor2  gate312(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate313(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate314(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );

  xor2  gate357(.a(N180), .b(N203), .O(gate61inter0));
  nand2 gate358(.a(gate61inter0), .b(s_28), .O(gate61inter1));
  and2  gate359(.a(N180), .b(N203), .O(gate61inter2));
  inv1  gate360(.a(s_28), .O(gate61inter3));
  inv1  gate361(.a(s_29), .O(gate61inter4));
  nand2 gate362(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate363(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate364(.a(N203), .O(gate61inter7));
  inv1  gate365(.a(N180), .O(gate61inter8));
  nand2 gate366(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate367(.a(s_29), .b(gate61inter3), .O(gate61inter10));
  nor2  gate368(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate369(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate370(.a(gate61inter12), .b(gate61inter1), .O(N251));
nand2 gate62( .a(N213), .b(N37), .O(N254) );

  xor2  gate371(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate372(.a(gate63inter0), .b(s_30), .O(gate63inter1));
  and2  gate373(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate374(.a(s_30), .O(gate63inter3));
  inv1  gate375(.a(s_31), .O(gate63inter4));
  nand2 gate376(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate377(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate378(.a(N213), .O(gate63inter7));
  inv1  gate379(.a(N50), .O(gate63inter8));
  nand2 gate380(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate381(.a(s_31), .b(gate63inter3), .O(gate63inter10));
  nor2  gate382(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate383(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate384(.a(gate63inter12), .b(gate63inter1), .O(N255));
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate161(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate162(.a(gate65inter0), .b(s_0), .O(gate65inter1));
  and2  gate163(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate164(.a(s_0), .O(gate65inter3));
  inv1  gate165(.a(s_1), .O(gate65inter4));
  nand2 gate166(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate167(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate168(.a(N213), .O(gate65inter7));
  inv1  gate169(.a(N76), .O(gate65inter8));
  nand2 gate170(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate171(.a(s_1), .b(gate65inter3), .O(gate65inter10));
  nor2  gate172(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate173(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate174(.a(gate65inter12), .b(gate65inter1), .O(N257));

  xor2  gate385(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate386(.a(gate66inter0), .b(s_32), .O(gate66inter1));
  and2  gate387(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate388(.a(s_32), .O(gate66inter3));
  inv1  gate389(.a(s_33), .O(gate66inter4));
  nand2 gate390(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate391(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate392(.a(N213), .O(gate66inter7));
  inv1  gate393(.a(N89), .O(gate66inter8));
  nand2 gate394(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate395(.a(s_33), .b(gate66inter3), .O(gate66inter10));
  nor2  gate396(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate397(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate398(.a(gate66inter12), .b(gate66inter1), .O(N258));

  xor2  gate903(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate904(.a(gate67inter0), .b(s_106), .O(gate67inter1));
  and2  gate905(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate906(.a(s_106), .O(gate67inter3));
  inv1  gate907(.a(s_107), .O(gate67inter4));
  nand2 gate908(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate909(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate910(.a(N213), .O(gate67inter7));
  inv1  gate911(.a(N102), .O(gate67inter8));
  nand2 gate912(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate913(.a(s_107), .b(gate67inter3), .O(gate67inter10));
  nor2  gate914(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate915(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate916(.a(gate67inter12), .b(gate67inter1), .O(N259));

  xor2  gate553(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate554(.a(gate68inter0), .b(s_56), .O(gate68inter1));
  and2  gate555(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate556(.a(s_56), .O(gate68inter3));
  inv1  gate557(.a(s_57), .O(gate68inter4));
  nand2 gate558(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate559(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate560(.a(N224), .O(gate68inter7));
  inv1  gate561(.a(N157), .O(gate68inter8));
  nand2 gate562(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate563(.a(s_57), .b(gate68inter3), .O(gate68inter10));
  nor2  gate564(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate565(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate566(.a(gate68inter12), .b(gate68inter1), .O(N260));

  xor2  gate539(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate540(.a(gate69inter0), .b(s_54), .O(gate69inter1));
  and2  gate541(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate542(.a(s_54), .O(gate69inter3));
  inv1  gate543(.a(s_55), .O(gate69inter4));
  nand2 gate544(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate545(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate546(.a(N224), .O(gate69inter7));
  inv1  gate547(.a(N158), .O(gate69inter8));
  nand2 gate548(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate549(.a(s_55), .b(gate69inter3), .O(gate69inter10));
  nor2  gate550(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate551(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate552(.a(gate69inter12), .b(gate69inter1), .O(N263));

  xor2  gate875(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate876(.a(gate70inter0), .b(s_102), .O(gate70inter1));
  and2  gate877(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate878(.a(s_102), .O(gate70inter3));
  inv1  gate879(.a(s_103), .O(gate70inter4));
  nand2 gate880(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate881(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate882(.a(N227), .O(gate70inter7));
  inv1  gate883(.a(N183), .O(gate70inter8));
  nand2 gate884(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate885(.a(s_103), .b(gate70inter3), .O(gate70inter10));
  nor2  gate886(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate887(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate888(.a(gate70inter12), .b(gate70inter1), .O(N264));

  xor2  gate805(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate806(.a(gate71inter0), .b(s_92), .O(gate71inter1));
  and2  gate807(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate808(.a(s_92), .O(gate71inter3));
  inv1  gate809(.a(s_93), .O(gate71inter4));
  nand2 gate810(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate811(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate812(.a(N230), .O(gate71inter7));
  inv1  gate813(.a(N185), .O(gate71inter8));
  nand2 gate814(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate815(.a(s_93), .b(gate71inter3), .O(gate71inter10));
  nor2  gate816(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate817(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate818(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );

  xor2  gate889(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate890(.a(gate74inter0), .b(s_104), .O(gate74inter1));
  and2  gate891(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate892(.a(s_104), .O(gate74inter3));
  inv1  gate893(.a(s_105), .O(gate74inter4));
  nand2 gate894(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate895(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate896(.a(N239), .O(gate74inter7));
  inv1  gate897(.a(N191), .O(gate74inter8));
  nand2 gate898(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate899(.a(s_105), .b(gate74inter3), .O(gate74inter10));
  nor2  gate900(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate901(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate902(.a(gate74inter12), .b(gate74inter1), .O(N276));
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate847(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate848(.a(gate78inter0), .b(s_98), .O(gate78inter1));
  and2  gate849(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate850(.a(s_98), .O(gate78inter3));
  inv1  gate851(.a(s_99), .O(gate78inter4));
  nand2 gate852(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate853(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate854(.a(N227), .O(gate78inter7));
  inv1  gate855(.a(N184), .O(gate78inter8));
  nand2 gate856(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate857(.a(s_99), .b(gate78inter3), .O(gate78inter10));
  nor2  gate858(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate859(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate860(.a(gate78inter12), .b(gate78inter1), .O(N288));

  xor2  gate441(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate442(.a(gate79inter0), .b(s_40), .O(gate79inter1));
  and2  gate443(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate444(.a(s_40), .O(gate79inter3));
  inv1  gate445(.a(s_41), .O(gate79inter4));
  nand2 gate446(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate447(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate448(.a(N230), .O(gate79inter7));
  inv1  gate449(.a(N186), .O(gate79inter8));
  nand2 gate450(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate451(.a(s_41), .b(gate79inter3), .O(gate79inter10));
  nor2  gate452(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate453(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate454(.a(gate79inter12), .b(gate79inter1), .O(N289));

  xor2  gate455(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate456(.a(gate80inter0), .b(s_42), .O(gate80inter1));
  and2  gate457(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate458(.a(s_42), .O(gate80inter3));
  inv1  gate459(.a(s_43), .O(gate80inter4));
  nand2 gate460(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate461(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate462(.a(N233), .O(gate80inter7));
  inv1  gate463(.a(N188), .O(gate80inter8));
  nand2 gate464(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate465(.a(s_43), .b(gate80inter3), .O(gate80inter10));
  nor2  gate466(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate467(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate468(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );

  xor2  gate651(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate652(.a(gate85inter0), .b(s_70), .O(gate85inter1));
  and2  gate653(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate654(.a(s_70), .O(gate85inter3));
  inv1  gate655(.a(s_71), .O(gate85inter4));
  nand2 gate656(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate657(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate658(.a(N251), .O(gate85inter7));
  inv1  gate659(.a(N198), .O(gate85inter8));
  nand2 gate660(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate661(.a(s_71), .b(gate85inter3), .O(gate85inter10));
  nor2  gate662(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate663(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate664(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );

  xor2  gate819(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate820(.a(gate101inter0), .b(s_94), .O(gate101inter1));
  and2  gate821(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate822(.a(s_94), .O(gate101inter3));
  inv1  gate823(.a(s_95), .O(gate101inter4));
  nand2 gate824(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate825(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate826(.a(N309), .O(gate101inter7));
  inv1  gate827(.a(N267), .O(gate101inter8));
  nand2 gate828(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate829(.a(s_95), .b(gate101inter3), .O(gate101inter10));
  nor2  gate830(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate831(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate832(.a(gate101inter12), .b(gate101inter1), .O(N332));

  xor2  gate707(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate708(.a(gate102inter0), .b(s_78), .O(gate102inter1));
  and2  gate709(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate710(.a(s_78), .O(gate102inter3));
  inv1  gate711(.a(s_79), .O(gate102inter4));
  nand2 gate712(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate713(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate714(.a(N309), .O(gate102inter7));
  inv1  gate715(.a(N270), .O(gate102inter8));
  nand2 gate716(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate717(.a(s_79), .b(gate102inter3), .O(gate102inter10));
  nor2  gate718(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate719(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate720(.a(gate102inter12), .b(gate102inter1), .O(N333));

  xor2  gate833(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate834(.a(gate103inter0), .b(s_96), .O(gate103inter1));
  and2  gate835(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate836(.a(s_96), .O(gate103inter3));
  inv1  gate837(.a(s_97), .O(gate103inter4));
  nand2 gate838(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate839(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate840(.a(N8), .O(gate103inter7));
  inv1  gate841(.a(N319), .O(gate103inter8));
  nand2 gate842(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate843(.a(s_97), .b(gate103inter3), .O(gate103inter10));
  nor2  gate844(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate845(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate846(.a(gate103inter12), .b(gate103inter1), .O(N334));

  xor2  gate273(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate274(.a(gate104inter0), .b(s_16), .O(gate104inter1));
  and2  gate275(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate276(.a(s_16), .O(gate104inter3));
  inv1  gate277(.a(s_17), .O(gate104inter4));
  nand2 gate278(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate279(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate280(.a(N309), .O(gate104inter7));
  inv1  gate281(.a(N273), .O(gate104inter8));
  nand2 gate282(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate283(.a(s_17), .b(gate104inter3), .O(gate104inter10));
  nor2  gate284(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate285(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate286(.a(gate104inter12), .b(gate104inter1), .O(N335));

  xor2  gate917(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate918(.a(gate105inter0), .b(s_108), .O(gate105inter1));
  and2  gate919(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate920(.a(s_108), .O(gate105inter3));
  inv1  gate921(.a(s_109), .O(gate105inter4));
  nand2 gate922(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate923(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate924(.a(N319), .O(gate105inter7));
  inv1  gate925(.a(N21), .O(gate105inter8));
  nand2 gate926(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate927(.a(s_109), .b(gate105inter3), .O(gate105inter10));
  nor2  gate928(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate929(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate930(.a(gate105inter12), .b(gate105inter1), .O(N336));

  xor2  gate581(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate582(.a(gate106inter0), .b(s_60), .O(gate106inter1));
  and2  gate583(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate584(.a(s_60), .O(gate106inter3));
  inv1  gate585(.a(s_61), .O(gate106inter4));
  nand2 gate586(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate587(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate588(.a(N309), .O(gate106inter7));
  inv1  gate589(.a(N276), .O(gate106inter8));
  nand2 gate590(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate591(.a(s_61), .b(gate106inter3), .O(gate106inter10));
  nor2  gate592(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate593(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate594(.a(gate106inter12), .b(gate106inter1), .O(N337));

  xor2  gate287(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate288(.a(gate107inter0), .b(s_18), .O(gate107inter1));
  and2  gate289(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate290(.a(s_18), .O(gate107inter3));
  inv1  gate291(.a(s_19), .O(gate107inter4));
  nand2 gate292(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate293(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate294(.a(N319), .O(gate107inter7));
  inv1  gate295(.a(N34), .O(gate107inter8));
  nand2 gate296(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate297(.a(s_19), .b(gate107inter3), .O(gate107inter10));
  nor2  gate298(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate299(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate300(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );

  xor2  gate721(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate722(.a(gate109inter0), .b(s_80), .O(gate109inter1));
  and2  gate723(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate724(.a(s_80), .O(gate109inter3));
  inv1  gate725(.a(s_81), .O(gate109inter4));
  nand2 gate726(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate727(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate728(.a(N319), .O(gate109inter7));
  inv1  gate729(.a(N47), .O(gate109inter8));
  nand2 gate730(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate731(.a(s_81), .b(gate109inter3), .O(gate109inter10));
  nor2  gate732(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate733(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate734(.a(gate109inter12), .b(gate109inter1), .O(N340));

  xor2  gate189(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate190(.a(gate110inter0), .b(s_4), .O(gate110inter1));
  and2  gate191(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate192(.a(s_4), .O(gate110inter3));
  inv1  gate193(.a(s_5), .O(gate110inter4));
  nand2 gate194(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate195(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate196(.a(N309), .O(gate110inter7));
  inv1  gate197(.a(N282), .O(gate110inter8));
  nand2 gate198(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate199(.a(s_5), .b(gate110inter3), .O(gate110inter10));
  nor2  gate200(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate201(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate202(.a(gate110inter12), .b(gate110inter1), .O(N341));

  xor2  gate777(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate778(.a(gate111inter0), .b(s_88), .O(gate111inter1));
  and2  gate779(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate780(.a(s_88), .O(gate111inter3));
  inv1  gate781(.a(s_89), .O(gate111inter4));
  nand2 gate782(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate783(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate784(.a(N319), .O(gate111inter7));
  inv1  gate785(.a(N60), .O(gate111inter8));
  nand2 gate786(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate787(.a(s_89), .b(gate111inter3), .O(gate111inter10));
  nor2  gate788(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate789(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate790(.a(gate111inter12), .b(gate111inter1), .O(N342));

  xor2  gate637(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate638(.a(gate112inter0), .b(s_68), .O(gate112inter1));
  and2  gate639(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate640(.a(s_68), .O(gate112inter3));
  inv1  gate641(.a(s_69), .O(gate112inter4));
  nand2 gate642(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate643(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate644(.a(N309), .O(gate112inter7));
  inv1  gate645(.a(N285), .O(gate112inter8));
  nand2 gate646(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate647(.a(s_69), .b(gate112inter3), .O(gate112inter10));
  nor2  gate648(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate649(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate650(.a(gate112inter12), .b(gate112inter1), .O(N343));

  xor2  gate497(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate498(.a(gate113inter0), .b(s_48), .O(gate113inter1));
  and2  gate499(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate500(.a(s_48), .O(gate113inter3));
  inv1  gate501(.a(s_49), .O(gate113inter4));
  nand2 gate502(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate503(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate504(.a(N319), .O(gate113inter7));
  inv1  gate505(.a(N73), .O(gate113inter8));
  nand2 gate506(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate507(.a(s_49), .b(gate113inter3), .O(gate113inter10));
  nor2  gate508(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate509(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate510(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate693(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate694(.a(gate115inter0), .b(s_76), .O(gate115inter1));
  and2  gate695(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate696(.a(s_76), .O(gate115inter3));
  inv1  gate697(.a(s_77), .O(gate115inter4));
  nand2 gate698(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate699(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate700(.a(N319), .O(gate115inter7));
  inv1  gate701(.a(N99), .O(gate115inter8));
  nand2 gate702(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate703(.a(s_77), .b(gate115inter3), .O(gate115inter10));
  nor2  gate704(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate705(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate706(.a(gate115inter12), .b(gate115inter1), .O(N346));

  xor2  gate623(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate624(.a(gate116inter0), .b(s_66), .O(gate116inter1));
  and2  gate625(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate626(.a(s_66), .O(gate116inter3));
  inv1  gate627(.a(s_67), .O(gate116inter4));
  nand2 gate628(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate629(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate630(.a(N319), .O(gate116inter7));
  inv1  gate631(.a(N112), .O(gate116inter8));
  nand2 gate632(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate633(.a(s_67), .b(gate116inter3), .O(gate116inter10));
  nor2  gate634(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate635(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate636(.a(gate116inter12), .b(gate116inter1), .O(N347));
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate931(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate932(.a(gate118inter0), .b(s_110), .O(gate118inter1));
  and2  gate933(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate934(.a(s_110), .O(gate118inter3));
  inv1  gate935(.a(s_111), .O(gate118inter4));
  nand2 gate936(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate937(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate938(.a(N331), .O(gate118inter7));
  inv1  gate939(.a(N301), .O(gate118inter8));
  nand2 gate940(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate941(.a(s_111), .b(gate118inter3), .O(gate118inter10));
  nor2  gate942(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate943(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate944(.a(gate118inter12), .b(gate118inter1), .O(N349));
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate259(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate260(.a(gate120inter0), .b(s_14), .O(gate120inter1));
  and2  gate261(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate262(.a(s_14), .O(gate120inter3));
  inv1  gate263(.a(s_15), .O(gate120inter4));
  nand2 gate264(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate265(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate266(.a(N333), .O(gate120inter7));
  inv1  gate267(.a(N303), .O(gate120inter8));
  nand2 gate268(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate269(.a(s_15), .b(gate120inter3), .O(gate120inter10));
  nor2  gate270(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate271(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate272(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );

  xor2  gate413(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate414(.a(gate123inter0), .b(s_36), .O(gate123inter1));
  and2  gate415(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate416(.a(s_36), .O(gate123inter3));
  inv1  gate417(.a(s_37), .O(gate123inter4));
  nand2 gate418(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate419(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate420(.a(N339), .O(gate123inter7));
  inv1  gate421(.a(N306), .O(gate123inter8));
  nand2 gate422(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate423(.a(s_37), .b(gate123inter3), .O(gate123inter10));
  nor2  gate424(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate425(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate426(.a(gate123inter12), .b(gate123inter1), .O(N354));
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate343(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate344(.a(gate131inter0), .b(s_26), .O(gate131inter1));
  and2  gate345(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate346(.a(s_26), .O(gate131inter3));
  inv1  gate347(.a(s_27), .O(gate131inter4));
  nand2 gate348(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate349(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate350(.a(N360), .O(gate131inter7));
  inv1  gate351(.a(N40), .O(gate131inter8));
  nand2 gate352(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate353(.a(s_27), .b(gate131inter3), .O(gate131inter10));
  nor2  gate354(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate355(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate356(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate861(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate862(.a(gate136inter0), .b(s_100), .O(gate136inter1));
  and2  gate863(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate864(.a(s_100), .O(gate136inter3));
  inv1  gate865(.a(s_101), .O(gate136inter4));
  nand2 gate866(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate867(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate868(.a(N360), .O(gate136inter7));
  inv1  gate869(.a(N105), .O(gate136inter8));
  nand2 gate870(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate871(.a(s_101), .b(gate136inter3), .O(gate136inter10));
  nor2  gate872(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate873(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate874(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate315(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate316(.a(gate153inter0), .b(s_22), .O(gate153inter1));
  and2  gate317(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate318(.a(s_22), .O(gate153inter3));
  inv1  gate319(.a(s_23), .O(gate153inter4));
  nand2 gate320(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate321(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate322(.a(N415), .O(gate153inter7));
  inv1  gate323(.a(N416), .O(gate153inter8));
  nand2 gate324(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate325(.a(s_23), .b(gate153inter3), .O(gate153inter10));
  nor2  gate326(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate327(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate328(.a(gate153inter12), .b(gate153inter1), .O(N421));

  xor2  gate469(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate470(.a(gate154inter0), .b(s_44), .O(gate154inter1));
  and2  gate471(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate472(.a(s_44), .O(gate154inter3));
  inv1  gate473(.a(s_45), .O(gate154inter4));
  nand2 gate474(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate475(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate476(.a(N386), .O(gate154inter7));
  inv1  gate477(.a(N417), .O(gate154inter8));
  nand2 gate478(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate479(.a(s_45), .b(gate154inter3), .O(gate154inter10));
  nor2  gate480(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate481(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate482(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule