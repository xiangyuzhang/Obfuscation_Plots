module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1051(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1052(.a(gate13inter0), .b(s_72), .O(gate13inter1));
  and2  gate1053(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1054(.a(s_72), .O(gate13inter3));
  inv1  gate1055(.a(s_73), .O(gate13inter4));
  nand2 gate1056(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1057(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1058(.a(G9), .O(gate13inter7));
  inv1  gate1059(.a(G10), .O(gate13inter8));
  nand2 gate1060(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1061(.a(s_73), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1062(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1063(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1064(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1471(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1472(.a(gate18inter0), .b(s_132), .O(gate18inter1));
  and2  gate1473(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1474(.a(s_132), .O(gate18inter3));
  inv1  gate1475(.a(s_133), .O(gate18inter4));
  nand2 gate1476(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1477(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1478(.a(G19), .O(gate18inter7));
  inv1  gate1479(.a(G20), .O(gate18inter8));
  nand2 gate1480(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1481(.a(s_133), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1482(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1483(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1484(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1163(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1164(.a(gate29inter0), .b(s_88), .O(gate29inter1));
  and2  gate1165(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1166(.a(s_88), .O(gate29inter3));
  inv1  gate1167(.a(s_89), .O(gate29inter4));
  nand2 gate1168(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1169(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1170(.a(G3), .O(gate29inter7));
  inv1  gate1171(.a(G7), .O(gate29inter8));
  nand2 gate1172(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1173(.a(s_89), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1174(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1175(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1176(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate953(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate954(.a(gate34inter0), .b(s_58), .O(gate34inter1));
  and2  gate955(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate956(.a(s_58), .O(gate34inter3));
  inv1  gate957(.a(s_59), .O(gate34inter4));
  nand2 gate958(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate959(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate960(.a(G25), .O(gate34inter7));
  inv1  gate961(.a(G29), .O(gate34inter8));
  nand2 gate962(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate963(.a(s_59), .b(gate34inter3), .O(gate34inter10));
  nor2  gate964(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate965(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate966(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1261(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1262(.a(gate35inter0), .b(s_102), .O(gate35inter1));
  and2  gate1263(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1264(.a(s_102), .O(gate35inter3));
  inv1  gate1265(.a(s_103), .O(gate35inter4));
  nand2 gate1266(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1267(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1268(.a(G18), .O(gate35inter7));
  inv1  gate1269(.a(G22), .O(gate35inter8));
  nand2 gate1270(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1271(.a(s_103), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1272(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1273(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1274(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate981(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate982(.a(gate38inter0), .b(s_62), .O(gate38inter1));
  and2  gate983(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate984(.a(s_62), .O(gate38inter3));
  inv1  gate985(.a(s_63), .O(gate38inter4));
  nand2 gate986(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate987(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate988(.a(G27), .O(gate38inter7));
  inv1  gate989(.a(G31), .O(gate38inter8));
  nand2 gate990(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate991(.a(s_63), .b(gate38inter3), .O(gate38inter10));
  nor2  gate992(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate993(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate994(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate645(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate646(.a(gate39inter0), .b(s_14), .O(gate39inter1));
  and2  gate647(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate648(.a(s_14), .O(gate39inter3));
  inv1  gate649(.a(s_15), .O(gate39inter4));
  nand2 gate650(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate651(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate652(.a(G20), .O(gate39inter7));
  inv1  gate653(.a(G24), .O(gate39inter8));
  nand2 gate654(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate655(.a(s_15), .b(gate39inter3), .O(gate39inter10));
  nor2  gate656(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate657(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate658(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1219(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1220(.a(gate40inter0), .b(s_96), .O(gate40inter1));
  and2  gate1221(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1222(.a(s_96), .O(gate40inter3));
  inv1  gate1223(.a(s_97), .O(gate40inter4));
  nand2 gate1224(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1225(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1226(.a(G28), .O(gate40inter7));
  inv1  gate1227(.a(G32), .O(gate40inter8));
  nand2 gate1228(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1229(.a(s_97), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1230(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1231(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1232(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate911(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate912(.a(gate46inter0), .b(s_52), .O(gate46inter1));
  and2  gate913(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate914(.a(s_52), .O(gate46inter3));
  inv1  gate915(.a(s_53), .O(gate46inter4));
  nand2 gate916(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate917(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate918(.a(G6), .O(gate46inter7));
  inv1  gate919(.a(G272), .O(gate46inter8));
  nand2 gate920(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate921(.a(s_53), .b(gate46inter3), .O(gate46inter10));
  nor2  gate922(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate923(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate924(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1597(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1598(.a(gate75inter0), .b(s_150), .O(gate75inter1));
  and2  gate1599(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1600(.a(s_150), .O(gate75inter3));
  inv1  gate1601(.a(s_151), .O(gate75inter4));
  nand2 gate1602(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1603(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1604(.a(G9), .O(gate75inter7));
  inv1  gate1605(.a(G317), .O(gate75inter8));
  nand2 gate1606(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1607(.a(s_151), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1608(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1609(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1610(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate603(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate604(.a(gate78inter0), .b(s_8), .O(gate78inter1));
  and2  gate605(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate606(.a(s_8), .O(gate78inter3));
  inv1  gate607(.a(s_9), .O(gate78inter4));
  nand2 gate608(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate609(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate610(.a(G6), .O(gate78inter7));
  inv1  gate611(.a(G320), .O(gate78inter8));
  nand2 gate612(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate613(.a(s_9), .b(gate78inter3), .O(gate78inter10));
  nor2  gate614(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate615(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate616(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1205(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1206(.a(gate82inter0), .b(s_94), .O(gate82inter1));
  and2  gate1207(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1208(.a(s_94), .O(gate82inter3));
  inv1  gate1209(.a(s_95), .O(gate82inter4));
  nand2 gate1210(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1211(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1212(.a(G7), .O(gate82inter7));
  inv1  gate1213(.a(G326), .O(gate82inter8));
  nand2 gate1214(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1215(.a(s_95), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1216(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1217(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1218(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1625(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1626(.a(gate86inter0), .b(s_154), .O(gate86inter1));
  and2  gate1627(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1628(.a(s_154), .O(gate86inter3));
  inv1  gate1629(.a(s_155), .O(gate86inter4));
  nand2 gate1630(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1631(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1632(.a(G8), .O(gate86inter7));
  inv1  gate1633(.a(G332), .O(gate86inter8));
  nand2 gate1634(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1635(.a(s_155), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1636(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1637(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1638(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1345(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1346(.a(gate87inter0), .b(s_114), .O(gate87inter1));
  and2  gate1347(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1348(.a(s_114), .O(gate87inter3));
  inv1  gate1349(.a(s_115), .O(gate87inter4));
  nand2 gate1350(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1351(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1352(.a(G12), .O(gate87inter7));
  inv1  gate1353(.a(G335), .O(gate87inter8));
  nand2 gate1354(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1355(.a(s_115), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1356(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1357(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1358(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate701(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate702(.a(gate93inter0), .b(s_22), .O(gate93inter1));
  and2  gate703(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate704(.a(s_22), .O(gate93inter3));
  inv1  gate705(.a(s_23), .O(gate93inter4));
  nand2 gate706(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate707(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate708(.a(G18), .O(gate93inter7));
  inv1  gate709(.a(G344), .O(gate93inter8));
  nand2 gate710(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate711(.a(s_23), .b(gate93inter3), .O(gate93inter10));
  nor2  gate712(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate713(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate714(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate589(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate590(.a(gate96inter0), .b(s_6), .O(gate96inter1));
  and2  gate591(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate592(.a(s_6), .O(gate96inter3));
  inv1  gate593(.a(s_7), .O(gate96inter4));
  nand2 gate594(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate595(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate596(.a(G30), .O(gate96inter7));
  inv1  gate597(.a(G347), .O(gate96inter8));
  nand2 gate598(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate599(.a(s_7), .b(gate96inter3), .O(gate96inter10));
  nor2  gate600(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate601(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate602(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1723(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1724(.a(gate101inter0), .b(s_168), .O(gate101inter1));
  and2  gate1725(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1726(.a(s_168), .O(gate101inter3));
  inv1  gate1727(.a(s_169), .O(gate101inter4));
  nand2 gate1728(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1729(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1730(.a(G20), .O(gate101inter7));
  inv1  gate1731(.a(G356), .O(gate101inter8));
  nand2 gate1732(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1733(.a(s_169), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1734(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1735(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1736(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1317(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1318(.a(gate107inter0), .b(s_110), .O(gate107inter1));
  and2  gate1319(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1320(.a(s_110), .O(gate107inter3));
  inv1  gate1321(.a(s_111), .O(gate107inter4));
  nand2 gate1322(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1323(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1324(.a(G366), .O(gate107inter7));
  inv1  gate1325(.a(G367), .O(gate107inter8));
  nand2 gate1326(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1327(.a(s_111), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1328(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1329(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1330(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1093(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1094(.a(gate108inter0), .b(s_78), .O(gate108inter1));
  and2  gate1095(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1096(.a(s_78), .O(gate108inter3));
  inv1  gate1097(.a(s_79), .O(gate108inter4));
  nand2 gate1098(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1099(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1100(.a(G368), .O(gate108inter7));
  inv1  gate1101(.a(G369), .O(gate108inter8));
  nand2 gate1102(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1103(.a(s_79), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1104(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1105(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1106(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate939(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate940(.a(gate110inter0), .b(s_56), .O(gate110inter1));
  and2  gate941(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate942(.a(s_56), .O(gate110inter3));
  inv1  gate943(.a(s_57), .O(gate110inter4));
  nand2 gate944(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate945(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate946(.a(G372), .O(gate110inter7));
  inv1  gate947(.a(G373), .O(gate110inter8));
  nand2 gate948(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate949(.a(s_57), .b(gate110inter3), .O(gate110inter10));
  nor2  gate950(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate951(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate952(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1443(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1444(.a(gate111inter0), .b(s_128), .O(gate111inter1));
  and2  gate1445(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1446(.a(s_128), .O(gate111inter3));
  inv1  gate1447(.a(s_129), .O(gate111inter4));
  nand2 gate1448(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1449(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1450(.a(G374), .O(gate111inter7));
  inv1  gate1451(.a(G375), .O(gate111inter8));
  nand2 gate1452(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1453(.a(s_129), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1454(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1455(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1456(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1275(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1276(.a(gate119inter0), .b(s_104), .O(gate119inter1));
  and2  gate1277(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1278(.a(s_104), .O(gate119inter3));
  inv1  gate1279(.a(s_105), .O(gate119inter4));
  nand2 gate1280(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1281(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1282(.a(G390), .O(gate119inter7));
  inv1  gate1283(.a(G391), .O(gate119inter8));
  nand2 gate1284(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1285(.a(s_105), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1286(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1287(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1288(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1737(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1738(.a(gate123inter0), .b(s_170), .O(gate123inter1));
  and2  gate1739(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1740(.a(s_170), .O(gate123inter3));
  inv1  gate1741(.a(s_171), .O(gate123inter4));
  nand2 gate1742(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1743(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1744(.a(G398), .O(gate123inter7));
  inv1  gate1745(.a(G399), .O(gate123inter8));
  nand2 gate1746(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1747(.a(s_171), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1748(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1749(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1750(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1247(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1248(.a(gate127inter0), .b(s_100), .O(gate127inter1));
  and2  gate1249(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1250(.a(s_100), .O(gate127inter3));
  inv1  gate1251(.a(s_101), .O(gate127inter4));
  nand2 gate1252(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1253(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1254(.a(G406), .O(gate127inter7));
  inv1  gate1255(.a(G407), .O(gate127inter8));
  nand2 gate1256(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1257(.a(s_101), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1258(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1259(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1260(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate813(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate814(.a(gate133inter0), .b(s_38), .O(gate133inter1));
  and2  gate815(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate816(.a(s_38), .O(gate133inter3));
  inv1  gate817(.a(s_39), .O(gate133inter4));
  nand2 gate818(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate819(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate820(.a(G418), .O(gate133inter7));
  inv1  gate821(.a(G419), .O(gate133inter8));
  nand2 gate822(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate823(.a(s_39), .b(gate133inter3), .O(gate133inter10));
  nor2  gate824(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate825(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate826(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1065(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1066(.a(gate135inter0), .b(s_74), .O(gate135inter1));
  and2  gate1067(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1068(.a(s_74), .O(gate135inter3));
  inv1  gate1069(.a(s_75), .O(gate135inter4));
  nand2 gate1070(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1071(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1072(.a(G422), .O(gate135inter7));
  inv1  gate1073(.a(G423), .O(gate135inter8));
  nand2 gate1074(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1075(.a(s_75), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1076(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1077(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1078(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1135(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1136(.a(gate137inter0), .b(s_84), .O(gate137inter1));
  and2  gate1137(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1138(.a(s_84), .O(gate137inter3));
  inv1  gate1139(.a(s_85), .O(gate137inter4));
  nand2 gate1140(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1141(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1142(.a(G426), .O(gate137inter7));
  inv1  gate1143(.a(G429), .O(gate137inter8));
  nand2 gate1144(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1145(.a(s_85), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1146(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1147(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1148(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate841(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate842(.a(gate151inter0), .b(s_42), .O(gate151inter1));
  and2  gate843(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate844(.a(s_42), .O(gate151inter3));
  inv1  gate845(.a(s_43), .O(gate151inter4));
  nand2 gate846(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate847(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate848(.a(G510), .O(gate151inter7));
  inv1  gate849(.a(G513), .O(gate151inter8));
  nand2 gate850(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate851(.a(s_43), .b(gate151inter3), .O(gate151inter10));
  nor2  gate852(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate853(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate854(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate883(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate884(.a(gate153inter0), .b(s_48), .O(gate153inter1));
  and2  gate885(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate886(.a(s_48), .O(gate153inter3));
  inv1  gate887(.a(s_49), .O(gate153inter4));
  nand2 gate888(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate889(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate890(.a(G426), .O(gate153inter7));
  inv1  gate891(.a(G522), .O(gate153inter8));
  nand2 gate892(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate893(.a(s_49), .b(gate153inter3), .O(gate153inter10));
  nor2  gate894(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate895(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate896(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1639(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1640(.a(gate166inter0), .b(s_156), .O(gate166inter1));
  and2  gate1641(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1642(.a(s_156), .O(gate166inter3));
  inv1  gate1643(.a(s_157), .O(gate166inter4));
  nand2 gate1644(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1645(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1646(.a(G465), .O(gate166inter7));
  inv1  gate1647(.a(G540), .O(gate166inter8));
  nand2 gate1648(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1649(.a(s_157), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1650(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1651(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1652(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1009(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1010(.a(gate168inter0), .b(s_66), .O(gate168inter1));
  and2  gate1011(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1012(.a(s_66), .O(gate168inter3));
  inv1  gate1013(.a(s_67), .O(gate168inter4));
  nand2 gate1014(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1015(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1016(.a(G471), .O(gate168inter7));
  inv1  gate1017(.a(G543), .O(gate168inter8));
  nand2 gate1018(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1019(.a(s_67), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1020(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1021(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1022(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1401(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1402(.a(gate173inter0), .b(s_122), .O(gate173inter1));
  and2  gate1403(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1404(.a(s_122), .O(gate173inter3));
  inv1  gate1405(.a(s_123), .O(gate173inter4));
  nand2 gate1406(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1407(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1408(.a(G486), .O(gate173inter7));
  inv1  gate1409(.a(G552), .O(gate173inter8));
  nand2 gate1410(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1411(.a(s_123), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1412(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1413(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1414(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate757(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate758(.a(gate174inter0), .b(s_30), .O(gate174inter1));
  and2  gate759(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate760(.a(s_30), .O(gate174inter3));
  inv1  gate761(.a(s_31), .O(gate174inter4));
  nand2 gate762(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate763(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate764(.a(G489), .O(gate174inter7));
  inv1  gate765(.a(G552), .O(gate174inter8));
  nand2 gate766(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate767(.a(s_31), .b(gate174inter3), .O(gate174inter10));
  nor2  gate768(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate769(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate770(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate771(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate772(.a(gate176inter0), .b(s_32), .O(gate176inter1));
  and2  gate773(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate774(.a(s_32), .O(gate176inter3));
  inv1  gate775(.a(s_33), .O(gate176inter4));
  nand2 gate776(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate777(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate778(.a(G495), .O(gate176inter7));
  inv1  gate779(.a(G555), .O(gate176inter8));
  nand2 gate780(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate781(.a(s_33), .b(gate176inter3), .O(gate176inter10));
  nor2  gate782(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate783(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate784(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1667(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1668(.a(gate186inter0), .b(s_160), .O(gate186inter1));
  and2  gate1669(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1670(.a(s_160), .O(gate186inter3));
  inv1  gate1671(.a(s_161), .O(gate186inter4));
  nand2 gate1672(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1673(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1674(.a(G572), .O(gate186inter7));
  inv1  gate1675(.a(G573), .O(gate186inter8));
  nand2 gate1676(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1677(.a(s_161), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1678(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1679(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1680(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1485(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1486(.a(gate187inter0), .b(s_134), .O(gate187inter1));
  and2  gate1487(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1488(.a(s_134), .O(gate187inter3));
  inv1  gate1489(.a(s_135), .O(gate187inter4));
  nand2 gate1490(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1491(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1492(.a(G574), .O(gate187inter7));
  inv1  gate1493(.a(G575), .O(gate187inter8));
  nand2 gate1494(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1495(.a(s_135), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1496(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1497(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1498(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate967(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate968(.a(gate188inter0), .b(s_60), .O(gate188inter1));
  and2  gate969(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate970(.a(s_60), .O(gate188inter3));
  inv1  gate971(.a(s_61), .O(gate188inter4));
  nand2 gate972(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate973(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate974(.a(G576), .O(gate188inter7));
  inv1  gate975(.a(G577), .O(gate188inter8));
  nand2 gate976(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate977(.a(s_61), .b(gate188inter3), .O(gate188inter10));
  nor2  gate978(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate979(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate980(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate897(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate898(.a(gate198inter0), .b(s_50), .O(gate198inter1));
  and2  gate899(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate900(.a(s_50), .O(gate198inter3));
  inv1  gate901(.a(s_51), .O(gate198inter4));
  nand2 gate902(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate903(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate904(.a(G596), .O(gate198inter7));
  inv1  gate905(.a(G597), .O(gate198inter8));
  nand2 gate906(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate907(.a(s_51), .b(gate198inter3), .O(gate198inter10));
  nor2  gate908(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate909(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate910(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1513(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1514(.a(gate200inter0), .b(s_138), .O(gate200inter1));
  and2  gate1515(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1516(.a(s_138), .O(gate200inter3));
  inv1  gate1517(.a(s_139), .O(gate200inter4));
  nand2 gate1518(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1519(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1520(.a(G600), .O(gate200inter7));
  inv1  gate1521(.a(G601), .O(gate200inter8));
  nand2 gate1522(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1523(.a(s_139), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1524(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1525(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1526(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate631(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate632(.a(gate202inter0), .b(s_12), .O(gate202inter1));
  and2  gate633(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate634(.a(s_12), .O(gate202inter3));
  inv1  gate635(.a(s_13), .O(gate202inter4));
  nand2 gate636(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate637(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate638(.a(G612), .O(gate202inter7));
  inv1  gate639(.a(G617), .O(gate202inter8));
  nand2 gate640(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate641(.a(s_13), .b(gate202inter3), .O(gate202inter10));
  nor2  gate642(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate643(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate644(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1079(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1080(.a(gate207inter0), .b(s_76), .O(gate207inter1));
  and2  gate1081(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1082(.a(s_76), .O(gate207inter3));
  inv1  gate1083(.a(s_77), .O(gate207inter4));
  nand2 gate1084(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1085(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1086(.a(G622), .O(gate207inter7));
  inv1  gate1087(.a(G632), .O(gate207inter8));
  nand2 gate1088(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1089(.a(s_77), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1090(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1091(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1092(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1373(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1374(.a(gate223inter0), .b(s_118), .O(gate223inter1));
  and2  gate1375(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1376(.a(s_118), .O(gate223inter3));
  inv1  gate1377(.a(s_119), .O(gate223inter4));
  nand2 gate1378(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1379(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1380(.a(G627), .O(gate223inter7));
  inv1  gate1381(.a(G687), .O(gate223inter8));
  nand2 gate1382(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1383(.a(s_119), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1384(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1385(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1386(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate827(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate828(.a(gate229inter0), .b(s_40), .O(gate229inter1));
  and2  gate829(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate830(.a(s_40), .O(gate229inter3));
  inv1  gate831(.a(s_41), .O(gate229inter4));
  nand2 gate832(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate833(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate834(.a(G698), .O(gate229inter7));
  inv1  gate835(.a(G699), .O(gate229inter8));
  nand2 gate836(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate837(.a(s_41), .b(gate229inter3), .O(gate229inter10));
  nor2  gate838(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate839(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate840(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1457(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1458(.a(gate236inter0), .b(s_130), .O(gate236inter1));
  and2  gate1459(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1460(.a(s_130), .O(gate236inter3));
  inv1  gate1461(.a(s_131), .O(gate236inter4));
  nand2 gate1462(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1463(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1464(.a(G251), .O(gate236inter7));
  inv1  gate1465(.a(G727), .O(gate236inter8));
  nand2 gate1466(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1467(.a(s_131), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1468(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1469(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1470(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1023(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1024(.a(gate238inter0), .b(s_68), .O(gate238inter1));
  and2  gate1025(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1026(.a(s_68), .O(gate238inter3));
  inv1  gate1027(.a(s_69), .O(gate238inter4));
  nand2 gate1028(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1029(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1030(.a(G257), .O(gate238inter7));
  inv1  gate1031(.a(G709), .O(gate238inter8));
  nand2 gate1032(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1033(.a(s_69), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1034(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1035(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1036(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1583(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1584(.a(gate240inter0), .b(s_148), .O(gate240inter1));
  and2  gate1585(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1586(.a(s_148), .O(gate240inter3));
  inv1  gate1587(.a(s_149), .O(gate240inter4));
  nand2 gate1588(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1589(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1590(.a(G263), .O(gate240inter7));
  inv1  gate1591(.a(G715), .O(gate240inter8));
  nand2 gate1592(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1593(.a(s_149), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1594(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1595(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1596(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1499(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1500(.a(gate241inter0), .b(s_136), .O(gate241inter1));
  and2  gate1501(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1502(.a(s_136), .O(gate241inter3));
  inv1  gate1503(.a(s_137), .O(gate241inter4));
  nand2 gate1504(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1505(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1506(.a(G242), .O(gate241inter7));
  inv1  gate1507(.a(G730), .O(gate241inter8));
  nand2 gate1508(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1509(.a(s_137), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1510(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1511(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1512(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate925(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate926(.a(gate249inter0), .b(s_54), .O(gate249inter1));
  and2  gate927(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate928(.a(s_54), .O(gate249inter3));
  inv1  gate929(.a(s_55), .O(gate249inter4));
  nand2 gate930(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate931(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate932(.a(G254), .O(gate249inter7));
  inv1  gate933(.a(G742), .O(gate249inter8));
  nand2 gate934(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate935(.a(s_55), .b(gate249inter3), .O(gate249inter10));
  nor2  gate936(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate937(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate938(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate729(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate730(.a(gate252inter0), .b(s_26), .O(gate252inter1));
  and2  gate731(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate732(.a(s_26), .O(gate252inter3));
  inv1  gate733(.a(s_27), .O(gate252inter4));
  nand2 gate734(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate735(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate736(.a(G709), .O(gate252inter7));
  inv1  gate737(.a(G745), .O(gate252inter8));
  nand2 gate738(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate739(.a(s_27), .b(gate252inter3), .O(gate252inter10));
  nor2  gate740(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate741(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate742(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1359(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1360(.a(gate264inter0), .b(s_116), .O(gate264inter1));
  and2  gate1361(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1362(.a(s_116), .O(gate264inter3));
  inv1  gate1363(.a(s_117), .O(gate264inter4));
  nand2 gate1364(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1365(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1366(.a(G768), .O(gate264inter7));
  inv1  gate1367(.a(G769), .O(gate264inter8));
  nand2 gate1368(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1369(.a(s_117), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1370(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1371(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1372(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1569(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1570(.a(gate266inter0), .b(s_146), .O(gate266inter1));
  and2  gate1571(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1572(.a(s_146), .O(gate266inter3));
  inv1  gate1573(.a(s_147), .O(gate266inter4));
  nand2 gate1574(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1575(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1576(.a(G645), .O(gate266inter7));
  inv1  gate1577(.a(G773), .O(gate266inter8));
  nand2 gate1578(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1579(.a(s_147), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1580(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1581(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1582(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1429(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1430(.a(gate269inter0), .b(s_126), .O(gate269inter1));
  and2  gate1431(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1432(.a(s_126), .O(gate269inter3));
  inv1  gate1433(.a(s_127), .O(gate269inter4));
  nand2 gate1434(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1435(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1436(.a(G654), .O(gate269inter7));
  inv1  gate1437(.a(G782), .O(gate269inter8));
  nand2 gate1438(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1439(.a(s_127), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1440(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1441(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1442(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate659(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate660(.a(gate271inter0), .b(s_16), .O(gate271inter1));
  and2  gate661(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate662(.a(s_16), .O(gate271inter3));
  inv1  gate663(.a(s_17), .O(gate271inter4));
  nand2 gate664(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate665(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate666(.a(G660), .O(gate271inter7));
  inv1  gate667(.a(G788), .O(gate271inter8));
  nand2 gate668(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate669(.a(s_17), .b(gate271inter3), .O(gate271inter10));
  nor2  gate670(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate671(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate672(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1303(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1304(.a(gate274inter0), .b(s_108), .O(gate274inter1));
  and2  gate1305(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1306(.a(s_108), .O(gate274inter3));
  inv1  gate1307(.a(s_109), .O(gate274inter4));
  nand2 gate1308(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1309(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1310(.a(G770), .O(gate274inter7));
  inv1  gate1311(.a(G794), .O(gate274inter8));
  nand2 gate1312(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1313(.a(s_109), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1314(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1315(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1316(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate785(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate786(.a(gate277inter0), .b(s_34), .O(gate277inter1));
  and2  gate787(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate788(.a(s_34), .O(gate277inter3));
  inv1  gate789(.a(s_35), .O(gate277inter4));
  nand2 gate790(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate791(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate792(.a(G648), .O(gate277inter7));
  inv1  gate793(.a(G800), .O(gate277inter8));
  nand2 gate794(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate795(.a(s_35), .b(gate277inter3), .O(gate277inter10));
  nor2  gate796(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate797(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate798(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1191(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1192(.a(gate288inter0), .b(s_92), .O(gate288inter1));
  and2  gate1193(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1194(.a(s_92), .O(gate288inter3));
  inv1  gate1195(.a(s_93), .O(gate288inter4));
  nand2 gate1196(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1197(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1198(.a(G791), .O(gate288inter7));
  inv1  gate1199(.a(G815), .O(gate288inter8));
  nand2 gate1200(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1201(.a(s_93), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1202(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1203(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1204(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1177(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1178(.a(gate291inter0), .b(s_90), .O(gate291inter1));
  and2  gate1179(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1180(.a(s_90), .O(gate291inter3));
  inv1  gate1181(.a(s_91), .O(gate291inter4));
  nand2 gate1182(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1183(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1184(.a(G822), .O(gate291inter7));
  inv1  gate1185(.a(G823), .O(gate291inter8));
  nand2 gate1186(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1187(.a(s_91), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1188(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1189(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1190(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1233(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1234(.a(gate295inter0), .b(s_98), .O(gate295inter1));
  and2  gate1235(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1236(.a(s_98), .O(gate295inter3));
  inv1  gate1237(.a(s_99), .O(gate295inter4));
  nand2 gate1238(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1239(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1240(.a(G830), .O(gate295inter7));
  inv1  gate1241(.a(G831), .O(gate295inter8));
  nand2 gate1242(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1243(.a(s_99), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1244(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1245(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1246(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1331(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1332(.a(gate296inter0), .b(s_112), .O(gate296inter1));
  and2  gate1333(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1334(.a(s_112), .O(gate296inter3));
  inv1  gate1335(.a(s_113), .O(gate296inter4));
  nand2 gate1336(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1337(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1338(.a(G826), .O(gate296inter7));
  inv1  gate1339(.a(G827), .O(gate296inter8));
  nand2 gate1340(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1341(.a(s_113), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1342(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1343(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1344(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1149(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1150(.a(gate387inter0), .b(s_86), .O(gate387inter1));
  and2  gate1151(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1152(.a(s_86), .O(gate387inter3));
  inv1  gate1153(.a(s_87), .O(gate387inter4));
  nand2 gate1154(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1155(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1156(.a(G1), .O(gate387inter7));
  inv1  gate1157(.a(G1036), .O(gate387inter8));
  nand2 gate1158(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1159(.a(s_87), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1160(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1161(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1162(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1387(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1388(.a(gate396inter0), .b(s_120), .O(gate396inter1));
  and2  gate1389(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1390(.a(s_120), .O(gate396inter3));
  inv1  gate1391(.a(s_121), .O(gate396inter4));
  nand2 gate1392(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1393(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1394(.a(G10), .O(gate396inter7));
  inv1  gate1395(.a(G1063), .O(gate396inter8));
  nand2 gate1396(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1397(.a(s_121), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1398(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1399(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1400(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1107(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1108(.a(gate399inter0), .b(s_80), .O(gate399inter1));
  and2  gate1109(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1110(.a(s_80), .O(gate399inter3));
  inv1  gate1111(.a(s_81), .O(gate399inter4));
  nand2 gate1112(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1113(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1114(.a(G13), .O(gate399inter7));
  inv1  gate1115(.a(G1072), .O(gate399inter8));
  nand2 gate1116(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1117(.a(s_81), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1118(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1119(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1120(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate547(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate548(.a(gate403inter0), .b(s_0), .O(gate403inter1));
  and2  gate549(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate550(.a(s_0), .O(gate403inter3));
  inv1  gate551(.a(s_1), .O(gate403inter4));
  nand2 gate552(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate553(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate554(.a(G17), .O(gate403inter7));
  inv1  gate555(.a(G1084), .O(gate403inter8));
  nand2 gate556(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate557(.a(s_1), .b(gate403inter3), .O(gate403inter10));
  nor2  gate558(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate559(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate560(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1541(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1542(.a(gate407inter0), .b(s_142), .O(gate407inter1));
  and2  gate1543(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1544(.a(s_142), .O(gate407inter3));
  inv1  gate1545(.a(s_143), .O(gate407inter4));
  nand2 gate1546(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1547(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1548(.a(G21), .O(gate407inter7));
  inv1  gate1549(.a(G1096), .O(gate407inter8));
  nand2 gate1550(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1551(.a(s_143), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1552(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1553(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1554(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate673(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate674(.a(gate418inter0), .b(s_18), .O(gate418inter1));
  and2  gate675(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate676(.a(s_18), .O(gate418inter3));
  inv1  gate677(.a(s_19), .O(gate418inter4));
  nand2 gate678(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate679(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate680(.a(G32), .O(gate418inter7));
  inv1  gate681(.a(G1129), .O(gate418inter8));
  nand2 gate682(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate683(.a(s_19), .b(gate418inter3), .O(gate418inter10));
  nor2  gate684(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate685(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate686(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1695(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1696(.a(gate420inter0), .b(s_164), .O(gate420inter1));
  and2  gate1697(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1698(.a(s_164), .O(gate420inter3));
  inv1  gate1699(.a(s_165), .O(gate420inter4));
  nand2 gate1700(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1701(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1702(.a(G1036), .O(gate420inter7));
  inv1  gate1703(.a(G1132), .O(gate420inter8));
  nand2 gate1704(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1705(.a(s_165), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1706(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1707(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1708(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1121(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1122(.a(gate422inter0), .b(s_82), .O(gate422inter1));
  and2  gate1123(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1124(.a(s_82), .O(gate422inter3));
  inv1  gate1125(.a(s_83), .O(gate422inter4));
  nand2 gate1126(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1127(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1128(.a(G1039), .O(gate422inter7));
  inv1  gate1129(.a(G1135), .O(gate422inter8));
  nand2 gate1130(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1131(.a(s_83), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1132(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1133(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1134(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1415(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1416(.a(gate428inter0), .b(s_124), .O(gate428inter1));
  and2  gate1417(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1418(.a(s_124), .O(gate428inter3));
  inv1  gate1419(.a(s_125), .O(gate428inter4));
  nand2 gate1420(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1421(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1422(.a(G1048), .O(gate428inter7));
  inv1  gate1423(.a(G1144), .O(gate428inter8));
  nand2 gate1424(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1425(.a(s_125), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1426(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1427(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1428(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1527(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1528(.a(gate430inter0), .b(s_140), .O(gate430inter1));
  and2  gate1529(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1530(.a(s_140), .O(gate430inter3));
  inv1  gate1531(.a(s_141), .O(gate430inter4));
  nand2 gate1532(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1533(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1534(.a(G1051), .O(gate430inter7));
  inv1  gate1535(.a(G1147), .O(gate430inter8));
  nand2 gate1536(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1537(.a(s_141), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1538(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1539(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1540(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate575(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate576(.a(gate434inter0), .b(s_4), .O(gate434inter1));
  and2  gate577(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate578(.a(s_4), .O(gate434inter3));
  inv1  gate579(.a(s_5), .O(gate434inter4));
  nand2 gate580(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate581(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate582(.a(G1057), .O(gate434inter7));
  inv1  gate583(.a(G1153), .O(gate434inter8));
  nand2 gate584(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate585(.a(s_5), .b(gate434inter3), .O(gate434inter10));
  nor2  gate586(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate587(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate588(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate715(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate716(.a(gate436inter0), .b(s_24), .O(gate436inter1));
  and2  gate717(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate718(.a(s_24), .O(gate436inter3));
  inv1  gate719(.a(s_25), .O(gate436inter4));
  nand2 gate720(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate721(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate722(.a(G1060), .O(gate436inter7));
  inv1  gate723(.a(G1156), .O(gate436inter8));
  nand2 gate724(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate725(.a(s_25), .b(gate436inter3), .O(gate436inter10));
  nor2  gate726(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate727(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate728(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1289(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1290(.a(gate438inter0), .b(s_106), .O(gate438inter1));
  and2  gate1291(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1292(.a(s_106), .O(gate438inter3));
  inv1  gate1293(.a(s_107), .O(gate438inter4));
  nand2 gate1294(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1295(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1296(.a(G1063), .O(gate438inter7));
  inv1  gate1297(.a(G1159), .O(gate438inter8));
  nand2 gate1298(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1299(.a(s_107), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1300(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1301(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1302(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate687(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate688(.a(gate439inter0), .b(s_20), .O(gate439inter1));
  and2  gate689(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate690(.a(s_20), .O(gate439inter3));
  inv1  gate691(.a(s_21), .O(gate439inter4));
  nand2 gate692(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate693(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate694(.a(G11), .O(gate439inter7));
  inv1  gate695(.a(G1162), .O(gate439inter8));
  nand2 gate696(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate697(.a(s_21), .b(gate439inter3), .O(gate439inter10));
  nor2  gate698(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate699(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate700(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate869(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate870(.a(gate448inter0), .b(s_46), .O(gate448inter1));
  and2  gate871(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate872(.a(s_46), .O(gate448inter3));
  inv1  gate873(.a(s_47), .O(gate448inter4));
  nand2 gate874(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate875(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate876(.a(G1078), .O(gate448inter7));
  inv1  gate877(.a(G1174), .O(gate448inter8));
  nand2 gate878(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate879(.a(s_47), .b(gate448inter3), .O(gate448inter10));
  nor2  gate880(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate881(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate882(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1681(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1682(.a(gate450inter0), .b(s_162), .O(gate450inter1));
  and2  gate1683(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1684(.a(s_162), .O(gate450inter3));
  inv1  gate1685(.a(s_163), .O(gate450inter4));
  nand2 gate1686(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1687(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1688(.a(G1081), .O(gate450inter7));
  inv1  gate1689(.a(G1177), .O(gate450inter8));
  nand2 gate1690(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1691(.a(s_163), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1692(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1693(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1694(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate561(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate562(.a(gate457inter0), .b(s_2), .O(gate457inter1));
  and2  gate563(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate564(.a(s_2), .O(gate457inter3));
  inv1  gate565(.a(s_3), .O(gate457inter4));
  nand2 gate566(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate567(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate568(.a(G20), .O(gate457inter7));
  inv1  gate569(.a(G1189), .O(gate457inter8));
  nand2 gate570(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate571(.a(s_3), .b(gate457inter3), .O(gate457inter10));
  nor2  gate572(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate573(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate574(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate995(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate996(.a(gate461inter0), .b(s_64), .O(gate461inter1));
  and2  gate997(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate998(.a(s_64), .O(gate461inter3));
  inv1  gate999(.a(s_65), .O(gate461inter4));
  nand2 gate1000(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1001(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1002(.a(G22), .O(gate461inter7));
  inv1  gate1003(.a(G1195), .O(gate461inter8));
  nand2 gate1004(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1005(.a(s_65), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1006(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1007(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1008(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1037(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1038(.a(gate466inter0), .b(s_70), .O(gate466inter1));
  and2  gate1039(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1040(.a(s_70), .O(gate466inter3));
  inv1  gate1041(.a(s_71), .O(gate466inter4));
  nand2 gate1042(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1043(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1044(.a(G1105), .O(gate466inter7));
  inv1  gate1045(.a(G1201), .O(gate466inter8));
  nand2 gate1046(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1047(.a(s_71), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1048(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1049(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1050(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate799(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate800(.a(gate475inter0), .b(s_36), .O(gate475inter1));
  and2  gate801(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate802(.a(s_36), .O(gate475inter3));
  inv1  gate803(.a(s_37), .O(gate475inter4));
  nand2 gate804(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate805(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate806(.a(G29), .O(gate475inter7));
  inv1  gate807(.a(G1216), .O(gate475inter8));
  nand2 gate808(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate809(.a(s_37), .b(gate475inter3), .O(gate475inter10));
  nor2  gate810(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate811(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate812(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1611(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1612(.a(gate477inter0), .b(s_152), .O(gate477inter1));
  and2  gate1613(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1614(.a(s_152), .O(gate477inter3));
  inv1  gate1615(.a(s_153), .O(gate477inter4));
  nand2 gate1616(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1617(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1618(.a(G30), .O(gate477inter7));
  inv1  gate1619(.a(G1219), .O(gate477inter8));
  nand2 gate1620(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1621(.a(s_153), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1622(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1623(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1624(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1653(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1654(.a(gate489inter0), .b(s_158), .O(gate489inter1));
  and2  gate1655(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1656(.a(s_158), .O(gate489inter3));
  inv1  gate1657(.a(s_159), .O(gate489inter4));
  nand2 gate1658(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1659(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1660(.a(G1240), .O(gate489inter7));
  inv1  gate1661(.a(G1241), .O(gate489inter8));
  nand2 gate1662(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1663(.a(s_159), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1664(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1665(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1666(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate743(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate744(.a(gate498inter0), .b(s_28), .O(gate498inter1));
  and2  gate745(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate746(.a(s_28), .O(gate498inter3));
  inv1  gate747(.a(s_29), .O(gate498inter4));
  nand2 gate748(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate749(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate750(.a(G1258), .O(gate498inter7));
  inv1  gate751(.a(G1259), .O(gate498inter8));
  nand2 gate752(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate753(.a(s_29), .b(gate498inter3), .O(gate498inter10));
  nor2  gate754(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate755(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate756(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1709(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1710(.a(gate506inter0), .b(s_166), .O(gate506inter1));
  and2  gate1711(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1712(.a(s_166), .O(gate506inter3));
  inv1  gate1713(.a(s_167), .O(gate506inter4));
  nand2 gate1714(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1715(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1716(.a(G1274), .O(gate506inter7));
  inv1  gate1717(.a(G1275), .O(gate506inter8));
  nand2 gate1718(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1719(.a(s_167), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1720(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1721(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1722(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1555(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1556(.a(gate508inter0), .b(s_144), .O(gate508inter1));
  and2  gate1557(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1558(.a(s_144), .O(gate508inter3));
  inv1  gate1559(.a(s_145), .O(gate508inter4));
  nand2 gate1560(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1561(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1562(.a(G1278), .O(gate508inter7));
  inv1  gate1563(.a(G1279), .O(gate508inter8));
  nand2 gate1564(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1565(.a(s_145), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1566(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1567(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1568(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate855(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate856(.a(gate510inter0), .b(s_44), .O(gate510inter1));
  and2  gate857(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate858(.a(s_44), .O(gate510inter3));
  inv1  gate859(.a(s_45), .O(gate510inter4));
  nand2 gate860(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate861(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate862(.a(G1282), .O(gate510inter7));
  inv1  gate863(.a(G1283), .O(gate510inter8));
  nand2 gate864(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate865(.a(s_45), .b(gate510inter3), .O(gate510inter10));
  nor2  gate866(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate867(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate868(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate617(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate618(.a(gate512inter0), .b(s_10), .O(gate512inter1));
  and2  gate619(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate620(.a(s_10), .O(gate512inter3));
  inv1  gate621(.a(s_11), .O(gate512inter4));
  nand2 gate622(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate623(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate624(.a(G1286), .O(gate512inter7));
  inv1  gate625(.a(G1287), .O(gate512inter8));
  nand2 gate626(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate627(.a(s_11), .b(gate512inter3), .O(gate512inter10));
  nor2  gate628(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate629(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate630(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule