module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate441(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate442(.a(gate6inter0), .b(s_34), .O(gate6inter1));
  and2  gate443(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate444(.a(s_34), .O(gate6inter3));
  inv1  gate445(.a(s_35), .O(gate6inter4));
  nand2 gate446(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate447(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate448(.a(N41), .O(gate6inter7));
  inv1  gate449(.a(N45), .O(gate6inter8));
  nand2 gate450(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate451(.a(s_35), .b(gate6inter3), .O(gate6inter10));
  nor2  gate452(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate453(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate454(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );

  xor2  gate413(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate414(.a(gate10inter0), .b(s_30), .O(gate10inter1));
  and2  gate415(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate416(.a(s_30), .O(gate10inter3));
  inv1  gate417(.a(s_31), .O(gate10inter4));
  nand2 gate418(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate419(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate420(.a(N73), .O(gate10inter7));
  inv1  gate421(.a(N77), .O(gate10inter8));
  nand2 gate422(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate423(.a(s_31), .b(gate10inter3), .O(gate10inter10));
  nor2  gate424(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate425(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate426(.a(gate10inter12), .b(gate10inter1), .O(N259));
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );

  xor2  gate273(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate274(.a(gate16inter0), .b(s_10), .O(gate16inter1));
  and2  gate275(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate276(.a(s_10), .O(gate16inter3));
  inv1  gate277(.a(s_11), .O(gate16inter4));
  nand2 gate278(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate279(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate280(.a(N121), .O(gate16inter7));
  inv1  gate281(.a(N125), .O(gate16inter8));
  nand2 gate282(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate283(.a(s_11), .b(gate16inter3), .O(gate16inter10));
  nor2  gate284(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate285(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate286(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate329(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate330(.a(gate25inter0), .b(s_18), .O(gate25inter1));
  and2  gate331(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate332(.a(s_18), .O(gate25inter3));
  inv1  gate333(.a(s_19), .O(gate25inter4));
  nand2 gate334(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate335(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate336(.a(N1), .O(gate25inter7));
  inv1  gate337(.a(N17), .O(gate25inter8));
  nand2 gate338(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate339(.a(s_19), .b(gate25inter3), .O(gate25inter10));
  nor2  gate340(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate341(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate342(.a(gate25inter12), .b(gate25inter1), .O(N274));
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );

  xor2  gate315(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate316(.a(gate31inter0), .b(s_16), .O(gate31inter1));
  and2  gate317(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate318(.a(s_16), .O(gate31inter3));
  inv1  gate319(.a(s_17), .O(gate31inter4));
  nand2 gate320(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate321(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate322(.a(N13), .O(gate31inter7));
  inv1  gate323(.a(N29), .O(gate31inter8));
  nand2 gate324(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate325(.a(s_17), .b(gate31inter3), .O(gate31inter10));
  nor2  gate326(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate327(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate328(.a(gate31inter12), .b(gate31inter1), .O(N280));
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );

  xor2  gate301(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate302(.a(gate36inter0), .b(s_14), .O(gate36inter1));
  and2  gate303(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate304(.a(s_14), .O(gate36inter3));
  inv1  gate305(.a(s_15), .O(gate36inter4));
  nand2 gate306(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate307(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate308(.a(N101), .O(gate36inter7));
  inv1  gate309(.a(N117), .O(gate36inter8));
  nand2 gate310(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate311(.a(s_15), .b(gate36inter3), .O(gate36inter10));
  nor2  gate312(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate313(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate314(.a(gate36inter12), .b(gate36inter1), .O(N285));
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );

  xor2  gate469(.a(N93), .b(N77), .O(gate39inter0));
  nand2 gate470(.a(gate39inter0), .b(s_38), .O(gate39inter1));
  and2  gate471(.a(N93), .b(N77), .O(gate39inter2));
  inv1  gate472(.a(s_38), .O(gate39inter3));
  inv1  gate473(.a(s_39), .O(gate39inter4));
  nand2 gate474(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate475(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate476(.a(N77), .O(gate39inter7));
  inv1  gate477(.a(N93), .O(gate39inter8));
  nand2 gate478(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate479(.a(s_39), .b(gate39inter3), .O(gate39inter10));
  nor2  gate480(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate481(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate482(.a(gate39inter12), .b(gate39inter1), .O(N288));

  xor2  gate399(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate400(.a(gate40inter0), .b(s_28), .O(gate40inter1));
  and2  gate401(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate402(.a(s_28), .O(gate40inter3));
  inv1  gate403(.a(s_29), .O(gate40inter4));
  nand2 gate404(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate405(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate406(.a(N109), .O(gate40inter7));
  inv1  gate407(.a(N125), .O(gate40inter8));
  nand2 gate408(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate409(.a(s_29), .b(gate40inter3), .O(gate40inter10));
  nor2  gate410(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate411(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate412(.a(gate40inter12), .b(gate40inter1), .O(N289));
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );

  xor2  gate371(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate372(.a(gate49inter0), .b(s_24), .O(gate49inter1));
  and2  gate373(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate374(.a(s_24), .O(gate49inter3));
  inv1  gate375(.a(s_25), .O(gate49inter4));
  nand2 gate376(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate377(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate378(.a(N274), .O(gate49inter7));
  inv1  gate379(.a(N275), .O(gate49inter8));
  nand2 gate380(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate381(.a(s_25), .b(gate49inter3), .O(gate49inter10));
  nor2  gate382(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate383(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate384(.a(gate49inter12), .b(gate49inter1), .O(N314));
xor2 gate50( .a(N276), .b(N277), .O(N315) );

  xor2  gate427(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate428(.a(gate51inter0), .b(s_32), .O(gate51inter1));
  and2  gate429(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate430(.a(s_32), .O(gate51inter3));
  inv1  gate431(.a(s_33), .O(gate51inter4));
  nand2 gate432(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate433(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate434(.a(N278), .O(gate51inter7));
  inv1  gate435(.a(N279), .O(gate51inter8));
  nand2 gate436(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate437(.a(s_33), .b(gate51inter3), .O(gate51inter10));
  nor2  gate438(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate439(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate440(.a(gate51inter12), .b(gate51inter1), .O(N316));
xor2 gate52( .a(N280), .b(N281), .O(N317) );

  xor2  gate287(.a(N283), .b(N282), .O(gate53inter0));
  nand2 gate288(.a(gate53inter0), .b(s_12), .O(gate53inter1));
  and2  gate289(.a(N283), .b(N282), .O(gate53inter2));
  inv1  gate290(.a(s_12), .O(gate53inter3));
  inv1  gate291(.a(s_13), .O(gate53inter4));
  nand2 gate292(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate293(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate294(.a(N282), .O(gate53inter7));
  inv1  gate295(.a(N283), .O(gate53inter8));
  nand2 gate296(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate297(.a(s_13), .b(gate53inter3), .O(gate53inter10));
  nor2  gate298(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate299(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate300(.a(gate53inter12), .b(gate53inter1), .O(N318));
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );

  xor2  gate455(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate456(.a(gate58inter0), .b(s_36), .O(gate58inter1));
  and2  gate457(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate458(.a(s_36), .O(gate58inter3));
  inv1  gate459(.a(s_37), .O(gate58inter4));
  nand2 gate460(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate461(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate462(.a(N296), .O(gate58inter7));
  inv1  gate463(.a(N299), .O(gate58inter8));
  nand2 gate464(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate465(.a(s_37), .b(gate58inter3), .O(gate58inter10));
  nor2  gate466(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate467(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate468(.a(gate58inter12), .b(gate58inter1), .O(N339));
xor2 gate59( .a(N290), .b(N296), .O(N340) );

  xor2  gate483(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate484(.a(gate60inter0), .b(s_40), .O(gate60inter1));
  and2  gate485(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate486(.a(s_40), .O(gate60inter3));
  inv1  gate487(.a(s_41), .O(gate60inter4));
  nand2 gate488(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate489(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate490(.a(N293), .O(gate60inter7));
  inv1  gate491(.a(N299), .O(gate60inter8));
  nand2 gate492(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate493(.a(s_41), .b(gate60inter3), .O(gate60inter10));
  nor2  gate494(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate495(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate496(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );

  xor2  gate245(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate246(.a(gate77inter0), .b(s_6), .O(gate77inter1));
  and2  gate247(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate248(.a(s_6), .O(gate77inter3));
  inv1  gate249(.a(s_7), .O(gate77inter4));
  nand2 gate250(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate251(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate252(.a(N318), .O(gate77inter7));
  inv1  gate253(.a(N350), .O(gate77inter8));
  nand2 gate254(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate255(.a(s_7), .b(gate77inter3), .O(gate77inter10));
  nor2  gate256(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate257(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate258(.a(gate77inter12), .b(gate77inter1), .O(N406));
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate203(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate204(.a(gate172inter0), .b(s_0), .O(gate172inter1));
  and2  gate205(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate206(.a(s_0), .O(gate172inter3));
  inv1  gate207(.a(s_1), .O(gate172inter4));
  nand2 gate208(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate209(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate210(.a(N5), .O(gate172inter7));
  inv1  gate211(.a(N693), .O(gate172inter8));
  nand2 gate212(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate213(.a(s_1), .b(gate172inter3), .O(gate172inter10));
  nor2  gate214(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate215(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate216(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate217(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate218(.a(gate177inter0), .b(s_2), .O(gate177inter1));
  and2  gate219(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate220(.a(s_2), .O(gate177inter3));
  inv1  gate221(.a(s_3), .O(gate177inter4));
  nand2 gate222(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate223(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate224(.a(N25), .O(gate177inter7));
  inv1  gate225(.a(N698), .O(gate177inter8));
  nand2 gate226(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate227(.a(s_3), .b(gate177inter3), .O(gate177inter10));
  nor2  gate228(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate229(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate230(.a(gate177inter12), .b(gate177inter1), .O(N730));
xor2 gate178( .a(N29), .b(N699), .O(N731) );

  xor2  gate343(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate344(.a(gate179inter0), .b(s_20), .O(gate179inter1));
  and2  gate345(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate346(.a(s_20), .O(gate179inter3));
  inv1  gate347(.a(s_21), .O(gate179inter4));
  nand2 gate348(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate349(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate350(.a(N33), .O(gate179inter7));
  inv1  gate351(.a(N700), .O(gate179inter8));
  nand2 gate352(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate353(.a(s_21), .b(gate179inter3), .O(gate179inter10));
  nor2  gate354(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate355(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate356(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );

  xor2  gate385(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate386(.a(gate182inter0), .b(s_26), .O(gate182inter1));
  and2  gate387(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate388(.a(s_26), .O(gate182inter3));
  inv1  gate389(.a(s_27), .O(gate182inter4));
  nand2 gate390(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate391(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate392(.a(N45), .O(gate182inter7));
  inv1  gate393(.a(N703), .O(gate182inter8));
  nand2 gate394(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate395(.a(s_27), .b(gate182inter3), .O(gate182inter10));
  nor2  gate396(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate397(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate398(.a(gate182inter12), .b(gate182inter1), .O(N735));
xor2 gate183( .a(N49), .b(N704), .O(N736) );

  xor2  gate259(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate260(.a(gate184inter0), .b(s_8), .O(gate184inter1));
  and2  gate261(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate262(.a(s_8), .O(gate184inter3));
  inv1  gate263(.a(s_9), .O(gate184inter4));
  nand2 gate264(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate265(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate266(.a(N53), .O(gate184inter7));
  inv1  gate267(.a(N705), .O(gate184inter8));
  nand2 gate268(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate269(.a(s_9), .b(gate184inter3), .O(gate184inter10));
  nor2  gate270(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate271(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate272(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );

  xor2  gate357(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate358(.a(gate192inter0), .b(s_22), .O(gate192inter1));
  and2  gate359(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate360(.a(s_22), .O(gate192inter3));
  inv1  gate361(.a(s_23), .O(gate192inter4));
  nand2 gate362(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate363(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate364(.a(N85), .O(gate192inter7));
  inv1  gate365(.a(N713), .O(gate192inter8));
  nand2 gate366(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate367(.a(s_23), .b(gate192inter3), .O(gate192inter10));
  nor2  gate368(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate369(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate370(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );

  xor2  gate231(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate232(.a(gate194inter0), .b(s_4), .O(gate194inter1));
  and2  gate233(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate234(.a(s_4), .O(gate194inter3));
  inv1  gate235(.a(s_5), .O(gate194inter4));
  nand2 gate236(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate237(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate238(.a(N93), .O(gate194inter7));
  inv1  gate239(.a(N715), .O(gate194inter8));
  nand2 gate240(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate241(.a(s_5), .b(gate194inter3), .O(gate194inter10));
  nor2  gate242(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate243(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate244(.a(gate194inter12), .b(gate194inter1), .O(N747));
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule