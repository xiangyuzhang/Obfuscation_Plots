module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1695(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1696(.a(gate9inter0), .b(s_164), .O(gate9inter1));
  and2  gate1697(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1698(.a(s_164), .O(gate9inter3));
  inv1  gate1699(.a(s_165), .O(gate9inter4));
  nand2 gate1700(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1701(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1702(.a(G1), .O(gate9inter7));
  inv1  gate1703(.a(G2), .O(gate9inter8));
  nand2 gate1704(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1705(.a(s_165), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1706(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1707(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1708(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1807(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1808(.a(gate11inter0), .b(s_180), .O(gate11inter1));
  and2  gate1809(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1810(.a(s_180), .O(gate11inter3));
  inv1  gate1811(.a(s_181), .O(gate11inter4));
  nand2 gate1812(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1813(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1814(.a(G5), .O(gate11inter7));
  inv1  gate1815(.a(G6), .O(gate11inter8));
  nand2 gate1816(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1817(.a(s_181), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1818(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1819(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1820(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2703(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2704(.a(gate19inter0), .b(s_308), .O(gate19inter1));
  and2  gate2705(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2706(.a(s_308), .O(gate19inter3));
  inv1  gate2707(.a(s_309), .O(gate19inter4));
  nand2 gate2708(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2709(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2710(.a(G21), .O(gate19inter7));
  inv1  gate2711(.a(G22), .O(gate19inter8));
  nand2 gate2712(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2713(.a(s_309), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2714(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2715(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2716(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2045(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2046(.a(gate20inter0), .b(s_214), .O(gate20inter1));
  and2  gate2047(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2048(.a(s_214), .O(gate20inter3));
  inv1  gate2049(.a(s_215), .O(gate20inter4));
  nand2 gate2050(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2051(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2052(.a(G23), .O(gate20inter7));
  inv1  gate2053(.a(G24), .O(gate20inter8));
  nand2 gate2054(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2055(.a(s_215), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2056(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2057(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2058(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2353(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2354(.a(gate24inter0), .b(s_258), .O(gate24inter1));
  and2  gate2355(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2356(.a(s_258), .O(gate24inter3));
  inv1  gate2357(.a(s_259), .O(gate24inter4));
  nand2 gate2358(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2359(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2360(.a(G31), .O(gate24inter7));
  inv1  gate2361(.a(G32), .O(gate24inter8));
  nand2 gate2362(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2363(.a(s_259), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2364(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2365(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2366(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate547(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate548(.a(gate27inter0), .b(s_0), .O(gate27inter1));
  and2  gate549(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate550(.a(s_0), .O(gate27inter3));
  inv1  gate551(.a(s_1), .O(gate27inter4));
  nand2 gate552(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate553(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate554(.a(G2), .O(gate27inter7));
  inv1  gate555(.a(G6), .O(gate27inter8));
  nand2 gate556(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate557(.a(s_1), .b(gate27inter3), .O(gate27inter10));
  nor2  gate558(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate559(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate560(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1163(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1164(.a(gate29inter0), .b(s_88), .O(gate29inter1));
  and2  gate1165(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1166(.a(s_88), .O(gate29inter3));
  inv1  gate1167(.a(s_89), .O(gate29inter4));
  nand2 gate1168(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1169(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1170(.a(G3), .O(gate29inter7));
  inv1  gate1171(.a(G7), .O(gate29inter8));
  nand2 gate1172(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1173(.a(s_89), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1174(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1175(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1176(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2143(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2144(.a(gate30inter0), .b(s_228), .O(gate30inter1));
  and2  gate2145(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2146(.a(s_228), .O(gate30inter3));
  inv1  gate2147(.a(s_229), .O(gate30inter4));
  nand2 gate2148(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2149(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2150(.a(G11), .O(gate30inter7));
  inv1  gate2151(.a(G15), .O(gate30inter8));
  nand2 gate2152(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2153(.a(s_229), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2154(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2155(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2156(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1891(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1892(.a(gate31inter0), .b(s_192), .O(gate31inter1));
  and2  gate1893(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1894(.a(s_192), .O(gate31inter3));
  inv1  gate1895(.a(s_193), .O(gate31inter4));
  nand2 gate1896(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1897(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1898(.a(G4), .O(gate31inter7));
  inv1  gate1899(.a(G8), .O(gate31inter8));
  nand2 gate1900(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1901(.a(s_193), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1902(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1903(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1904(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1975(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1976(.a(gate33inter0), .b(s_204), .O(gate33inter1));
  and2  gate1977(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1978(.a(s_204), .O(gate33inter3));
  inv1  gate1979(.a(s_205), .O(gate33inter4));
  nand2 gate1980(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1981(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1982(.a(G17), .O(gate33inter7));
  inv1  gate1983(.a(G21), .O(gate33inter8));
  nand2 gate1984(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1985(.a(s_205), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1986(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1987(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1988(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2843(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2844(.a(gate35inter0), .b(s_328), .O(gate35inter1));
  and2  gate2845(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2846(.a(s_328), .O(gate35inter3));
  inv1  gate2847(.a(s_329), .O(gate35inter4));
  nand2 gate2848(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2849(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2850(.a(G18), .O(gate35inter7));
  inv1  gate2851(.a(G22), .O(gate35inter8));
  nand2 gate2852(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2853(.a(s_329), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2854(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2855(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2856(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2255(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2256(.a(gate37inter0), .b(s_244), .O(gate37inter1));
  and2  gate2257(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2258(.a(s_244), .O(gate37inter3));
  inv1  gate2259(.a(s_245), .O(gate37inter4));
  nand2 gate2260(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2261(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2262(.a(G19), .O(gate37inter7));
  inv1  gate2263(.a(G23), .O(gate37inter8));
  nand2 gate2264(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2265(.a(s_245), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2266(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2267(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2268(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1527(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1528(.a(gate49inter0), .b(s_140), .O(gate49inter1));
  and2  gate1529(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1530(.a(s_140), .O(gate49inter3));
  inv1  gate1531(.a(s_141), .O(gate49inter4));
  nand2 gate1532(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1533(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1534(.a(G9), .O(gate49inter7));
  inv1  gate1535(.a(G278), .O(gate49inter8));
  nand2 gate1536(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1537(.a(s_141), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1538(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1539(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1540(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1415(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1416(.a(gate50inter0), .b(s_124), .O(gate50inter1));
  and2  gate1417(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1418(.a(s_124), .O(gate50inter3));
  inv1  gate1419(.a(s_125), .O(gate50inter4));
  nand2 gate1420(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1421(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1422(.a(G10), .O(gate50inter7));
  inv1  gate1423(.a(G278), .O(gate50inter8));
  nand2 gate1424(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1425(.a(s_125), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1426(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1427(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1428(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate603(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate604(.a(gate53inter0), .b(s_8), .O(gate53inter1));
  and2  gate605(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate606(.a(s_8), .O(gate53inter3));
  inv1  gate607(.a(s_9), .O(gate53inter4));
  nand2 gate608(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate609(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate610(.a(G13), .O(gate53inter7));
  inv1  gate611(.a(G284), .O(gate53inter8));
  nand2 gate612(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate613(.a(s_9), .b(gate53inter3), .O(gate53inter10));
  nor2  gate614(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate615(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate616(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1597(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1598(.a(gate58inter0), .b(s_150), .O(gate58inter1));
  and2  gate1599(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1600(.a(s_150), .O(gate58inter3));
  inv1  gate1601(.a(s_151), .O(gate58inter4));
  nand2 gate1602(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1603(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1604(.a(G18), .O(gate58inter7));
  inv1  gate1605(.a(G290), .O(gate58inter8));
  nand2 gate1606(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1607(.a(s_151), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1608(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1609(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1610(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1919(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1920(.a(gate60inter0), .b(s_196), .O(gate60inter1));
  and2  gate1921(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1922(.a(s_196), .O(gate60inter3));
  inv1  gate1923(.a(s_197), .O(gate60inter4));
  nand2 gate1924(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1925(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1926(.a(G20), .O(gate60inter7));
  inv1  gate1927(.a(G293), .O(gate60inter8));
  nand2 gate1928(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1929(.a(s_197), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1930(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1931(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1932(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate925(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate926(.a(gate63inter0), .b(s_54), .O(gate63inter1));
  and2  gate927(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate928(.a(s_54), .O(gate63inter3));
  inv1  gate929(.a(s_55), .O(gate63inter4));
  nand2 gate930(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate931(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate932(.a(G23), .O(gate63inter7));
  inv1  gate933(.a(G299), .O(gate63inter8));
  nand2 gate934(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate935(.a(s_55), .b(gate63inter3), .O(gate63inter10));
  nor2  gate936(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate937(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate938(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2661(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2662(.a(gate64inter0), .b(s_302), .O(gate64inter1));
  and2  gate2663(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2664(.a(s_302), .O(gate64inter3));
  inv1  gate2665(.a(s_303), .O(gate64inter4));
  nand2 gate2666(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2667(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2668(.a(G24), .O(gate64inter7));
  inv1  gate2669(.a(G299), .O(gate64inter8));
  nand2 gate2670(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2671(.a(s_303), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2672(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2673(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2674(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1401(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1402(.a(gate65inter0), .b(s_122), .O(gate65inter1));
  and2  gate1403(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1404(.a(s_122), .O(gate65inter3));
  inv1  gate1405(.a(s_123), .O(gate65inter4));
  nand2 gate1406(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1407(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1408(.a(G25), .O(gate65inter7));
  inv1  gate1409(.a(G302), .O(gate65inter8));
  nand2 gate1410(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1411(.a(s_123), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1412(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1413(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1414(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1443(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1444(.a(gate67inter0), .b(s_128), .O(gate67inter1));
  and2  gate1445(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1446(.a(s_128), .O(gate67inter3));
  inv1  gate1447(.a(s_129), .O(gate67inter4));
  nand2 gate1448(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1449(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1450(.a(G27), .O(gate67inter7));
  inv1  gate1451(.a(G305), .O(gate67inter8));
  nand2 gate1452(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1453(.a(s_129), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1454(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1455(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1456(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2199(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2200(.a(gate72inter0), .b(s_236), .O(gate72inter1));
  and2  gate2201(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2202(.a(s_236), .O(gate72inter3));
  inv1  gate2203(.a(s_237), .O(gate72inter4));
  nand2 gate2204(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2205(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2206(.a(G32), .O(gate72inter7));
  inv1  gate2207(.a(G311), .O(gate72inter8));
  nand2 gate2208(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2209(.a(s_237), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2210(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2211(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2212(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1849(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1850(.a(gate76inter0), .b(s_186), .O(gate76inter1));
  and2  gate1851(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1852(.a(s_186), .O(gate76inter3));
  inv1  gate1853(.a(s_187), .O(gate76inter4));
  nand2 gate1854(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1855(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1856(.a(G13), .O(gate76inter7));
  inv1  gate1857(.a(G317), .O(gate76inter8));
  nand2 gate1858(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1859(.a(s_187), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1860(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1861(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1862(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2647(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2648(.a(gate81inter0), .b(s_300), .O(gate81inter1));
  and2  gate2649(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2650(.a(s_300), .O(gate81inter3));
  inv1  gate2651(.a(s_301), .O(gate81inter4));
  nand2 gate2652(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2653(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2654(.a(G3), .O(gate81inter7));
  inv1  gate2655(.a(G326), .O(gate81inter8));
  nand2 gate2656(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2657(.a(s_301), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2658(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2659(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2660(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2185(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2186(.a(gate87inter0), .b(s_234), .O(gate87inter1));
  and2  gate2187(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2188(.a(s_234), .O(gate87inter3));
  inv1  gate2189(.a(s_235), .O(gate87inter4));
  nand2 gate2190(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2191(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2192(.a(G12), .O(gate87inter7));
  inv1  gate2193(.a(G335), .O(gate87inter8));
  nand2 gate2194(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2195(.a(s_235), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2196(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2197(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2198(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate617(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate618(.a(gate88inter0), .b(s_10), .O(gate88inter1));
  and2  gate619(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate620(.a(s_10), .O(gate88inter3));
  inv1  gate621(.a(s_11), .O(gate88inter4));
  nand2 gate622(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate623(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate624(.a(G16), .O(gate88inter7));
  inv1  gate625(.a(G335), .O(gate88inter8));
  nand2 gate626(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate627(.a(s_11), .b(gate88inter3), .O(gate88inter10));
  nor2  gate628(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate629(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate630(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2227(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2228(.a(gate90inter0), .b(s_240), .O(gate90inter1));
  and2  gate2229(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2230(.a(s_240), .O(gate90inter3));
  inv1  gate2231(.a(s_241), .O(gate90inter4));
  nand2 gate2232(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2233(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2234(.a(G21), .O(gate90inter7));
  inv1  gate2235(.a(G338), .O(gate90inter8));
  nand2 gate2236(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2237(.a(s_241), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2238(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2239(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2240(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate869(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate870(.a(gate91inter0), .b(s_46), .O(gate91inter1));
  and2  gate871(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate872(.a(s_46), .O(gate91inter3));
  inv1  gate873(.a(s_47), .O(gate91inter4));
  nand2 gate874(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate875(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate876(.a(G25), .O(gate91inter7));
  inv1  gate877(.a(G341), .O(gate91inter8));
  nand2 gate878(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate879(.a(s_47), .b(gate91inter3), .O(gate91inter10));
  nor2  gate880(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate881(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate882(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1905(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1906(.a(gate94inter0), .b(s_194), .O(gate94inter1));
  and2  gate1907(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1908(.a(s_194), .O(gate94inter3));
  inv1  gate1909(.a(s_195), .O(gate94inter4));
  nand2 gate1910(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1911(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1912(.a(G22), .O(gate94inter7));
  inv1  gate1913(.a(G344), .O(gate94inter8));
  nand2 gate1914(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1915(.a(s_195), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1916(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1917(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1918(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate883(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate884(.a(gate95inter0), .b(s_48), .O(gate95inter1));
  and2  gate885(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate886(.a(s_48), .O(gate95inter3));
  inv1  gate887(.a(s_49), .O(gate95inter4));
  nand2 gate888(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate889(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate890(.a(G26), .O(gate95inter7));
  inv1  gate891(.a(G347), .O(gate95inter8));
  nand2 gate892(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate893(.a(s_49), .b(gate95inter3), .O(gate95inter10));
  nor2  gate894(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate895(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate896(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1779(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1780(.a(gate101inter0), .b(s_176), .O(gate101inter1));
  and2  gate1781(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1782(.a(s_176), .O(gate101inter3));
  inv1  gate1783(.a(s_177), .O(gate101inter4));
  nand2 gate1784(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1785(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1786(.a(G20), .O(gate101inter7));
  inv1  gate1787(.a(G356), .O(gate101inter8));
  nand2 gate1788(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1789(.a(s_177), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1790(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1791(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1792(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1947(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1948(.a(gate104inter0), .b(s_200), .O(gate104inter1));
  and2  gate1949(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1950(.a(s_200), .O(gate104inter3));
  inv1  gate1951(.a(s_201), .O(gate104inter4));
  nand2 gate1952(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1953(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1954(.a(G32), .O(gate104inter7));
  inv1  gate1955(.a(G359), .O(gate104inter8));
  nand2 gate1956(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1957(.a(s_201), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1958(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1959(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1960(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate953(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate954(.a(gate105inter0), .b(s_58), .O(gate105inter1));
  and2  gate955(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate956(.a(s_58), .O(gate105inter3));
  inv1  gate957(.a(s_59), .O(gate105inter4));
  nand2 gate958(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate959(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate960(.a(G362), .O(gate105inter7));
  inv1  gate961(.a(G363), .O(gate105inter8));
  nand2 gate962(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate963(.a(s_59), .b(gate105inter3), .O(gate105inter10));
  nor2  gate964(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate965(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate966(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1989(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1990(.a(gate107inter0), .b(s_206), .O(gate107inter1));
  and2  gate1991(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1992(.a(s_206), .O(gate107inter3));
  inv1  gate1993(.a(s_207), .O(gate107inter4));
  nand2 gate1994(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1995(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1996(.a(G366), .O(gate107inter7));
  inv1  gate1997(.a(G367), .O(gate107inter8));
  nand2 gate1998(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1999(.a(s_207), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2000(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2001(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2002(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1373(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1374(.a(gate111inter0), .b(s_118), .O(gate111inter1));
  and2  gate1375(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1376(.a(s_118), .O(gate111inter3));
  inv1  gate1377(.a(s_119), .O(gate111inter4));
  nand2 gate1378(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1379(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1380(.a(G374), .O(gate111inter7));
  inv1  gate1381(.a(G375), .O(gate111inter8));
  nand2 gate1382(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1383(.a(s_119), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1384(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1385(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1386(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate2283(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2284(.a(gate113inter0), .b(s_248), .O(gate113inter1));
  and2  gate2285(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2286(.a(s_248), .O(gate113inter3));
  inv1  gate2287(.a(s_249), .O(gate113inter4));
  nand2 gate2288(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2289(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2290(.a(G378), .O(gate113inter7));
  inv1  gate2291(.a(G379), .O(gate113inter8));
  nand2 gate2292(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2293(.a(s_249), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2294(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2295(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2296(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1023(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1024(.a(gate117inter0), .b(s_68), .O(gate117inter1));
  and2  gate1025(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1026(.a(s_68), .O(gate117inter3));
  inv1  gate1027(.a(s_69), .O(gate117inter4));
  nand2 gate1028(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1029(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1030(.a(G386), .O(gate117inter7));
  inv1  gate1031(.a(G387), .O(gate117inter8));
  nand2 gate1032(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1033(.a(s_69), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1034(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1035(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1036(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1317(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1318(.a(gate119inter0), .b(s_110), .O(gate119inter1));
  and2  gate1319(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1320(.a(s_110), .O(gate119inter3));
  inv1  gate1321(.a(s_111), .O(gate119inter4));
  nand2 gate1322(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1323(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1324(.a(G390), .O(gate119inter7));
  inv1  gate1325(.a(G391), .O(gate119inter8));
  nand2 gate1326(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1327(.a(s_111), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1328(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1329(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1330(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1387(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1388(.a(gate122inter0), .b(s_120), .O(gate122inter1));
  and2  gate1389(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1390(.a(s_120), .O(gate122inter3));
  inv1  gate1391(.a(s_121), .O(gate122inter4));
  nand2 gate1392(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1393(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1394(.a(G396), .O(gate122inter7));
  inv1  gate1395(.a(G397), .O(gate122inter8));
  nand2 gate1396(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1397(.a(s_121), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1398(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1399(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1400(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate2465(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2466(.a(gate123inter0), .b(s_274), .O(gate123inter1));
  and2  gate2467(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2468(.a(s_274), .O(gate123inter3));
  inv1  gate2469(.a(s_275), .O(gate123inter4));
  nand2 gate2470(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2471(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2472(.a(G398), .O(gate123inter7));
  inv1  gate2473(.a(G399), .O(gate123inter8));
  nand2 gate2474(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2475(.a(s_275), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2476(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2477(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2478(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate2059(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2060(.a(gate124inter0), .b(s_216), .O(gate124inter1));
  and2  gate2061(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2062(.a(s_216), .O(gate124inter3));
  inv1  gate2063(.a(s_217), .O(gate124inter4));
  nand2 gate2064(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2065(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2066(.a(G400), .O(gate124inter7));
  inv1  gate2067(.a(G401), .O(gate124inter8));
  nand2 gate2068(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2069(.a(s_217), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2070(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2071(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2072(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate2409(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2410(.a(gate125inter0), .b(s_266), .O(gate125inter1));
  and2  gate2411(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2412(.a(s_266), .O(gate125inter3));
  inv1  gate2413(.a(s_267), .O(gate125inter4));
  nand2 gate2414(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2415(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2416(.a(G402), .O(gate125inter7));
  inv1  gate2417(.a(G403), .O(gate125inter8));
  nand2 gate2418(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2419(.a(s_267), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2420(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2421(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2422(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1233(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1234(.a(gate134inter0), .b(s_98), .O(gate134inter1));
  and2  gate1235(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1236(.a(s_98), .O(gate134inter3));
  inv1  gate1237(.a(s_99), .O(gate134inter4));
  nand2 gate1238(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1239(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1240(.a(G420), .O(gate134inter7));
  inv1  gate1241(.a(G421), .O(gate134inter8));
  nand2 gate1242(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1243(.a(s_99), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1244(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1245(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1246(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate1653(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1654(.a(gate135inter0), .b(s_158), .O(gate135inter1));
  and2  gate1655(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1656(.a(s_158), .O(gate135inter3));
  inv1  gate1657(.a(s_159), .O(gate135inter4));
  nand2 gate1658(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1659(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1660(.a(G422), .O(gate135inter7));
  inv1  gate1661(.a(G423), .O(gate135inter8));
  nand2 gate1662(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1663(.a(s_159), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1664(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1665(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1666(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1793(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1794(.a(gate141inter0), .b(s_178), .O(gate141inter1));
  and2  gate1795(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1796(.a(s_178), .O(gate141inter3));
  inv1  gate1797(.a(s_179), .O(gate141inter4));
  nand2 gate1798(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1799(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1800(.a(G450), .O(gate141inter7));
  inv1  gate1801(.a(G453), .O(gate141inter8));
  nand2 gate1802(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1803(.a(s_179), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1804(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1805(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1806(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1961(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1962(.a(gate145inter0), .b(s_202), .O(gate145inter1));
  and2  gate1963(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1964(.a(s_202), .O(gate145inter3));
  inv1  gate1965(.a(s_203), .O(gate145inter4));
  nand2 gate1966(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1967(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1968(.a(G474), .O(gate145inter7));
  inv1  gate1969(.a(G477), .O(gate145inter8));
  nand2 gate1970(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1971(.a(s_203), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1972(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1973(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1974(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1639(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1640(.a(gate153inter0), .b(s_156), .O(gate153inter1));
  and2  gate1641(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1642(.a(s_156), .O(gate153inter3));
  inv1  gate1643(.a(s_157), .O(gate153inter4));
  nand2 gate1644(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1645(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1646(.a(G426), .O(gate153inter7));
  inv1  gate1647(.a(G522), .O(gate153inter8));
  nand2 gate1648(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1649(.a(s_157), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1650(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1651(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1652(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate701(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate702(.a(gate156inter0), .b(s_22), .O(gate156inter1));
  and2  gate703(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate704(.a(s_22), .O(gate156inter3));
  inv1  gate705(.a(s_23), .O(gate156inter4));
  nand2 gate706(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate707(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate708(.a(G435), .O(gate156inter7));
  inv1  gate709(.a(G525), .O(gate156inter8));
  nand2 gate710(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate711(.a(s_23), .b(gate156inter3), .O(gate156inter10));
  nor2  gate712(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate713(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate714(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate589(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate590(.a(gate159inter0), .b(s_6), .O(gate159inter1));
  and2  gate591(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate592(.a(s_6), .O(gate159inter3));
  inv1  gate593(.a(s_7), .O(gate159inter4));
  nand2 gate594(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate595(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate596(.a(G444), .O(gate159inter7));
  inv1  gate597(.a(G531), .O(gate159inter8));
  nand2 gate598(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate599(.a(s_7), .b(gate159inter3), .O(gate159inter10));
  nor2  gate600(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate601(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate602(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2395(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2396(.a(gate160inter0), .b(s_264), .O(gate160inter1));
  and2  gate2397(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2398(.a(s_264), .O(gate160inter3));
  inv1  gate2399(.a(s_265), .O(gate160inter4));
  nand2 gate2400(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2401(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2402(.a(G447), .O(gate160inter7));
  inv1  gate2403(.a(G531), .O(gate160inter8));
  nand2 gate2404(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2405(.a(s_265), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2406(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2407(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2408(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1121(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1122(.a(gate161inter0), .b(s_82), .O(gate161inter1));
  and2  gate1123(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1124(.a(s_82), .O(gate161inter3));
  inv1  gate1125(.a(s_83), .O(gate161inter4));
  nand2 gate1126(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1127(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1128(.a(G450), .O(gate161inter7));
  inv1  gate1129(.a(G534), .O(gate161inter8));
  nand2 gate1130(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1131(.a(s_83), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1132(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1133(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1134(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1135(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1136(.a(gate162inter0), .b(s_84), .O(gate162inter1));
  and2  gate1137(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1138(.a(s_84), .O(gate162inter3));
  inv1  gate1139(.a(s_85), .O(gate162inter4));
  nand2 gate1140(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1141(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1142(.a(G453), .O(gate162inter7));
  inv1  gate1143(.a(G534), .O(gate162inter8));
  nand2 gate1144(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1145(.a(s_85), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1146(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1147(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1148(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2017(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2018(.a(gate171inter0), .b(s_210), .O(gate171inter1));
  and2  gate2019(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2020(.a(s_210), .O(gate171inter3));
  inv1  gate2021(.a(s_211), .O(gate171inter4));
  nand2 gate2022(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2023(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2024(.a(G480), .O(gate171inter7));
  inv1  gate2025(.a(G549), .O(gate171inter8));
  nand2 gate2026(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2027(.a(s_211), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2028(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2029(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2030(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate967(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate968(.a(gate173inter0), .b(s_60), .O(gate173inter1));
  and2  gate969(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate970(.a(s_60), .O(gate173inter3));
  inv1  gate971(.a(s_61), .O(gate173inter4));
  nand2 gate972(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate973(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate974(.a(G486), .O(gate173inter7));
  inv1  gate975(.a(G552), .O(gate173inter8));
  nand2 gate976(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate977(.a(s_61), .b(gate173inter3), .O(gate173inter10));
  nor2  gate978(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate979(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate980(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1709(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1710(.a(gate175inter0), .b(s_166), .O(gate175inter1));
  and2  gate1711(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1712(.a(s_166), .O(gate175inter3));
  inv1  gate1713(.a(s_167), .O(gate175inter4));
  nand2 gate1714(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1715(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1716(.a(G492), .O(gate175inter7));
  inv1  gate1717(.a(G555), .O(gate175inter8));
  nand2 gate1718(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1719(.a(s_167), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1720(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1721(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1722(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1723(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1724(.a(gate177inter0), .b(s_168), .O(gate177inter1));
  and2  gate1725(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1726(.a(s_168), .O(gate177inter3));
  inv1  gate1727(.a(s_169), .O(gate177inter4));
  nand2 gate1728(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1729(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1730(.a(G498), .O(gate177inter7));
  inv1  gate1731(.a(G558), .O(gate177inter8));
  nand2 gate1732(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1733(.a(s_169), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1734(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1735(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1736(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2535(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2536(.a(gate181inter0), .b(s_284), .O(gate181inter1));
  and2  gate2537(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2538(.a(s_284), .O(gate181inter3));
  inv1  gate2539(.a(s_285), .O(gate181inter4));
  nand2 gate2540(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2541(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2542(.a(G510), .O(gate181inter7));
  inv1  gate2543(.a(G564), .O(gate181inter8));
  nand2 gate2544(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2545(.a(s_285), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2546(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2547(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2548(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1303(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1304(.a(gate184inter0), .b(s_108), .O(gate184inter1));
  and2  gate1305(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1306(.a(s_108), .O(gate184inter3));
  inv1  gate1307(.a(s_109), .O(gate184inter4));
  nand2 gate1308(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1309(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1310(.a(G519), .O(gate184inter7));
  inv1  gate1311(.a(G567), .O(gate184inter8));
  nand2 gate1312(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1313(.a(s_109), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1314(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1315(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1316(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2479(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2480(.a(gate185inter0), .b(s_276), .O(gate185inter1));
  and2  gate2481(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2482(.a(s_276), .O(gate185inter3));
  inv1  gate2483(.a(s_277), .O(gate185inter4));
  nand2 gate2484(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2485(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2486(.a(G570), .O(gate185inter7));
  inv1  gate2487(.a(G571), .O(gate185inter8));
  nand2 gate2488(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2489(.a(s_277), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2490(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2491(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2492(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate995(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate996(.a(gate187inter0), .b(s_64), .O(gate187inter1));
  and2  gate997(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate998(.a(s_64), .O(gate187inter3));
  inv1  gate999(.a(s_65), .O(gate187inter4));
  nand2 gate1000(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1001(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1002(.a(G574), .O(gate187inter7));
  inv1  gate1003(.a(G575), .O(gate187inter8));
  nand2 gate1004(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1005(.a(s_65), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1006(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1007(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1008(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1499(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1500(.a(gate189inter0), .b(s_136), .O(gate189inter1));
  and2  gate1501(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1502(.a(s_136), .O(gate189inter3));
  inv1  gate1503(.a(s_137), .O(gate189inter4));
  nand2 gate1504(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1505(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1506(.a(G578), .O(gate189inter7));
  inv1  gate1507(.a(G579), .O(gate189inter8));
  nand2 gate1508(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1509(.a(s_137), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1510(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1511(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1512(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate2563(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2564(.a(gate190inter0), .b(s_288), .O(gate190inter1));
  and2  gate2565(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2566(.a(s_288), .O(gate190inter3));
  inv1  gate2567(.a(s_289), .O(gate190inter4));
  nand2 gate2568(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2569(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2570(.a(G580), .O(gate190inter7));
  inv1  gate2571(.a(G581), .O(gate190inter8));
  nand2 gate2572(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2573(.a(s_289), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2574(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2575(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2576(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2115(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2116(.a(gate192inter0), .b(s_224), .O(gate192inter1));
  and2  gate2117(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2118(.a(s_224), .O(gate192inter3));
  inv1  gate2119(.a(s_225), .O(gate192inter4));
  nand2 gate2120(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2121(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2122(.a(G584), .O(gate192inter7));
  inv1  gate2123(.a(G585), .O(gate192inter8));
  nand2 gate2124(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2125(.a(s_225), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2126(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2127(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2128(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2633(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2634(.a(gate193inter0), .b(s_298), .O(gate193inter1));
  and2  gate2635(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2636(.a(s_298), .O(gate193inter3));
  inv1  gate2637(.a(s_299), .O(gate193inter4));
  nand2 gate2638(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2639(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2640(.a(G586), .O(gate193inter7));
  inv1  gate2641(.a(G587), .O(gate193inter8));
  nand2 gate2642(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2643(.a(s_299), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2644(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2645(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2646(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2451(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2452(.a(gate197inter0), .b(s_272), .O(gate197inter1));
  and2  gate2453(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2454(.a(s_272), .O(gate197inter3));
  inv1  gate2455(.a(s_273), .O(gate197inter4));
  nand2 gate2456(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2457(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2458(.a(G594), .O(gate197inter7));
  inv1  gate2459(.a(G595), .O(gate197inter8));
  nand2 gate2460(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2461(.a(s_273), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2462(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2463(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2464(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate827(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate828(.a(gate201inter0), .b(s_40), .O(gate201inter1));
  and2  gate829(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate830(.a(s_40), .O(gate201inter3));
  inv1  gate831(.a(s_41), .O(gate201inter4));
  nand2 gate832(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate833(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate834(.a(G602), .O(gate201inter7));
  inv1  gate835(.a(G607), .O(gate201inter8));
  nand2 gate836(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate837(.a(s_41), .b(gate201inter3), .O(gate201inter10));
  nor2  gate838(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate839(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate840(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1471(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1472(.a(gate202inter0), .b(s_132), .O(gate202inter1));
  and2  gate1473(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1474(.a(s_132), .O(gate202inter3));
  inv1  gate1475(.a(s_133), .O(gate202inter4));
  nand2 gate1476(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1477(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1478(.a(G612), .O(gate202inter7));
  inv1  gate1479(.a(G617), .O(gate202inter8));
  nand2 gate1480(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1481(.a(s_133), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1482(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1483(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1484(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate757(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate758(.a(gate204inter0), .b(s_30), .O(gate204inter1));
  and2  gate759(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate760(.a(s_30), .O(gate204inter3));
  inv1  gate761(.a(s_31), .O(gate204inter4));
  nand2 gate762(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate763(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate764(.a(G607), .O(gate204inter7));
  inv1  gate765(.a(G617), .O(gate204inter8));
  nand2 gate766(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate767(.a(s_31), .b(gate204inter3), .O(gate204inter10));
  nor2  gate768(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate769(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate770(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate771(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate772(.a(gate207inter0), .b(s_32), .O(gate207inter1));
  and2  gate773(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate774(.a(s_32), .O(gate207inter3));
  inv1  gate775(.a(s_33), .O(gate207inter4));
  nand2 gate776(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate777(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate778(.a(G622), .O(gate207inter7));
  inv1  gate779(.a(G632), .O(gate207inter8));
  nand2 gate780(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate781(.a(s_33), .b(gate207inter3), .O(gate207inter10));
  nor2  gate782(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate783(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate784(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate939(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate940(.a(gate213inter0), .b(s_56), .O(gate213inter1));
  and2  gate941(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate942(.a(s_56), .O(gate213inter3));
  inv1  gate943(.a(s_57), .O(gate213inter4));
  nand2 gate944(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate945(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate946(.a(G602), .O(gate213inter7));
  inv1  gate947(.a(G672), .O(gate213inter8));
  nand2 gate948(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate949(.a(s_57), .b(gate213inter3), .O(gate213inter10));
  nor2  gate950(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate951(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate952(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1751(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1752(.a(gate214inter0), .b(s_172), .O(gate214inter1));
  and2  gate1753(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1754(.a(s_172), .O(gate214inter3));
  inv1  gate1755(.a(s_173), .O(gate214inter4));
  nand2 gate1756(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1757(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1758(.a(G612), .O(gate214inter7));
  inv1  gate1759(.a(G672), .O(gate214inter8));
  nand2 gate1760(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1761(.a(s_173), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1762(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1763(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1764(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1079(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1080(.a(gate216inter0), .b(s_76), .O(gate216inter1));
  and2  gate1081(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1082(.a(s_76), .O(gate216inter3));
  inv1  gate1083(.a(s_77), .O(gate216inter4));
  nand2 gate1084(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1085(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1086(.a(G617), .O(gate216inter7));
  inv1  gate1087(.a(G675), .O(gate216inter8));
  nand2 gate1088(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1089(.a(s_77), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1090(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1091(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1092(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2087(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2088(.a(gate217inter0), .b(s_220), .O(gate217inter1));
  and2  gate2089(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2090(.a(s_220), .O(gate217inter3));
  inv1  gate2091(.a(s_221), .O(gate217inter4));
  nand2 gate2092(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2093(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2094(.a(G622), .O(gate217inter7));
  inv1  gate2095(.a(G678), .O(gate217inter8));
  nand2 gate2096(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2097(.a(s_221), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2098(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2099(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2100(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1457(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1458(.a(gate220inter0), .b(s_130), .O(gate220inter1));
  and2  gate1459(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1460(.a(s_130), .O(gate220inter3));
  inv1  gate1461(.a(s_131), .O(gate220inter4));
  nand2 gate1462(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1463(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1464(.a(G637), .O(gate220inter7));
  inv1  gate1465(.a(G681), .O(gate220inter8));
  nand2 gate1466(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1467(.a(s_131), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1468(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1469(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1470(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate743(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate744(.a(gate222inter0), .b(s_28), .O(gate222inter1));
  and2  gate745(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate746(.a(s_28), .O(gate222inter3));
  inv1  gate747(.a(s_29), .O(gate222inter4));
  nand2 gate748(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate749(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate750(.a(G632), .O(gate222inter7));
  inv1  gate751(.a(G684), .O(gate222inter8));
  nand2 gate752(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate753(.a(s_29), .b(gate222inter3), .O(gate222inter10));
  nor2  gate754(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate755(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate756(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate785(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate786(.a(gate224inter0), .b(s_34), .O(gate224inter1));
  and2  gate787(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate788(.a(s_34), .O(gate224inter3));
  inv1  gate789(.a(s_35), .O(gate224inter4));
  nand2 gate790(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate791(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate792(.a(G637), .O(gate224inter7));
  inv1  gate793(.a(G687), .O(gate224inter8));
  nand2 gate794(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate795(.a(s_35), .b(gate224inter3), .O(gate224inter10));
  nor2  gate796(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate797(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate798(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1191(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1192(.a(gate227inter0), .b(s_92), .O(gate227inter1));
  and2  gate1193(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1194(.a(s_92), .O(gate227inter3));
  inv1  gate1195(.a(s_93), .O(gate227inter4));
  nand2 gate1196(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1197(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1198(.a(G694), .O(gate227inter7));
  inv1  gate1199(.a(G695), .O(gate227inter8));
  nand2 gate1200(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1201(.a(s_93), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1202(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1203(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1204(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate687(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate688(.a(gate231inter0), .b(s_20), .O(gate231inter1));
  and2  gate689(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate690(.a(s_20), .O(gate231inter3));
  inv1  gate691(.a(s_21), .O(gate231inter4));
  nand2 gate692(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate693(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate694(.a(G702), .O(gate231inter7));
  inv1  gate695(.a(G703), .O(gate231inter8));
  nand2 gate696(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate697(.a(s_21), .b(gate231inter3), .O(gate231inter10));
  nor2  gate698(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate699(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate700(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2423(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2424(.a(gate236inter0), .b(s_268), .O(gate236inter1));
  and2  gate2425(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2426(.a(s_268), .O(gate236inter3));
  inv1  gate2427(.a(s_269), .O(gate236inter4));
  nand2 gate2428(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2429(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2430(.a(G251), .O(gate236inter7));
  inv1  gate2431(.a(G727), .O(gate236inter8));
  nand2 gate2432(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2433(.a(s_269), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2434(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2435(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2436(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate2577(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2578(.a(gate237inter0), .b(s_290), .O(gate237inter1));
  and2  gate2579(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2580(.a(s_290), .O(gate237inter3));
  inv1  gate2581(.a(s_291), .O(gate237inter4));
  nand2 gate2582(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2583(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2584(.a(G254), .O(gate237inter7));
  inv1  gate2585(.a(G706), .O(gate237inter8));
  nand2 gate2586(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2587(.a(s_291), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2588(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2589(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2590(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2731(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2732(.a(gate241inter0), .b(s_312), .O(gate241inter1));
  and2  gate2733(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2734(.a(s_312), .O(gate241inter3));
  inv1  gate2735(.a(s_313), .O(gate241inter4));
  nand2 gate2736(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2737(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2738(.a(G242), .O(gate241inter7));
  inv1  gate2739(.a(G730), .O(gate241inter8));
  nand2 gate2740(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2741(.a(s_313), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2742(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2743(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2744(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1331(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1332(.a(gate243inter0), .b(s_112), .O(gate243inter1));
  and2  gate1333(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1334(.a(s_112), .O(gate243inter3));
  inv1  gate1335(.a(s_113), .O(gate243inter4));
  nand2 gate1336(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1337(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1338(.a(G245), .O(gate243inter7));
  inv1  gate1339(.a(G733), .O(gate243inter8));
  nand2 gate1340(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1341(.a(s_113), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1342(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1343(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1344(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate673(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate674(.a(gate246inter0), .b(s_18), .O(gate246inter1));
  and2  gate675(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate676(.a(s_18), .O(gate246inter3));
  inv1  gate677(.a(s_19), .O(gate246inter4));
  nand2 gate678(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate679(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate680(.a(G724), .O(gate246inter7));
  inv1  gate681(.a(G736), .O(gate246inter8));
  nand2 gate682(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate683(.a(s_19), .b(gate246inter3), .O(gate246inter10));
  nor2  gate684(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate685(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate686(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1737(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1738(.a(gate249inter0), .b(s_170), .O(gate249inter1));
  and2  gate1739(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1740(.a(s_170), .O(gate249inter3));
  inv1  gate1741(.a(s_171), .O(gate249inter4));
  nand2 gate1742(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1743(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1744(.a(G254), .O(gate249inter7));
  inv1  gate1745(.a(G742), .O(gate249inter8));
  nand2 gate1746(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1747(.a(s_171), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1748(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1749(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1750(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1611(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1612(.a(gate252inter0), .b(s_152), .O(gate252inter1));
  and2  gate1613(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1614(.a(s_152), .O(gate252inter3));
  inv1  gate1615(.a(s_153), .O(gate252inter4));
  nand2 gate1616(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1617(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1618(.a(G709), .O(gate252inter7));
  inv1  gate1619(.a(G745), .O(gate252inter8));
  nand2 gate1620(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1621(.a(s_153), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1622(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1623(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1624(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2297(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2298(.a(gate254inter0), .b(s_250), .O(gate254inter1));
  and2  gate2299(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2300(.a(s_250), .O(gate254inter3));
  inv1  gate2301(.a(s_251), .O(gate254inter4));
  nand2 gate2302(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2303(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2304(.a(G712), .O(gate254inter7));
  inv1  gate2305(.a(G748), .O(gate254inter8));
  nand2 gate2306(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2307(.a(s_251), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2308(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2309(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2310(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1261(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1262(.a(gate258inter0), .b(s_102), .O(gate258inter1));
  and2  gate1263(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1264(.a(s_102), .O(gate258inter3));
  inv1  gate1265(.a(s_103), .O(gate258inter4));
  nand2 gate1266(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1267(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1268(.a(G756), .O(gate258inter7));
  inv1  gate1269(.a(G757), .O(gate258inter8));
  nand2 gate1270(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1271(.a(s_103), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1272(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1273(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1274(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate841(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate842(.a(gate259inter0), .b(s_42), .O(gate259inter1));
  and2  gate843(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate844(.a(s_42), .O(gate259inter3));
  inv1  gate845(.a(s_43), .O(gate259inter4));
  nand2 gate846(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate847(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate848(.a(G758), .O(gate259inter7));
  inv1  gate849(.a(G759), .O(gate259inter8));
  nand2 gate850(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate851(.a(s_43), .b(gate259inter3), .O(gate259inter10));
  nor2  gate852(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate853(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate854(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate2241(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2242(.a(gate260inter0), .b(s_242), .O(gate260inter1));
  and2  gate2243(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2244(.a(s_242), .O(gate260inter3));
  inv1  gate2245(.a(s_243), .O(gate260inter4));
  nand2 gate2246(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2247(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2248(.a(G760), .O(gate260inter7));
  inv1  gate2249(.a(G761), .O(gate260inter8));
  nand2 gate2250(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2251(.a(s_243), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2252(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2253(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2254(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate575(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate576(.a(gate264inter0), .b(s_4), .O(gate264inter1));
  and2  gate577(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate578(.a(s_4), .O(gate264inter3));
  inv1  gate579(.a(s_5), .O(gate264inter4));
  nand2 gate580(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate581(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate582(.a(G768), .O(gate264inter7));
  inv1  gate583(.a(G769), .O(gate264inter8));
  nand2 gate584(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate585(.a(s_5), .b(gate264inter3), .O(gate264inter10));
  nor2  gate586(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate587(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate588(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1275(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1276(.a(gate266inter0), .b(s_104), .O(gate266inter1));
  and2  gate1277(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1278(.a(s_104), .O(gate266inter3));
  inv1  gate1279(.a(s_105), .O(gate266inter4));
  nand2 gate1280(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1281(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1282(.a(G645), .O(gate266inter7));
  inv1  gate1283(.a(G773), .O(gate266inter8));
  nand2 gate1284(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1285(.a(s_105), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1286(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1287(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1288(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2591(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2592(.a(gate267inter0), .b(s_292), .O(gate267inter1));
  and2  gate2593(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2594(.a(s_292), .O(gate267inter3));
  inv1  gate2595(.a(s_293), .O(gate267inter4));
  nand2 gate2596(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2597(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2598(.a(G648), .O(gate267inter7));
  inv1  gate2599(.a(G776), .O(gate267inter8));
  nand2 gate2600(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2601(.a(s_293), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2602(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2603(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2604(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2437(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2438(.a(gate268inter0), .b(s_270), .O(gate268inter1));
  and2  gate2439(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2440(.a(s_270), .O(gate268inter3));
  inv1  gate2441(.a(s_271), .O(gate268inter4));
  nand2 gate2442(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2443(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2444(.a(G651), .O(gate268inter7));
  inv1  gate2445(.a(G779), .O(gate268inter8));
  nand2 gate2446(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2447(.a(s_271), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2448(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2449(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2450(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2675(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2676(.a(gate269inter0), .b(s_304), .O(gate269inter1));
  and2  gate2677(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2678(.a(s_304), .O(gate269inter3));
  inv1  gate2679(.a(s_305), .O(gate269inter4));
  nand2 gate2680(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2681(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2682(.a(G654), .O(gate269inter7));
  inv1  gate2683(.a(G782), .O(gate269inter8));
  nand2 gate2684(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2685(.a(s_305), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2686(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2687(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2688(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1583(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1584(.a(gate271inter0), .b(s_148), .O(gate271inter1));
  and2  gate1585(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1586(.a(s_148), .O(gate271inter3));
  inv1  gate1587(.a(s_149), .O(gate271inter4));
  nand2 gate1588(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1589(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1590(.a(G660), .O(gate271inter7));
  inv1  gate1591(.a(G788), .O(gate271inter8));
  nand2 gate1592(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1593(.a(s_149), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1594(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1595(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1596(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1149(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1150(.a(gate272inter0), .b(s_86), .O(gate272inter1));
  and2  gate1151(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1152(.a(s_86), .O(gate272inter3));
  inv1  gate1153(.a(s_87), .O(gate272inter4));
  nand2 gate1154(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1155(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1156(.a(G663), .O(gate272inter7));
  inv1  gate1157(.a(G791), .O(gate272inter8));
  nand2 gate1158(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1159(.a(s_87), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1160(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1161(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1162(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate855(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate856(.a(gate273inter0), .b(s_44), .O(gate273inter1));
  and2  gate857(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate858(.a(s_44), .O(gate273inter3));
  inv1  gate859(.a(s_45), .O(gate273inter4));
  nand2 gate860(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate861(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate862(.a(G642), .O(gate273inter7));
  inv1  gate863(.a(G794), .O(gate273inter8));
  nand2 gate864(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate865(.a(s_45), .b(gate273inter3), .O(gate273inter10));
  nor2  gate866(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate867(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate868(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2339(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2340(.a(gate275inter0), .b(s_256), .O(gate275inter1));
  and2  gate2341(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2342(.a(s_256), .O(gate275inter3));
  inv1  gate2343(.a(s_257), .O(gate275inter4));
  nand2 gate2344(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2345(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2346(.a(G645), .O(gate275inter7));
  inv1  gate2347(.a(G797), .O(gate275inter8));
  nand2 gate2348(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2349(.a(s_257), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2350(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2351(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2352(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2101(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2102(.a(gate278inter0), .b(s_222), .O(gate278inter1));
  and2  gate2103(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2104(.a(s_222), .O(gate278inter3));
  inv1  gate2105(.a(s_223), .O(gate278inter4));
  nand2 gate2106(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2107(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2108(.a(G776), .O(gate278inter7));
  inv1  gate2109(.a(G800), .O(gate278inter8));
  nand2 gate2110(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2111(.a(s_223), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2112(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2113(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2114(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1569(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1570(.a(gate280inter0), .b(s_146), .O(gate280inter1));
  and2  gate1571(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1572(.a(s_146), .O(gate280inter3));
  inv1  gate1573(.a(s_147), .O(gate280inter4));
  nand2 gate1574(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1575(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1576(.a(G779), .O(gate280inter7));
  inv1  gate1577(.a(G803), .O(gate280inter8));
  nand2 gate1578(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1579(.a(s_147), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1580(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1581(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1582(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1037(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1038(.a(gate281inter0), .b(s_70), .O(gate281inter1));
  and2  gate1039(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1040(.a(s_70), .O(gate281inter3));
  inv1  gate1041(.a(s_71), .O(gate281inter4));
  nand2 gate1042(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1043(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1044(.a(G654), .O(gate281inter7));
  inv1  gate1045(.a(G806), .O(gate281inter8));
  nand2 gate1046(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1047(.a(s_71), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1048(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1049(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1050(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2829(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2830(.a(gate282inter0), .b(s_326), .O(gate282inter1));
  and2  gate2831(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2832(.a(s_326), .O(gate282inter3));
  inv1  gate2833(.a(s_327), .O(gate282inter4));
  nand2 gate2834(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2835(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2836(.a(G782), .O(gate282inter7));
  inv1  gate2837(.a(G806), .O(gate282inter8));
  nand2 gate2838(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2839(.a(s_327), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2840(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2841(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2842(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1093(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1094(.a(gate284inter0), .b(s_78), .O(gate284inter1));
  and2  gate1095(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1096(.a(s_78), .O(gate284inter3));
  inv1  gate1097(.a(s_79), .O(gate284inter4));
  nand2 gate1098(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1099(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1100(.a(G785), .O(gate284inter7));
  inv1  gate1101(.a(G809), .O(gate284inter8));
  nand2 gate1102(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1103(.a(s_79), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1104(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1105(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1106(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2689(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2690(.a(gate287inter0), .b(s_306), .O(gate287inter1));
  and2  gate2691(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2692(.a(s_306), .O(gate287inter3));
  inv1  gate2693(.a(s_307), .O(gate287inter4));
  nand2 gate2694(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2695(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2696(.a(G663), .O(gate287inter7));
  inv1  gate2697(.a(G815), .O(gate287inter8));
  nand2 gate2698(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2699(.a(s_307), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2700(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2701(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2702(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1681(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1682(.a(gate288inter0), .b(s_162), .O(gate288inter1));
  and2  gate1683(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1684(.a(s_162), .O(gate288inter3));
  inv1  gate1685(.a(s_163), .O(gate288inter4));
  nand2 gate1686(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1687(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1688(.a(G791), .O(gate288inter7));
  inv1  gate1689(.a(G815), .O(gate288inter8));
  nand2 gate1690(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1691(.a(s_163), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1692(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1693(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1694(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1177(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1178(.a(gate290inter0), .b(s_90), .O(gate290inter1));
  and2  gate1179(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1180(.a(s_90), .O(gate290inter3));
  inv1  gate1181(.a(s_91), .O(gate290inter4));
  nand2 gate1182(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1183(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1184(.a(G820), .O(gate290inter7));
  inv1  gate1185(.a(G821), .O(gate290inter8));
  nand2 gate1186(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1187(.a(s_91), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1188(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1189(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1190(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1821(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1822(.a(gate293inter0), .b(s_182), .O(gate293inter1));
  and2  gate1823(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1824(.a(s_182), .O(gate293inter3));
  inv1  gate1825(.a(s_183), .O(gate293inter4));
  nand2 gate1826(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1827(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1828(.a(G828), .O(gate293inter7));
  inv1  gate1829(.a(G829), .O(gate293inter8));
  nand2 gate1830(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1831(.a(s_183), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1832(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1833(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1834(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1863(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1864(.a(gate294inter0), .b(s_188), .O(gate294inter1));
  and2  gate1865(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1866(.a(s_188), .O(gate294inter3));
  inv1  gate1867(.a(s_189), .O(gate294inter4));
  nand2 gate1868(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1869(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1870(.a(G832), .O(gate294inter7));
  inv1  gate1871(.a(G833), .O(gate294inter8));
  nand2 gate1872(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1873(.a(s_189), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1874(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1875(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1876(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1765(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1766(.a(gate388inter0), .b(s_174), .O(gate388inter1));
  and2  gate1767(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1768(.a(s_174), .O(gate388inter3));
  inv1  gate1769(.a(s_175), .O(gate388inter4));
  nand2 gate1770(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1771(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1772(.a(G2), .O(gate388inter7));
  inv1  gate1773(.a(G1039), .O(gate388inter8));
  nand2 gate1774(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1775(.a(s_175), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1776(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1777(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1778(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2213(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2214(.a(gate389inter0), .b(s_238), .O(gate389inter1));
  and2  gate2215(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2216(.a(s_238), .O(gate389inter3));
  inv1  gate2217(.a(s_239), .O(gate389inter4));
  nand2 gate2218(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2219(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2220(.a(G3), .O(gate389inter7));
  inv1  gate2221(.a(G1042), .O(gate389inter8));
  nand2 gate2222(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2223(.a(s_239), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2224(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2225(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2226(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2381(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2382(.a(gate396inter0), .b(s_262), .O(gate396inter1));
  and2  gate2383(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2384(.a(s_262), .O(gate396inter3));
  inv1  gate2385(.a(s_263), .O(gate396inter4));
  nand2 gate2386(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2387(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2388(.a(G10), .O(gate396inter7));
  inv1  gate2389(.a(G1063), .O(gate396inter8));
  nand2 gate2390(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2391(.a(s_263), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2392(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2393(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2394(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2605(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2606(.a(gate398inter0), .b(s_294), .O(gate398inter1));
  and2  gate2607(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2608(.a(s_294), .O(gate398inter3));
  inv1  gate2609(.a(s_295), .O(gate398inter4));
  nand2 gate2610(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2611(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2612(.a(G12), .O(gate398inter7));
  inv1  gate2613(.a(G1069), .O(gate398inter8));
  nand2 gate2614(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2615(.a(s_295), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2616(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2617(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2618(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate2367(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2368(.a(gate399inter0), .b(s_260), .O(gate399inter1));
  and2  gate2369(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2370(.a(s_260), .O(gate399inter3));
  inv1  gate2371(.a(s_261), .O(gate399inter4));
  nand2 gate2372(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2373(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2374(.a(G13), .O(gate399inter7));
  inv1  gate2375(.a(G1072), .O(gate399inter8));
  nand2 gate2376(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2377(.a(s_261), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2378(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2379(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2380(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate813(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate814(.a(gate400inter0), .b(s_38), .O(gate400inter1));
  and2  gate815(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate816(.a(s_38), .O(gate400inter3));
  inv1  gate817(.a(s_39), .O(gate400inter4));
  nand2 gate818(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate819(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate820(.a(G14), .O(gate400inter7));
  inv1  gate821(.a(G1075), .O(gate400inter8));
  nand2 gate822(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate823(.a(s_39), .b(gate400inter3), .O(gate400inter10));
  nor2  gate824(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate825(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate826(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1877(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1878(.a(gate403inter0), .b(s_190), .O(gate403inter1));
  and2  gate1879(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1880(.a(s_190), .O(gate403inter3));
  inv1  gate1881(.a(s_191), .O(gate403inter4));
  nand2 gate1882(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1883(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1884(.a(G17), .O(gate403inter7));
  inv1  gate1885(.a(G1084), .O(gate403inter8));
  nand2 gate1886(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1887(.a(s_191), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1888(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1889(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1890(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1247(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1248(.a(gate404inter0), .b(s_100), .O(gate404inter1));
  and2  gate1249(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1250(.a(s_100), .O(gate404inter3));
  inv1  gate1251(.a(s_101), .O(gate404inter4));
  nand2 gate1252(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1253(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1254(.a(G18), .O(gate404inter7));
  inv1  gate1255(.a(G1087), .O(gate404inter8));
  nand2 gate1256(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1257(.a(s_101), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1258(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1259(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1260(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1345(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1346(.a(gate407inter0), .b(s_114), .O(gate407inter1));
  and2  gate1347(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1348(.a(s_114), .O(gate407inter3));
  inv1  gate1349(.a(s_115), .O(gate407inter4));
  nand2 gate1350(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1351(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1352(.a(G21), .O(gate407inter7));
  inv1  gate1353(.a(G1096), .O(gate407inter8));
  nand2 gate1354(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1355(.a(s_115), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1356(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1357(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1358(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate2325(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2326(.a(gate408inter0), .b(s_254), .O(gate408inter1));
  and2  gate2327(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2328(.a(s_254), .O(gate408inter3));
  inv1  gate2329(.a(s_255), .O(gate408inter4));
  nand2 gate2330(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2331(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2332(.a(G22), .O(gate408inter7));
  inv1  gate2333(.a(G1099), .O(gate408inter8));
  nand2 gate2334(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2335(.a(s_255), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2336(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2337(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2338(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate631(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate632(.a(gate409inter0), .b(s_12), .O(gate409inter1));
  and2  gate633(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate634(.a(s_12), .O(gate409inter3));
  inv1  gate635(.a(s_13), .O(gate409inter4));
  nand2 gate636(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate637(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate638(.a(G23), .O(gate409inter7));
  inv1  gate639(.a(G1102), .O(gate409inter8));
  nand2 gate640(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate641(.a(s_13), .b(gate409inter3), .O(gate409inter10));
  nor2  gate642(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate643(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate644(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1835(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1836(.a(gate411inter0), .b(s_184), .O(gate411inter1));
  and2  gate1837(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1838(.a(s_184), .O(gate411inter3));
  inv1  gate1839(.a(s_185), .O(gate411inter4));
  nand2 gate1840(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1841(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1842(.a(G25), .O(gate411inter7));
  inv1  gate1843(.a(G1108), .O(gate411inter8));
  nand2 gate1844(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1845(.a(s_185), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1846(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1847(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1848(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2493(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2494(.a(gate413inter0), .b(s_278), .O(gate413inter1));
  and2  gate2495(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2496(.a(s_278), .O(gate413inter3));
  inv1  gate2497(.a(s_279), .O(gate413inter4));
  nand2 gate2498(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2499(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2500(.a(G27), .O(gate413inter7));
  inv1  gate2501(.a(G1114), .O(gate413inter8));
  nand2 gate2502(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2503(.a(s_279), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2504(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2505(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2506(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1205(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1206(.a(gate418inter0), .b(s_94), .O(gate418inter1));
  and2  gate1207(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1208(.a(s_94), .O(gate418inter3));
  inv1  gate1209(.a(s_95), .O(gate418inter4));
  nand2 gate1210(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1211(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1212(.a(G32), .O(gate418inter7));
  inv1  gate1213(.a(G1129), .O(gate418inter8));
  nand2 gate1214(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1215(.a(s_95), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1216(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1217(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1218(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate981(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate982(.a(gate420inter0), .b(s_62), .O(gate420inter1));
  and2  gate983(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate984(.a(s_62), .O(gate420inter3));
  inv1  gate985(.a(s_63), .O(gate420inter4));
  nand2 gate986(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate987(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate988(.a(G1036), .O(gate420inter7));
  inv1  gate989(.a(G1132), .O(gate420inter8));
  nand2 gate990(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate991(.a(s_63), .b(gate420inter3), .O(gate420inter10));
  nor2  gate992(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate993(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate994(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1667(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1668(.a(gate424inter0), .b(s_160), .O(gate424inter1));
  and2  gate1669(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1670(.a(s_160), .O(gate424inter3));
  inv1  gate1671(.a(s_161), .O(gate424inter4));
  nand2 gate1672(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1673(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1674(.a(G1042), .O(gate424inter7));
  inv1  gate1675(.a(G1138), .O(gate424inter8));
  nand2 gate1676(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1677(.a(s_161), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1678(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1679(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1680(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1289(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1290(.a(gate426inter0), .b(s_106), .O(gate426inter1));
  and2  gate1291(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1292(.a(s_106), .O(gate426inter3));
  inv1  gate1293(.a(s_107), .O(gate426inter4));
  nand2 gate1294(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1295(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1296(.a(G1045), .O(gate426inter7));
  inv1  gate1297(.a(G1141), .O(gate426inter8));
  nand2 gate1298(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1299(.a(s_107), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1300(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1301(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1302(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2269(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2270(.a(gate429inter0), .b(s_246), .O(gate429inter1));
  and2  gate2271(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2272(.a(s_246), .O(gate429inter3));
  inv1  gate2273(.a(s_247), .O(gate429inter4));
  nand2 gate2274(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2275(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2276(.a(G6), .O(gate429inter7));
  inv1  gate2277(.a(G1147), .O(gate429inter8));
  nand2 gate2278(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2279(.a(s_247), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2280(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2281(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2282(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate2157(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2158(.a(gate430inter0), .b(s_230), .O(gate430inter1));
  and2  gate2159(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2160(.a(s_230), .O(gate430inter3));
  inv1  gate2161(.a(s_231), .O(gate430inter4));
  nand2 gate2162(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2163(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2164(.a(G1051), .O(gate430inter7));
  inv1  gate2165(.a(G1147), .O(gate430inter8));
  nand2 gate2166(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2167(.a(s_231), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2168(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2169(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2170(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2031(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2032(.a(gate431inter0), .b(s_212), .O(gate431inter1));
  and2  gate2033(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2034(.a(s_212), .O(gate431inter3));
  inv1  gate2035(.a(s_213), .O(gate431inter4));
  nand2 gate2036(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2037(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2038(.a(G7), .O(gate431inter7));
  inv1  gate2039(.a(G1150), .O(gate431inter8));
  nand2 gate2040(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2041(.a(s_213), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2042(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2043(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2044(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1219(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1220(.a(gate432inter0), .b(s_96), .O(gate432inter1));
  and2  gate1221(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1222(.a(s_96), .O(gate432inter3));
  inv1  gate1223(.a(s_97), .O(gate432inter4));
  nand2 gate1224(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1225(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1226(.a(G1054), .O(gate432inter7));
  inv1  gate1227(.a(G1150), .O(gate432inter8));
  nand2 gate1228(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1229(.a(s_97), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1230(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1231(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1232(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2801(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2802(.a(gate434inter0), .b(s_322), .O(gate434inter1));
  and2  gate2803(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2804(.a(s_322), .O(gate434inter3));
  inv1  gate2805(.a(s_323), .O(gate434inter4));
  nand2 gate2806(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2807(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2808(.a(G1057), .O(gate434inter7));
  inv1  gate2809(.a(G1153), .O(gate434inter8));
  nand2 gate2810(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2811(.a(s_323), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2812(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2813(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2814(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate715(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate716(.a(gate436inter0), .b(s_24), .O(gate436inter1));
  and2  gate717(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate718(.a(s_24), .O(gate436inter3));
  inv1  gate719(.a(s_25), .O(gate436inter4));
  nand2 gate720(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate721(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate722(.a(G1060), .O(gate436inter7));
  inv1  gate723(.a(G1156), .O(gate436inter8));
  nand2 gate724(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate725(.a(s_25), .b(gate436inter3), .O(gate436inter10));
  nor2  gate726(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate727(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate728(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate2311(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2312(.a(gate437inter0), .b(s_252), .O(gate437inter1));
  and2  gate2313(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2314(.a(s_252), .O(gate437inter3));
  inv1  gate2315(.a(s_253), .O(gate437inter4));
  nand2 gate2316(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2317(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2318(.a(G10), .O(gate437inter7));
  inv1  gate2319(.a(G1159), .O(gate437inter8));
  nand2 gate2320(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2321(.a(s_253), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2322(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2323(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2324(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2171(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2172(.a(gate439inter0), .b(s_232), .O(gate439inter1));
  and2  gate2173(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2174(.a(s_232), .O(gate439inter3));
  inv1  gate2175(.a(s_233), .O(gate439inter4));
  nand2 gate2176(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2177(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2178(.a(G11), .O(gate439inter7));
  inv1  gate2179(.a(G1162), .O(gate439inter8));
  nand2 gate2180(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2181(.a(s_233), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2182(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2183(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2184(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2549(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2550(.a(gate442inter0), .b(s_286), .O(gate442inter1));
  and2  gate2551(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2552(.a(s_286), .O(gate442inter3));
  inv1  gate2553(.a(s_287), .O(gate442inter4));
  nand2 gate2554(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2555(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2556(.a(G1069), .O(gate442inter7));
  inv1  gate2557(.a(G1165), .O(gate442inter8));
  nand2 gate2558(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2559(.a(s_287), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2560(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2561(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2562(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1359(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1360(.a(gate444inter0), .b(s_116), .O(gate444inter1));
  and2  gate1361(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1362(.a(s_116), .O(gate444inter3));
  inv1  gate1363(.a(s_117), .O(gate444inter4));
  nand2 gate1364(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1365(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1366(.a(G1072), .O(gate444inter7));
  inv1  gate1367(.a(G1168), .O(gate444inter8));
  nand2 gate1368(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1369(.a(s_117), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1370(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1371(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1372(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate897(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate898(.a(gate448inter0), .b(s_50), .O(gate448inter1));
  and2  gate899(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate900(.a(s_50), .O(gate448inter3));
  inv1  gate901(.a(s_51), .O(gate448inter4));
  nand2 gate902(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate903(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate904(.a(G1078), .O(gate448inter7));
  inv1  gate905(.a(G1174), .O(gate448inter8));
  nand2 gate906(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate907(.a(s_51), .b(gate448inter3), .O(gate448inter10));
  nor2  gate908(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate909(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate910(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1513(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1514(.a(gate449inter0), .b(s_138), .O(gate449inter1));
  and2  gate1515(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1516(.a(s_138), .O(gate449inter3));
  inv1  gate1517(.a(s_139), .O(gate449inter4));
  nand2 gate1518(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1519(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1520(.a(G16), .O(gate449inter7));
  inv1  gate1521(.a(G1177), .O(gate449inter8));
  nand2 gate1522(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1523(.a(s_139), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1524(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1525(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1526(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate2773(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2774(.a(gate450inter0), .b(s_318), .O(gate450inter1));
  and2  gate2775(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2776(.a(s_318), .O(gate450inter3));
  inv1  gate2777(.a(s_319), .O(gate450inter4));
  nand2 gate2778(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2779(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2780(.a(G1081), .O(gate450inter7));
  inv1  gate2781(.a(G1177), .O(gate450inter8));
  nand2 gate2782(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2783(.a(s_319), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2784(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2785(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2786(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1485(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1486(.a(gate451inter0), .b(s_134), .O(gate451inter1));
  and2  gate1487(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1488(.a(s_134), .O(gate451inter3));
  inv1  gate1489(.a(s_135), .O(gate451inter4));
  nand2 gate1490(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1491(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1492(.a(G17), .O(gate451inter7));
  inv1  gate1493(.a(G1180), .O(gate451inter8));
  nand2 gate1494(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1495(.a(s_135), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1496(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1497(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1498(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate729(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate730(.a(gate453inter0), .b(s_26), .O(gate453inter1));
  and2  gate731(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate732(.a(s_26), .O(gate453inter3));
  inv1  gate733(.a(s_27), .O(gate453inter4));
  nand2 gate734(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate735(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate736(.a(G18), .O(gate453inter7));
  inv1  gate737(.a(G1183), .O(gate453inter8));
  nand2 gate738(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate739(.a(s_27), .b(gate453inter3), .O(gate453inter10));
  nor2  gate740(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate741(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate742(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2745(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2746(.a(gate457inter0), .b(s_314), .O(gate457inter1));
  and2  gate2747(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2748(.a(s_314), .O(gate457inter3));
  inv1  gate2749(.a(s_315), .O(gate457inter4));
  nand2 gate2750(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2751(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2752(.a(G20), .O(gate457inter7));
  inv1  gate2753(.a(G1189), .O(gate457inter8));
  nand2 gate2754(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2755(.a(s_315), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2756(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2757(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2758(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate911(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate912(.a(gate459inter0), .b(s_52), .O(gate459inter1));
  and2  gate913(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate914(.a(s_52), .O(gate459inter3));
  inv1  gate915(.a(s_53), .O(gate459inter4));
  nand2 gate916(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate917(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate918(.a(G21), .O(gate459inter7));
  inv1  gate919(.a(G1192), .O(gate459inter8));
  nand2 gate920(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate921(.a(s_53), .b(gate459inter3), .O(gate459inter10));
  nor2  gate922(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate923(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate924(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1009(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1010(.a(gate460inter0), .b(s_66), .O(gate460inter1));
  and2  gate1011(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1012(.a(s_66), .O(gate460inter3));
  inv1  gate1013(.a(s_67), .O(gate460inter4));
  nand2 gate1014(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1015(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1016(.a(G1096), .O(gate460inter7));
  inv1  gate1017(.a(G1192), .O(gate460inter8));
  nand2 gate1018(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1019(.a(s_67), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1020(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1021(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1022(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2787(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2788(.a(gate462inter0), .b(s_320), .O(gate462inter1));
  and2  gate2789(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2790(.a(s_320), .O(gate462inter3));
  inv1  gate2791(.a(s_321), .O(gate462inter4));
  nand2 gate2792(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2793(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2794(.a(G1099), .O(gate462inter7));
  inv1  gate2795(.a(G1195), .O(gate462inter8));
  nand2 gate2796(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2797(.a(s_321), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2798(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2799(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2800(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1107(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1108(.a(gate463inter0), .b(s_80), .O(gate463inter1));
  and2  gate1109(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1110(.a(s_80), .O(gate463inter3));
  inv1  gate1111(.a(s_81), .O(gate463inter4));
  nand2 gate1112(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1113(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1114(.a(G23), .O(gate463inter7));
  inv1  gate1115(.a(G1198), .O(gate463inter8));
  nand2 gate1116(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1117(.a(s_81), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1118(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1119(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1120(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1541(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1542(.a(gate466inter0), .b(s_142), .O(gate466inter1));
  and2  gate1543(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1544(.a(s_142), .O(gate466inter3));
  inv1  gate1545(.a(s_143), .O(gate466inter4));
  nand2 gate1546(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1547(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1548(.a(G1105), .O(gate466inter7));
  inv1  gate1549(.a(G1201), .O(gate466inter8));
  nand2 gate1550(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1551(.a(s_143), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1552(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1553(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1554(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2129(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2130(.a(gate467inter0), .b(s_226), .O(gate467inter1));
  and2  gate2131(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2132(.a(s_226), .O(gate467inter3));
  inv1  gate2133(.a(s_227), .O(gate467inter4));
  nand2 gate2134(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2135(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2136(.a(G25), .O(gate467inter7));
  inv1  gate2137(.a(G1204), .O(gate467inter8));
  nand2 gate2138(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2139(.a(s_227), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2140(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2141(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2142(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate2717(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2718(.a(gate468inter0), .b(s_310), .O(gate468inter1));
  and2  gate2719(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2720(.a(s_310), .O(gate468inter3));
  inv1  gate2721(.a(s_311), .O(gate468inter4));
  nand2 gate2722(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2723(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2724(.a(G1108), .O(gate468inter7));
  inv1  gate2725(.a(G1204), .O(gate468inter8));
  nand2 gate2726(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2727(.a(s_311), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2728(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2729(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2730(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1065(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1066(.a(gate470inter0), .b(s_74), .O(gate470inter1));
  and2  gate1067(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1068(.a(s_74), .O(gate470inter3));
  inv1  gate1069(.a(s_75), .O(gate470inter4));
  nand2 gate1070(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1071(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1072(.a(G1111), .O(gate470inter7));
  inv1  gate1073(.a(G1207), .O(gate470inter8));
  nand2 gate1074(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1075(.a(s_75), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1076(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1077(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1078(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1555(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1556(.a(gate472inter0), .b(s_144), .O(gate472inter1));
  and2  gate1557(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1558(.a(s_144), .O(gate472inter3));
  inv1  gate1559(.a(s_145), .O(gate472inter4));
  nand2 gate1560(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1561(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1562(.a(G1114), .O(gate472inter7));
  inv1  gate1563(.a(G1210), .O(gate472inter8));
  nand2 gate1564(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1565(.a(s_145), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1566(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1567(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1568(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate799(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate800(.a(gate479inter0), .b(s_36), .O(gate479inter1));
  and2  gate801(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate802(.a(s_36), .O(gate479inter3));
  inv1  gate803(.a(s_37), .O(gate479inter4));
  nand2 gate804(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate805(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate806(.a(G31), .O(gate479inter7));
  inv1  gate807(.a(G1222), .O(gate479inter8));
  nand2 gate808(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate809(.a(s_37), .b(gate479inter3), .O(gate479inter10));
  nor2  gate810(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate811(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate812(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1625(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1626(.a(gate484inter0), .b(s_154), .O(gate484inter1));
  and2  gate1627(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1628(.a(s_154), .O(gate484inter3));
  inv1  gate1629(.a(s_155), .O(gate484inter4));
  nand2 gate1630(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1631(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1632(.a(G1230), .O(gate484inter7));
  inv1  gate1633(.a(G1231), .O(gate484inter8));
  nand2 gate1634(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1635(.a(s_155), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1636(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1637(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1638(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2857(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2858(.a(gate488inter0), .b(s_330), .O(gate488inter1));
  and2  gate2859(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2860(.a(s_330), .O(gate488inter3));
  inv1  gate2861(.a(s_331), .O(gate488inter4));
  nand2 gate2862(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2863(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2864(.a(G1238), .O(gate488inter7));
  inv1  gate2865(.a(G1239), .O(gate488inter8));
  nand2 gate2866(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2867(.a(s_331), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2868(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2869(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2870(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate645(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate646(.a(gate490inter0), .b(s_14), .O(gate490inter1));
  and2  gate647(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate648(.a(s_14), .O(gate490inter3));
  inv1  gate649(.a(s_15), .O(gate490inter4));
  nand2 gate650(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate651(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate652(.a(G1242), .O(gate490inter7));
  inv1  gate653(.a(G1243), .O(gate490inter8));
  nand2 gate654(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate655(.a(s_15), .b(gate490inter3), .O(gate490inter10));
  nor2  gate656(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate657(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate658(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2507(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2508(.a(gate492inter0), .b(s_280), .O(gate492inter1));
  and2  gate2509(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2510(.a(s_280), .O(gate492inter3));
  inv1  gate2511(.a(s_281), .O(gate492inter4));
  nand2 gate2512(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2513(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2514(.a(G1246), .O(gate492inter7));
  inv1  gate2515(.a(G1247), .O(gate492inter8));
  nand2 gate2516(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2517(.a(s_281), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2518(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2519(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2520(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2073(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2074(.a(gate497inter0), .b(s_218), .O(gate497inter1));
  and2  gate2075(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2076(.a(s_218), .O(gate497inter3));
  inv1  gate2077(.a(s_219), .O(gate497inter4));
  nand2 gate2078(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2079(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2080(.a(G1256), .O(gate497inter7));
  inv1  gate2081(.a(G1257), .O(gate497inter8));
  nand2 gate2082(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2083(.a(s_219), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2084(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2085(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2086(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate659(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate660(.a(gate498inter0), .b(s_16), .O(gate498inter1));
  and2  gate661(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate662(.a(s_16), .O(gate498inter3));
  inv1  gate663(.a(s_17), .O(gate498inter4));
  nand2 gate664(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate665(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate666(.a(G1258), .O(gate498inter7));
  inv1  gate667(.a(G1259), .O(gate498inter8));
  nand2 gate668(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate669(.a(s_17), .b(gate498inter3), .O(gate498inter10));
  nor2  gate670(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate671(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate672(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2521(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2522(.a(gate501inter0), .b(s_282), .O(gate501inter1));
  and2  gate2523(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2524(.a(s_282), .O(gate501inter3));
  inv1  gate2525(.a(s_283), .O(gate501inter4));
  nand2 gate2526(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2527(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2528(.a(G1264), .O(gate501inter7));
  inv1  gate2529(.a(G1265), .O(gate501inter8));
  nand2 gate2530(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2531(.a(s_283), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2532(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2533(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2534(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1429(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1430(.a(gate502inter0), .b(s_126), .O(gate502inter1));
  and2  gate1431(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1432(.a(s_126), .O(gate502inter3));
  inv1  gate1433(.a(s_127), .O(gate502inter4));
  nand2 gate1434(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1435(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1436(.a(G1266), .O(gate502inter7));
  inv1  gate1437(.a(G1267), .O(gate502inter8));
  nand2 gate1438(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1439(.a(s_127), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1440(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1441(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1442(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1933(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1934(.a(gate503inter0), .b(s_198), .O(gate503inter1));
  and2  gate1935(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1936(.a(s_198), .O(gate503inter3));
  inv1  gate1937(.a(s_199), .O(gate503inter4));
  nand2 gate1938(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1939(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1940(.a(G1268), .O(gate503inter7));
  inv1  gate1941(.a(G1269), .O(gate503inter8));
  nand2 gate1942(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1943(.a(s_199), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1944(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1945(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1946(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2619(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2620(.a(gate505inter0), .b(s_296), .O(gate505inter1));
  and2  gate2621(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2622(.a(s_296), .O(gate505inter3));
  inv1  gate2623(.a(s_297), .O(gate505inter4));
  nand2 gate2624(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2625(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2626(.a(G1272), .O(gate505inter7));
  inv1  gate2627(.a(G1273), .O(gate505inter8));
  nand2 gate2628(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2629(.a(s_297), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2630(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2631(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2632(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate561(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate562(.a(gate507inter0), .b(s_2), .O(gate507inter1));
  and2  gate563(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate564(.a(s_2), .O(gate507inter3));
  inv1  gate565(.a(s_3), .O(gate507inter4));
  nand2 gate566(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate567(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate568(.a(G1276), .O(gate507inter7));
  inv1  gate569(.a(G1277), .O(gate507inter8));
  nand2 gate570(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate571(.a(s_3), .b(gate507inter3), .O(gate507inter10));
  nor2  gate572(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate573(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate574(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2759(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2760(.a(gate508inter0), .b(s_316), .O(gate508inter1));
  and2  gate2761(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2762(.a(s_316), .O(gate508inter3));
  inv1  gate2763(.a(s_317), .O(gate508inter4));
  nand2 gate2764(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2765(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2766(.a(G1278), .O(gate508inter7));
  inv1  gate2767(.a(G1279), .O(gate508inter8));
  nand2 gate2768(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2769(.a(s_317), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2770(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2771(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2772(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1051(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1052(.a(gate511inter0), .b(s_72), .O(gate511inter1));
  and2  gate1053(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1054(.a(s_72), .O(gate511inter3));
  inv1  gate1055(.a(s_73), .O(gate511inter4));
  nand2 gate1056(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1057(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1058(.a(G1284), .O(gate511inter7));
  inv1  gate1059(.a(G1285), .O(gate511inter8));
  nand2 gate1060(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1061(.a(s_73), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1062(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1063(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1064(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2003(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2004(.a(gate513inter0), .b(s_208), .O(gate513inter1));
  and2  gate2005(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2006(.a(s_208), .O(gate513inter3));
  inv1  gate2007(.a(s_209), .O(gate513inter4));
  nand2 gate2008(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2009(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2010(.a(G1288), .O(gate513inter7));
  inv1  gate2011(.a(G1289), .O(gate513inter8));
  nand2 gate2012(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2013(.a(s_209), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2014(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2015(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2016(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate2815(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2816(.a(gate514inter0), .b(s_324), .O(gate514inter1));
  and2  gate2817(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2818(.a(s_324), .O(gate514inter3));
  inv1  gate2819(.a(s_325), .O(gate514inter4));
  nand2 gate2820(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2821(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2822(.a(G1290), .O(gate514inter7));
  inv1  gate2823(.a(G1291), .O(gate514inter8));
  nand2 gate2824(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2825(.a(s_325), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2826(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2827(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2828(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule