module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2367(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2368(.a(gate10inter0), .b(s_260), .O(gate10inter1));
  and2  gate2369(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2370(.a(s_260), .O(gate10inter3));
  inv1  gate2371(.a(s_261), .O(gate10inter4));
  nand2 gate2372(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2373(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2374(.a(G3), .O(gate10inter7));
  inv1  gate2375(.a(G4), .O(gate10inter8));
  nand2 gate2376(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2377(.a(s_261), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2378(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2379(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2380(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2479(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2480(.a(gate12inter0), .b(s_276), .O(gate12inter1));
  and2  gate2481(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2482(.a(s_276), .O(gate12inter3));
  inv1  gate2483(.a(s_277), .O(gate12inter4));
  nand2 gate2484(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2485(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2486(.a(G7), .O(gate12inter7));
  inv1  gate2487(.a(G8), .O(gate12inter8));
  nand2 gate2488(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2489(.a(s_277), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2490(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2491(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2492(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1233(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1234(.a(gate16inter0), .b(s_98), .O(gate16inter1));
  and2  gate1235(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1236(.a(s_98), .O(gate16inter3));
  inv1  gate1237(.a(s_99), .O(gate16inter4));
  nand2 gate1238(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1239(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1240(.a(G15), .O(gate16inter7));
  inv1  gate1241(.a(G16), .O(gate16inter8));
  nand2 gate1242(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1243(.a(s_99), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1244(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1245(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1246(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate659(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate660(.a(gate18inter0), .b(s_16), .O(gate18inter1));
  and2  gate661(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate662(.a(s_16), .O(gate18inter3));
  inv1  gate663(.a(s_17), .O(gate18inter4));
  nand2 gate664(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate665(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate666(.a(G19), .O(gate18inter7));
  inv1  gate667(.a(G20), .O(gate18inter8));
  nand2 gate668(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate669(.a(s_17), .b(gate18inter3), .O(gate18inter10));
  nor2  gate670(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate671(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate672(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1793(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1794(.a(gate20inter0), .b(s_178), .O(gate20inter1));
  and2  gate1795(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1796(.a(s_178), .O(gate20inter3));
  inv1  gate1797(.a(s_179), .O(gate20inter4));
  nand2 gate1798(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1799(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1800(.a(G23), .O(gate20inter7));
  inv1  gate1801(.a(G24), .O(gate20inter8));
  nand2 gate1802(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1803(.a(s_179), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1804(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1805(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1806(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2619(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2620(.a(gate22inter0), .b(s_296), .O(gate22inter1));
  and2  gate2621(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2622(.a(s_296), .O(gate22inter3));
  inv1  gate2623(.a(s_297), .O(gate22inter4));
  nand2 gate2624(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2625(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2626(.a(G27), .O(gate22inter7));
  inv1  gate2627(.a(G28), .O(gate22inter8));
  nand2 gate2628(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2629(.a(s_297), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2630(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2631(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2632(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1415(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1416(.a(gate24inter0), .b(s_124), .O(gate24inter1));
  and2  gate1417(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1418(.a(s_124), .O(gate24inter3));
  inv1  gate1419(.a(s_125), .O(gate24inter4));
  nand2 gate1420(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1421(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1422(.a(G31), .O(gate24inter7));
  inv1  gate1423(.a(G32), .O(gate24inter8));
  nand2 gate1424(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1425(.a(s_125), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1426(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1427(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1428(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1177(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1178(.a(gate32inter0), .b(s_90), .O(gate32inter1));
  and2  gate1179(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1180(.a(s_90), .O(gate32inter3));
  inv1  gate1181(.a(s_91), .O(gate32inter4));
  nand2 gate1182(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1183(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1184(.a(G12), .O(gate32inter7));
  inv1  gate1185(.a(G16), .O(gate32inter8));
  nand2 gate1186(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1187(.a(s_91), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1188(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1189(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1190(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate617(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate618(.a(gate35inter0), .b(s_10), .O(gate35inter1));
  and2  gate619(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate620(.a(s_10), .O(gate35inter3));
  inv1  gate621(.a(s_11), .O(gate35inter4));
  nand2 gate622(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate623(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate624(.a(G18), .O(gate35inter7));
  inv1  gate625(.a(G22), .O(gate35inter8));
  nand2 gate626(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate627(.a(s_11), .b(gate35inter3), .O(gate35inter10));
  nor2  gate628(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate629(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate630(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1121(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1122(.a(gate46inter0), .b(s_82), .O(gate46inter1));
  and2  gate1123(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1124(.a(s_82), .O(gate46inter3));
  inv1  gate1125(.a(s_83), .O(gate46inter4));
  nand2 gate1126(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1127(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1128(.a(G6), .O(gate46inter7));
  inv1  gate1129(.a(G272), .O(gate46inter8));
  nand2 gate1130(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1131(.a(s_83), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1132(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1133(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1134(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2171(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2172(.a(gate47inter0), .b(s_232), .O(gate47inter1));
  and2  gate2173(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2174(.a(s_232), .O(gate47inter3));
  inv1  gate2175(.a(s_233), .O(gate47inter4));
  nand2 gate2176(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2177(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2178(.a(G7), .O(gate47inter7));
  inv1  gate2179(.a(G275), .O(gate47inter8));
  nand2 gate2180(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2181(.a(s_233), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2182(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2183(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2184(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate645(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate646(.a(gate53inter0), .b(s_14), .O(gate53inter1));
  and2  gate647(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate648(.a(s_14), .O(gate53inter3));
  inv1  gate649(.a(s_15), .O(gate53inter4));
  nand2 gate650(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate651(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate652(.a(G13), .O(gate53inter7));
  inv1  gate653(.a(G284), .O(gate53inter8));
  nand2 gate654(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate655(.a(s_15), .b(gate53inter3), .O(gate53inter10));
  nor2  gate656(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate657(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate658(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate687(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate688(.a(gate54inter0), .b(s_20), .O(gate54inter1));
  and2  gate689(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate690(.a(s_20), .O(gate54inter3));
  inv1  gate691(.a(s_21), .O(gate54inter4));
  nand2 gate692(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate693(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate694(.a(G14), .O(gate54inter7));
  inv1  gate695(.a(G284), .O(gate54inter8));
  nand2 gate696(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate697(.a(s_21), .b(gate54inter3), .O(gate54inter10));
  nor2  gate698(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate699(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate700(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2563(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2564(.a(gate58inter0), .b(s_288), .O(gate58inter1));
  and2  gate2565(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2566(.a(s_288), .O(gate58inter3));
  inv1  gate2567(.a(s_289), .O(gate58inter4));
  nand2 gate2568(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2569(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2570(.a(G18), .O(gate58inter7));
  inv1  gate2571(.a(G290), .O(gate58inter8));
  nand2 gate2572(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2573(.a(s_289), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2574(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2575(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2576(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate939(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate940(.a(gate60inter0), .b(s_56), .O(gate60inter1));
  and2  gate941(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate942(.a(s_56), .O(gate60inter3));
  inv1  gate943(.a(s_57), .O(gate60inter4));
  nand2 gate944(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate945(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate946(.a(G20), .O(gate60inter7));
  inv1  gate947(.a(G293), .O(gate60inter8));
  nand2 gate948(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate949(.a(s_57), .b(gate60inter3), .O(gate60inter10));
  nor2  gate950(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate951(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate952(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1555(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1556(.a(gate61inter0), .b(s_144), .O(gate61inter1));
  and2  gate1557(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1558(.a(s_144), .O(gate61inter3));
  inv1  gate1559(.a(s_145), .O(gate61inter4));
  nand2 gate1560(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1561(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1562(.a(G21), .O(gate61inter7));
  inv1  gate1563(.a(G296), .O(gate61inter8));
  nand2 gate1564(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1565(.a(s_145), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1566(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1567(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1568(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate953(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate954(.a(gate64inter0), .b(s_58), .O(gate64inter1));
  and2  gate955(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate956(.a(s_58), .O(gate64inter3));
  inv1  gate957(.a(s_59), .O(gate64inter4));
  nand2 gate958(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate959(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate960(.a(G24), .O(gate64inter7));
  inv1  gate961(.a(G299), .O(gate64inter8));
  nand2 gate962(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate963(.a(s_59), .b(gate64inter3), .O(gate64inter10));
  nor2  gate964(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate965(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate966(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1499(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1500(.a(gate70inter0), .b(s_136), .O(gate70inter1));
  and2  gate1501(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1502(.a(s_136), .O(gate70inter3));
  inv1  gate1503(.a(s_137), .O(gate70inter4));
  nand2 gate1504(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1505(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1506(.a(G30), .O(gate70inter7));
  inv1  gate1507(.a(G308), .O(gate70inter8));
  nand2 gate1508(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1509(.a(s_137), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1510(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1511(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1512(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2353(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2354(.a(gate72inter0), .b(s_258), .O(gate72inter1));
  and2  gate2355(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2356(.a(s_258), .O(gate72inter3));
  inv1  gate2357(.a(s_259), .O(gate72inter4));
  nand2 gate2358(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2359(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2360(.a(G32), .O(gate72inter7));
  inv1  gate2361(.a(G311), .O(gate72inter8));
  nand2 gate2362(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2363(.a(s_259), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2364(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2365(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2366(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate2199(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2200(.a(gate73inter0), .b(s_236), .O(gate73inter1));
  and2  gate2201(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2202(.a(s_236), .O(gate73inter3));
  inv1  gate2203(.a(s_237), .O(gate73inter4));
  nand2 gate2204(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2205(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2206(.a(G1), .O(gate73inter7));
  inv1  gate2207(.a(G314), .O(gate73inter8));
  nand2 gate2208(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2209(.a(s_237), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2210(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2211(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2212(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1961(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1962(.a(gate75inter0), .b(s_202), .O(gate75inter1));
  and2  gate1963(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1964(.a(s_202), .O(gate75inter3));
  inv1  gate1965(.a(s_203), .O(gate75inter4));
  nand2 gate1966(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1967(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1968(.a(G9), .O(gate75inter7));
  inv1  gate1969(.a(G317), .O(gate75inter8));
  nand2 gate1970(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1971(.a(s_203), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1972(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1973(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1974(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2227(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2228(.a(gate89inter0), .b(s_240), .O(gate89inter1));
  and2  gate2229(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2230(.a(s_240), .O(gate89inter3));
  inv1  gate2231(.a(s_241), .O(gate89inter4));
  nand2 gate2232(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2233(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2234(.a(G17), .O(gate89inter7));
  inv1  gate2235(.a(G338), .O(gate89inter8));
  nand2 gate2236(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2237(.a(s_241), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2238(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2239(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2240(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1625(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1626(.a(gate92inter0), .b(s_154), .O(gate92inter1));
  and2  gate1627(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1628(.a(s_154), .O(gate92inter3));
  inv1  gate1629(.a(s_155), .O(gate92inter4));
  nand2 gate1630(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1631(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1632(.a(G29), .O(gate92inter7));
  inv1  gate1633(.a(G341), .O(gate92inter8));
  nand2 gate1634(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1635(.a(s_155), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1636(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1637(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1638(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2493(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2494(.a(gate96inter0), .b(s_278), .O(gate96inter1));
  and2  gate2495(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2496(.a(s_278), .O(gate96inter3));
  inv1  gate2497(.a(s_279), .O(gate96inter4));
  nand2 gate2498(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2499(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2500(.a(G30), .O(gate96inter7));
  inv1  gate2501(.a(G347), .O(gate96inter8));
  nand2 gate2502(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2503(.a(s_279), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2504(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2505(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2506(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate757(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate758(.a(gate103inter0), .b(s_30), .O(gate103inter1));
  and2  gate759(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate760(.a(s_30), .O(gate103inter3));
  inv1  gate761(.a(s_31), .O(gate103inter4));
  nand2 gate762(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate763(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate764(.a(G28), .O(gate103inter7));
  inv1  gate765(.a(G359), .O(gate103inter8));
  nand2 gate766(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate767(.a(s_31), .b(gate103inter3), .O(gate103inter10));
  nor2  gate768(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate769(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate770(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2073(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2074(.a(gate107inter0), .b(s_218), .O(gate107inter1));
  and2  gate2075(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2076(.a(s_218), .O(gate107inter3));
  inv1  gate2077(.a(s_219), .O(gate107inter4));
  nand2 gate2078(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2079(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2080(.a(G366), .O(gate107inter7));
  inv1  gate2081(.a(G367), .O(gate107inter8));
  nand2 gate2082(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2083(.a(s_219), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2084(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2085(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2086(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate2185(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2186(.a(gate108inter0), .b(s_234), .O(gate108inter1));
  and2  gate2187(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2188(.a(s_234), .O(gate108inter3));
  inv1  gate2189(.a(s_235), .O(gate108inter4));
  nand2 gate2190(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2191(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2192(.a(G368), .O(gate108inter7));
  inv1  gate2193(.a(G369), .O(gate108inter8));
  nand2 gate2194(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2195(.a(s_235), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2196(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2197(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2198(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate2325(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2326(.a(gate109inter0), .b(s_254), .O(gate109inter1));
  and2  gate2327(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2328(.a(s_254), .O(gate109inter3));
  inv1  gate2329(.a(s_255), .O(gate109inter4));
  nand2 gate2330(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2331(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2332(.a(G370), .O(gate109inter7));
  inv1  gate2333(.a(G371), .O(gate109inter8));
  nand2 gate2334(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2335(.a(s_255), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2336(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2337(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2338(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1835(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1836(.a(gate110inter0), .b(s_184), .O(gate110inter1));
  and2  gate1837(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1838(.a(s_184), .O(gate110inter3));
  inv1  gate1839(.a(s_185), .O(gate110inter4));
  nand2 gate1840(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1841(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1842(.a(G372), .O(gate110inter7));
  inv1  gate1843(.a(G373), .O(gate110inter8));
  nand2 gate1844(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1845(.a(s_185), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1846(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1847(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1848(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1975(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1976(.a(gate114inter0), .b(s_204), .O(gate114inter1));
  and2  gate1977(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1978(.a(s_204), .O(gate114inter3));
  inv1  gate1979(.a(s_205), .O(gate114inter4));
  nand2 gate1980(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1981(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1982(.a(G380), .O(gate114inter7));
  inv1  gate1983(.a(G381), .O(gate114inter8));
  nand2 gate1984(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1985(.a(s_205), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1986(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1987(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1988(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate729(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate730(.a(gate116inter0), .b(s_26), .O(gate116inter1));
  and2  gate731(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate732(.a(s_26), .O(gate116inter3));
  inv1  gate733(.a(s_27), .O(gate116inter4));
  nand2 gate734(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate735(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate736(.a(G384), .O(gate116inter7));
  inv1  gate737(.a(G385), .O(gate116inter8));
  nand2 gate738(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate739(.a(s_27), .b(gate116inter3), .O(gate116inter10));
  nor2  gate740(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate741(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate742(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1611(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1612(.a(gate120inter0), .b(s_152), .O(gate120inter1));
  and2  gate1613(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1614(.a(s_152), .O(gate120inter3));
  inv1  gate1615(.a(s_153), .O(gate120inter4));
  nand2 gate1616(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1617(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1618(.a(G392), .O(gate120inter7));
  inv1  gate1619(.a(G393), .O(gate120inter8));
  nand2 gate1620(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1621(.a(s_153), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1622(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1623(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1624(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2423(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2424(.a(gate123inter0), .b(s_268), .O(gate123inter1));
  and2  gate2425(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2426(.a(s_268), .O(gate123inter3));
  inv1  gate2427(.a(s_269), .O(gate123inter4));
  nand2 gate2428(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2429(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2430(.a(G398), .O(gate123inter7));
  inv1  gate2431(.a(G399), .O(gate123inter8));
  nand2 gate2432(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2433(.a(s_269), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2434(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2435(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2436(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1443(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1444(.a(gate124inter0), .b(s_128), .O(gate124inter1));
  and2  gate1445(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1446(.a(s_128), .O(gate124inter3));
  inv1  gate1447(.a(s_129), .O(gate124inter4));
  nand2 gate1448(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1449(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1450(.a(G400), .O(gate124inter7));
  inv1  gate1451(.a(G401), .O(gate124inter8));
  nand2 gate1452(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1453(.a(s_129), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1454(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1455(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1456(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1877(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1878(.a(gate126inter0), .b(s_190), .O(gate126inter1));
  and2  gate1879(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1880(.a(s_190), .O(gate126inter3));
  inv1  gate1881(.a(s_191), .O(gate126inter4));
  nand2 gate1882(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1883(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1884(.a(G404), .O(gate126inter7));
  inv1  gate1885(.a(G405), .O(gate126inter8));
  nand2 gate1886(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1887(.a(s_191), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1888(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1889(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1890(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2605(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2606(.a(gate128inter0), .b(s_294), .O(gate128inter1));
  and2  gate2607(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2608(.a(s_294), .O(gate128inter3));
  inv1  gate2609(.a(s_295), .O(gate128inter4));
  nand2 gate2610(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2611(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2612(.a(G408), .O(gate128inter7));
  inv1  gate2613(.a(G409), .O(gate128inter8));
  nand2 gate2614(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2615(.a(s_295), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2616(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2617(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2618(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2311(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2312(.a(gate138inter0), .b(s_252), .O(gate138inter1));
  and2  gate2313(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2314(.a(s_252), .O(gate138inter3));
  inv1  gate2315(.a(s_253), .O(gate138inter4));
  nand2 gate2316(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2317(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2318(.a(G432), .O(gate138inter7));
  inv1  gate2319(.a(G435), .O(gate138inter8));
  nand2 gate2320(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2321(.a(s_253), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2322(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2323(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2324(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2535(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2536(.a(gate141inter0), .b(s_284), .O(gate141inter1));
  and2  gate2537(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2538(.a(s_284), .O(gate141inter3));
  inv1  gate2539(.a(s_285), .O(gate141inter4));
  nand2 gate2540(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2541(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2542(.a(G450), .O(gate141inter7));
  inv1  gate2543(.a(G453), .O(gate141inter8));
  nand2 gate2544(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2545(.a(s_285), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2546(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2547(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2548(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1569(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1570(.a(gate145inter0), .b(s_146), .O(gate145inter1));
  and2  gate1571(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1572(.a(s_146), .O(gate145inter3));
  inv1  gate1573(.a(s_147), .O(gate145inter4));
  nand2 gate1574(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1575(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1576(.a(G474), .O(gate145inter7));
  inv1  gate1577(.a(G477), .O(gate145inter8));
  nand2 gate1578(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1579(.a(s_147), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1580(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1581(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1582(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1009(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1010(.a(gate149inter0), .b(s_66), .O(gate149inter1));
  and2  gate1011(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1012(.a(s_66), .O(gate149inter3));
  inv1  gate1013(.a(s_67), .O(gate149inter4));
  nand2 gate1014(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1015(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1016(.a(G498), .O(gate149inter7));
  inv1  gate1017(.a(G501), .O(gate149inter8));
  nand2 gate1018(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1019(.a(s_67), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1020(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1021(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1022(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1779(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1780(.a(gate150inter0), .b(s_176), .O(gate150inter1));
  and2  gate1781(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1782(.a(s_176), .O(gate150inter3));
  inv1  gate1783(.a(s_177), .O(gate150inter4));
  nand2 gate1784(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1785(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1786(.a(G504), .O(gate150inter7));
  inv1  gate1787(.a(G507), .O(gate150inter8));
  nand2 gate1788(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1789(.a(s_177), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1790(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1791(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1792(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1919(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1920(.a(gate151inter0), .b(s_196), .O(gate151inter1));
  and2  gate1921(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1922(.a(s_196), .O(gate151inter3));
  inv1  gate1923(.a(s_197), .O(gate151inter4));
  nand2 gate1924(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1925(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1926(.a(G510), .O(gate151inter7));
  inv1  gate1927(.a(G513), .O(gate151inter8));
  nand2 gate1928(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1929(.a(s_197), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1930(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1931(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1932(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate561(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate562(.a(gate152inter0), .b(s_2), .O(gate152inter1));
  and2  gate563(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate564(.a(s_2), .O(gate152inter3));
  inv1  gate565(.a(s_3), .O(gate152inter4));
  nand2 gate566(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate567(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate568(.a(G516), .O(gate152inter7));
  inv1  gate569(.a(G519), .O(gate152inter8));
  nand2 gate570(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate571(.a(s_3), .b(gate152inter3), .O(gate152inter10));
  nor2  gate572(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate573(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate574(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate883(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate884(.a(gate154inter0), .b(s_48), .O(gate154inter1));
  and2  gate885(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate886(.a(s_48), .O(gate154inter3));
  inv1  gate887(.a(s_49), .O(gate154inter4));
  nand2 gate888(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate889(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate890(.a(G429), .O(gate154inter7));
  inv1  gate891(.a(G522), .O(gate154inter8));
  nand2 gate892(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate893(.a(s_49), .b(gate154inter3), .O(gate154inter10));
  nor2  gate894(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate895(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate896(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2549(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2550(.a(gate156inter0), .b(s_286), .O(gate156inter1));
  and2  gate2551(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2552(.a(s_286), .O(gate156inter3));
  inv1  gate2553(.a(s_287), .O(gate156inter4));
  nand2 gate2554(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2555(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2556(.a(G435), .O(gate156inter7));
  inv1  gate2557(.a(G525), .O(gate156inter8));
  nand2 gate2558(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2559(.a(s_287), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2560(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2561(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2562(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1891(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1892(.a(gate158inter0), .b(s_192), .O(gate158inter1));
  and2  gate1893(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1894(.a(s_192), .O(gate158inter3));
  inv1  gate1895(.a(s_193), .O(gate158inter4));
  nand2 gate1896(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1897(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1898(.a(G441), .O(gate158inter7));
  inv1  gate1899(.a(G528), .O(gate158inter8));
  nand2 gate1900(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1901(.a(s_193), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1902(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1903(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1904(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2241(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2242(.a(gate160inter0), .b(s_242), .O(gate160inter1));
  and2  gate2243(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2244(.a(s_242), .O(gate160inter3));
  inv1  gate2245(.a(s_243), .O(gate160inter4));
  nand2 gate2246(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2247(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2248(.a(G447), .O(gate160inter7));
  inv1  gate2249(.a(G531), .O(gate160inter8));
  nand2 gate2250(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2251(.a(s_243), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2252(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2253(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2254(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1737(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1738(.a(gate161inter0), .b(s_170), .O(gate161inter1));
  and2  gate1739(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1740(.a(s_170), .O(gate161inter3));
  inv1  gate1741(.a(s_171), .O(gate161inter4));
  nand2 gate1742(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1743(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1744(.a(G450), .O(gate161inter7));
  inv1  gate1745(.a(G534), .O(gate161inter8));
  nand2 gate1746(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1747(.a(s_171), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1748(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1749(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1750(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1807(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1808(.a(gate164inter0), .b(s_180), .O(gate164inter1));
  and2  gate1809(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1810(.a(s_180), .O(gate164inter3));
  inv1  gate1811(.a(s_181), .O(gate164inter4));
  nand2 gate1812(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1813(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1814(.a(G459), .O(gate164inter7));
  inv1  gate1815(.a(G537), .O(gate164inter8));
  nand2 gate1816(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1817(.a(s_181), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1818(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1819(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1820(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate2269(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2270(.a(gate165inter0), .b(s_246), .O(gate165inter1));
  and2  gate2271(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2272(.a(s_246), .O(gate165inter3));
  inv1  gate2273(.a(s_247), .O(gate165inter4));
  nand2 gate2274(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2275(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2276(.a(G462), .O(gate165inter7));
  inv1  gate2277(.a(G540), .O(gate165inter8));
  nand2 gate2278(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2279(.a(s_247), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2280(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2281(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2282(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2087(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2088(.a(gate168inter0), .b(s_220), .O(gate168inter1));
  and2  gate2089(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2090(.a(s_220), .O(gate168inter3));
  inv1  gate2091(.a(s_221), .O(gate168inter4));
  nand2 gate2092(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2093(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2094(.a(G471), .O(gate168inter7));
  inv1  gate2095(.a(G543), .O(gate168inter8));
  nand2 gate2096(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2097(.a(s_221), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2098(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2099(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2100(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2143(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2144(.a(gate170inter0), .b(s_228), .O(gate170inter1));
  and2  gate2145(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2146(.a(s_228), .O(gate170inter3));
  inv1  gate2147(.a(s_229), .O(gate170inter4));
  nand2 gate2148(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2149(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2150(.a(G477), .O(gate170inter7));
  inv1  gate2151(.a(G546), .O(gate170inter8));
  nand2 gate2152(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2153(.a(s_229), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2154(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2155(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2156(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2451(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2452(.a(gate173inter0), .b(s_272), .O(gate173inter1));
  and2  gate2453(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2454(.a(s_272), .O(gate173inter3));
  inv1  gate2455(.a(s_273), .O(gate173inter4));
  nand2 gate2456(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2457(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2458(.a(G486), .O(gate173inter7));
  inv1  gate2459(.a(G552), .O(gate173inter8));
  nand2 gate2460(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2461(.a(s_273), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2462(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2463(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2464(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2101(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2102(.a(gate176inter0), .b(s_222), .O(gate176inter1));
  and2  gate2103(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2104(.a(s_222), .O(gate176inter3));
  inv1  gate2105(.a(s_223), .O(gate176inter4));
  nand2 gate2106(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2107(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2108(.a(G495), .O(gate176inter7));
  inv1  gate2109(.a(G555), .O(gate176inter8));
  nand2 gate2110(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2111(.a(s_223), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2112(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2113(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2114(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate1933(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1934(.a(gate177inter0), .b(s_198), .O(gate177inter1));
  and2  gate1935(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1936(.a(s_198), .O(gate177inter3));
  inv1  gate1937(.a(s_199), .O(gate177inter4));
  nand2 gate1938(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1939(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1940(.a(G498), .O(gate177inter7));
  inv1  gate1941(.a(G558), .O(gate177inter8));
  nand2 gate1942(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1943(.a(s_199), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1944(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1945(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1946(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1247(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1248(.a(gate187inter0), .b(s_100), .O(gate187inter1));
  and2  gate1249(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1250(.a(s_100), .O(gate187inter3));
  inv1  gate1251(.a(s_101), .O(gate187inter4));
  nand2 gate1252(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1253(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1254(.a(G574), .O(gate187inter7));
  inv1  gate1255(.a(G575), .O(gate187inter8));
  nand2 gate1256(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1257(.a(s_101), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1258(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1259(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1260(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1345(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1346(.a(gate188inter0), .b(s_114), .O(gate188inter1));
  and2  gate1347(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1348(.a(s_114), .O(gate188inter3));
  inv1  gate1349(.a(s_115), .O(gate188inter4));
  nand2 gate1350(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1351(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1352(.a(G576), .O(gate188inter7));
  inv1  gate1353(.a(G577), .O(gate188inter8));
  nand2 gate1354(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1355(.a(s_115), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1356(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1357(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1358(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1401(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1402(.a(gate191inter0), .b(s_122), .O(gate191inter1));
  and2  gate1403(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1404(.a(s_122), .O(gate191inter3));
  inv1  gate1405(.a(s_123), .O(gate191inter4));
  nand2 gate1406(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1407(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1408(.a(G582), .O(gate191inter7));
  inv1  gate1409(.a(G583), .O(gate191inter8));
  nand2 gate1410(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1411(.a(s_123), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1412(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1413(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1414(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1373(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1374(.a(gate193inter0), .b(s_118), .O(gate193inter1));
  and2  gate1375(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1376(.a(s_118), .O(gate193inter3));
  inv1  gate1377(.a(s_119), .O(gate193inter4));
  nand2 gate1378(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1379(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1380(.a(G586), .O(gate193inter7));
  inv1  gate1381(.a(G587), .O(gate193inter8));
  nand2 gate1382(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1383(.a(s_119), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1384(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1385(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1386(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2213(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2214(.a(gate195inter0), .b(s_238), .O(gate195inter1));
  and2  gate2215(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2216(.a(s_238), .O(gate195inter3));
  inv1  gate2217(.a(s_239), .O(gate195inter4));
  nand2 gate2218(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2219(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2220(.a(G590), .O(gate195inter7));
  inv1  gate2221(.a(G591), .O(gate195inter8));
  nand2 gate2222(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2223(.a(s_239), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2224(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2225(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2226(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate575(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate576(.a(gate197inter0), .b(s_4), .O(gate197inter1));
  and2  gate577(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate578(.a(s_4), .O(gate197inter3));
  inv1  gate579(.a(s_5), .O(gate197inter4));
  nand2 gate580(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate581(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate582(.a(G594), .O(gate197inter7));
  inv1  gate583(.a(G595), .O(gate197inter8));
  nand2 gate584(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate585(.a(s_5), .b(gate197inter3), .O(gate197inter10));
  nor2  gate586(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate587(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate588(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2115(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2116(.a(gate201inter0), .b(s_224), .O(gate201inter1));
  and2  gate2117(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2118(.a(s_224), .O(gate201inter3));
  inv1  gate2119(.a(s_225), .O(gate201inter4));
  nand2 gate2120(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2121(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2122(.a(G602), .O(gate201inter7));
  inv1  gate2123(.a(G607), .O(gate201inter8));
  nand2 gate2124(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2125(.a(s_225), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2126(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2127(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2128(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate827(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate828(.a(gate203inter0), .b(s_40), .O(gate203inter1));
  and2  gate829(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate830(.a(s_40), .O(gate203inter3));
  inv1  gate831(.a(s_41), .O(gate203inter4));
  nand2 gate832(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate833(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate834(.a(G602), .O(gate203inter7));
  inv1  gate835(.a(G612), .O(gate203inter8));
  nand2 gate836(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate837(.a(s_41), .b(gate203inter3), .O(gate203inter10));
  nor2  gate838(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate839(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate840(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate589(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate590(.a(gate204inter0), .b(s_6), .O(gate204inter1));
  and2  gate591(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate592(.a(s_6), .O(gate204inter3));
  inv1  gate593(.a(s_7), .O(gate204inter4));
  nand2 gate594(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate595(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate596(.a(G607), .O(gate204inter7));
  inv1  gate597(.a(G617), .O(gate204inter8));
  nand2 gate598(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate599(.a(s_7), .b(gate204inter3), .O(gate204inter10));
  nor2  gate600(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate601(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate602(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1037(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1038(.a(gate206inter0), .b(s_70), .O(gate206inter1));
  and2  gate1039(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1040(.a(s_70), .O(gate206inter3));
  inv1  gate1041(.a(s_71), .O(gate206inter4));
  nand2 gate1042(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1043(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1044(.a(G632), .O(gate206inter7));
  inv1  gate1045(.a(G637), .O(gate206inter8));
  nand2 gate1046(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1047(.a(s_71), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1048(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1049(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1050(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2465(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2466(.a(gate210inter0), .b(s_274), .O(gate210inter1));
  and2  gate2467(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2468(.a(s_274), .O(gate210inter3));
  inv1  gate2469(.a(s_275), .O(gate210inter4));
  nand2 gate2470(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2471(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2472(.a(G607), .O(gate210inter7));
  inv1  gate2473(.a(G666), .O(gate210inter8));
  nand2 gate2474(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2475(.a(s_275), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2476(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2477(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2478(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1205(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1206(.a(gate211inter0), .b(s_94), .O(gate211inter1));
  and2  gate1207(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1208(.a(s_94), .O(gate211inter3));
  inv1  gate1209(.a(s_95), .O(gate211inter4));
  nand2 gate1210(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1211(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1212(.a(G612), .O(gate211inter7));
  inv1  gate1213(.a(G669), .O(gate211inter8));
  nand2 gate1214(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1215(.a(s_95), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1216(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1217(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1218(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2381(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2382(.a(gate212inter0), .b(s_262), .O(gate212inter1));
  and2  gate2383(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2384(.a(s_262), .O(gate212inter3));
  inv1  gate2385(.a(s_263), .O(gate212inter4));
  nand2 gate2386(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2387(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2388(.a(G617), .O(gate212inter7));
  inv1  gate2389(.a(G669), .O(gate212inter8));
  nand2 gate2390(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2391(.a(s_263), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2392(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2393(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2394(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1317(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1318(.a(gate213inter0), .b(s_110), .O(gate213inter1));
  and2  gate1319(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1320(.a(s_110), .O(gate213inter3));
  inv1  gate1321(.a(s_111), .O(gate213inter4));
  nand2 gate1322(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1323(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1324(.a(G602), .O(gate213inter7));
  inv1  gate1325(.a(G672), .O(gate213inter8));
  nand2 gate1326(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1327(.a(s_111), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1328(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1329(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1330(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1541(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1542(.a(gate215inter0), .b(s_142), .O(gate215inter1));
  and2  gate1543(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1544(.a(s_142), .O(gate215inter3));
  inv1  gate1545(.a(s_143), .O(gate215inter4));
  nand2 gate1546(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1547(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1548(.a(G607), .O(gate215inter7));
  inv1  gate1549(.a(G675), .O(gate215inter8));
  nand2 gate1550(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1551(.a(s_143), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1552(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1553(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1554(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate911(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate912(.a(gate216inter0), .b(s_52), .O(gate216inter1));
  and2  gate913(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate914(.a(s_52), .O(gate216inter3));
  inv1  gate915(.a(s_53), .O(gate216inter4));
  nand2 gate916(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate917(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate918(.a(G617), .O(gate216inter7));
  inv1  gate919(.a(G675), .O(gate216inter8));
  nand2 gate920(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate921(.a(s_53), .b(gate216inter3), .O(gate216inter10));
  nor2  gate922(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate923(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate924(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1471(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1472(.a(gate218inter0), .b(s_132), .O(gate218inter1));
  and2  gate1473(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1474(.a(s_132), .O(gate218inter3));
  inv1  gate1475(.a(s_133), .O(gate218inter4));
  nand2 gate1476(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1477(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1478(.a(G627), .O(gate218inter7));
  inv1  gate1479(.a(G678), .O(gate218inter8));
  nand2 gate1480(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1481(.a(s_133), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1482(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1483(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1484(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate813(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate814(.a(gate219inter0), .b(s_38), .O(gate219inter1));
  and2  gate815(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate816(.a(s_38), .O(gate219inter3));
  inv1  gate817(.a(s_39), .O(gate219inter4));
  nand2 gate818(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate819(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate820(.a(G632), .O(gate219inter7));
  inv1  gate821(.a(G681), .O(gate219inter8));
  nand2 gate822(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate823(.a(s_39), .b(gate219inter3), .O(gate219inter10));
  nor2  gate824(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate825(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate826(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate2031(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2032(.a(gate221inter0), .b(s_212), .O(gate221inter1));
  and2  gate2033(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2034(.a(s_212), .O(gate221inter3));
  inv1  gate2035(.a(s_213), .O(gate221inter4));
  nand2 gate2036(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2037(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2038(.a(G622), .O(gate221inter7));
  inv1  gate2039(.a(G684), .O(gate221inter8));
  nand2 gate2040(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2041(.a(s_213), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2042(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2043(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2044(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate2507(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2508(.a(gate222inter0), .b(s_280), .O(gate222inter1));
  and2  gate2509(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2510(.a(s_280), .O(gate222inter3));
  inv1  gate2511(.a(s_281), .O(gate222inter4));
  nand2 gate2512(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2513(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2514(.a(G632), .O(gate222inter7));
  inv1  gate2515(.a(G684), .O(gate222inter8));
  nand2 gate2516(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2517(.a(s_281), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2518(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2519(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2520(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1219(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1220(.a(gate226inter0), .b(s_96), .O(gate226inter1));
  and2  gate1221(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1222(.a(s_96), .O(gate226inter3));
  inv1  gate1223(.a(s_97), .O(gate226inter4));
  nand2 gate1224(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1225(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1226(.a(G692), .O(gate226inter7));
  inv1  gate1227(.a(G693), .O(gate226inter8));
  nand2 gate1228(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1229(.a(s_97), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1230(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1231(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1232(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2045(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2046(.a(gate228inter0), .b(s_214), .O(gate228inter1));
  and2  gate2047(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2048(.a(s_214), .O(gate228inter3));
  inv1  gate2049(.a(s_215), .O(gate228inter4));
  nand2 gate2050(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2051(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2052(.a(G696), .O(gate228inter7));
  inv1  gate2053(.a(G697), .O(gate228inter8));
  nand2 gate2054(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2055(.a(s_215), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2056(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2057(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2058(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1051(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1052(.a(gate236inter0), .b(s_72), .O(gate236inter1));
  and2  gate1053(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1054(.a(s_72), .O(gate236inter3));
  inv1  gate1055(.a(s_73), .O(gate236inter4));
  nand2 gate1056(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1057(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1058(.a(G251), .O(gate236inter7));
  inv1  gate1059(.a(G727), .O(gate236inter8));
  nand2 gate1060(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1061(.a(s_73), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1062(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1063(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1064(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1989(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1990(.a(gate237inter0), .b(s_206), .O(gate237inter1));
  and2  gate1991(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1992(.a(s_206), .O(gate237inter3));
  inv1  gate1993(.a(s_207), .O(gate237inter4));
  nand2 gate1994(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1995(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1996(.a(G254), .O(gate237inter7));
  inv1  gate1997(.a(G706), .O(gate237inter8));
  nand2 gate1998(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1999(.a(s_207), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2000(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2001(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2002(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2339(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2340(.a(gate245inter0), .b(s_256), .O(gate245inter1));
  and2  gate2341(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2342(.a(s_256), .O(gate245inter3));
  inv1  gate2343(.a(s_257), .O(gate245inter4));
  nand2 gate2344(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2345(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2346(.a(G248), .O(gate245inter7));
  inv1  gate2347(.a(G736), .O(gate245inter8));
  nand2 gate2348(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2349(.a(s_257), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2350(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2351(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2352(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1275(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1276(.a(gate249inter0), .b(s_104), .O(gate249inter1));
  and2  gate1277(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1278(.a(s_104), .O(gate249inter3));
  inv1  gate1279(.a(s_105), .O(gate249inter4));
  nand2 gate1280(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1281(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1282(.a(G254), .O(gate249inter7));
  inv1  gate1283(.a(G742), .O(gate249inter8));
  nand2 gate1284(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1285(.a(s_105), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1286(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1287(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1288(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1765(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1766(.a(gate250inter0), .b(s_174), .O(gate250inter1));
  and2  gate1767(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1768(.a(s_174), .O(gate250inter3));
  inv1  gate1769(.a(s_175), .O(gate250inter4));
  nand2 gate1770(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1771(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1772(.a(G706), .O(gate250inter7));
  inv1  gate1773(.a(G742), .O(gate250inter8));
  nand2 gate1774(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1775(.a(s_175), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1776(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1777(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1778(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1303(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1304(.a(gate251inter0), .b(s_108), .O(gate251inter1));
  and2  gate1305(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1306(.a(s_108), .O(gate251inter3));
  inv1  gate1307(.a(s_109), .O(gate251inter4));
  nand2 gate1308(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1309(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1310(.a(G257), .O(gate251inter7));
  inv1  gate1311(.a(G745), .O(gate251inter8));
  nand2 gate1312(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1313(.a(s_109), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1314(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1315(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1316(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1149(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1150(.a(gate252inter0), .b(s_86), .O(gate252inter1));
  and2  gate1151(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1152(.a(s_86), .O(gate252inter3));
  inv1  gate1153(.a(s_87), .O(gate252inter4));
  nand2 gate1154(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1155(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1156(.a(G709), .O(gate252inter7));
  inv1  gate1157(.a(G745), .O(gate252inter8));
  nand2 gate1158(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1159(.a(s_87), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1160(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1161(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1162(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1681(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1682(.a(gate256inter0), .b(s_162), .O(gate256inter1));
  and2  gate1683(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1684(.a(s_162), .O(gate256inter3));
  inv1  gate1685(.a(s_163), .O(gate256inter4));
  nand2 gate1686(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1687(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1688(.a(G715), .O(gate256inter7));
  inv1  gate1689(.a(G751), .O(gate256inter8));
  nand2 gate1690(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1691(.a(s_163), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1692(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1693(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1694(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1023(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1024(.a(gate258inter0), .b(s_68), .O(gate258inter1));
  and2  gate1025(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1026(.a(s_68), .O(gate258inter3));
  inv1  gate1027(.a(s_69), .O(gate258inter4));
  nand2 gate1028(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1029(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1030(.a(G756), .O(gate258inter7));
  inv1  gate1031(.a(G757), .O(gate258inter8));
  nand2 gate1032(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1033(.a(s_69), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1034(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1035(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1036(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate995(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate996(.a(gate261inter0), .b(s_64), .O(gate261inter1));
  and2  gate997(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate998(.a(s_64), .O(gate261inter3));
  inv1  gate999(.a(s_65), .O(gate261inter4));
  nand2 gate1000(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1001(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1002(.a(G762), .O(gate261inter7));
  inv1  gate1003(.a(G763), .O(gate261inter8));
  nand2 gate1004(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1005(.a(s_65), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1006(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1007(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1008(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1191(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1192(.a(gate264inter0), .b(s_92), .O(gate264inter1));
  and2  gate1193(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1194(.a(s_92), .O(gate264inter3));
  inv1  gate1195(.a(s_93), .O(gate264inter4));
  nand2 gate1196(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1197(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1198(.a(G768), .O(gate264inter7));
  inv1  gate1199(.a(G769), .O(gate264inter8));
  nand2 gate1200(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1201(.a(s_93), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1202(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1203(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1204(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate855(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate856(.a(gate265inter0), .b(s_44), .O(gate265inter1));
  and2  gate857(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate858(.a(s_44), .O(gate265inter3));
  inv1  gate859(.a(s_45), .O(gate265inter4));
  nand2 gate860(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate861(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate862(.a(G642), .O(gate265inter7));
  inv1  gate863(.a(G770), .O(gate265inter8));
  nand2 gate864(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate865(.a(s_45), .b(gate265inter3), .O(gate265inter10));
  nor2  gate866(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate867(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate868(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1653(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1654(.a(gate267inter0), .b(s_158), .O(gate267inter1));
  and2  gate1655(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1656(.a(s_158), .O(gate267inter3));
  inv1  gate1657(.a(s_159), .O(gate267inter4));
  nand2 gate1658(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1659(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1660(.a(G648), .O(gate267inter7));
  inv1  gate1661(.a(G776), .O(gate267inter8));
  nand2 gate1662(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1663(.a(s_159), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1664(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1665(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1666(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate673(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate674(.a(gate268inter0), .b(s_18), .O(gate268inter1));
  and2  gate675(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate676(.a(s_18), .O(gate268inter3));
  inv1  gate677(.a(s_19), .O(gate268inter4));
  nand2 gate678(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate679(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate680(.a(G651), .O(gate268inter7));
  inv1  gate681(.a(G779), .O(gate268inter8));
  nand2 gate682(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate683(.a(s_19), .b(gate268inter3), .O(gate268inter10));
  nor2  gate684(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate685(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate686(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2521(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2522(.a(gate270inter0), .b(s_282), .O(gate270inter1));
  and2  gate2523(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2524(.a(s_282), .O(gate270inter3));
  inv1  gate2525(.a(s_283), .O(gate270inter4));
  nand2 gate2526(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2527(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2528(.a(G657), .O(gate270inter7));
  inv1  gate2529(.a(G785), .O(gate270inter8));
  nand2 gate2530(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2531(.a(s_283), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2532(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2533(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2534(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2157(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2158(.a(gate276inter0), .b(s_230), .O(gate276inter1));
  and2  gate2159(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2160(.a(s_230), .O(gate276inter3));
  inv1  gate2161(.a(s_231), .O(gate276inter4));
  nand2 gate2162(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2163(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2164(.a(G773), .O(gate276inter7));
  inv1  gate2165(.a(G797), .O(gate276inter8));
  nand2 gate2166(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2167(.a(s_231), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2168(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2169(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2170(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1093(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1094(.a(gate277inter0), .b(s_78), .O(gate277inter1));
  and2  gate1095(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1096(.a(s_78), .O(gate277inter3));
  inv1  gate1097(.a(s_79), .O(gate277inter4));
  nand2 gate1098(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1099(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1100(.a(G648), .O(gate277inter7));
  inv1  gate1101(.a(G800), .O(gate277inter8));
  nand2 gate1102(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1103(.a(s_79), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1104(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1105(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1106(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1583(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1584(.a(gate278inter0), .b(s_148), .O(gate278inter1));
  and2  gate1585(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1586(.a(s_148), .O(gate278inter3));
  inv1  gate1587(.a(s_149), .O(gate278inter4));
  nand2 gate1588(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1589(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1590(.a(G776), .O(gate278inter7));
  inv1  gate1591(.a(G800), .O(gate278inter8));
  nand2 gate1592(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1593(.a(s_149), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1594(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1595(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1596(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1723(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1724(.a(gate280inter0), .b(s_168), .O(gate280inter1));
  and2  gate1725(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1726(.a(s_168), .O(gate280inter3));
  inv1  gate1727(.a(s_169), .O(gate280inter4));
  nand2 gate1728(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1729(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1730(.a(G779), .O(gate280inter7));
  inv1  gate1731(.a(G803), .O(gate280inter8));
  nand2 gate1732(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1733(.a(s_169), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1734(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1735(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1736(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1387(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1388(.a(gate284inter0), .b(s_120), .O(gate284inter1));
  and2  gate1389(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1390(.a(s_120), .O(gate284inter3));
  inv1  gate1391(.a(s_121), .O(gate284inter4));
  nand2 gate1392(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1393(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1394(.a(G785), .O(gate284inter7));
  inv1  gate1395(.a(G809), .O(gate284inter8));
  nand2 gate1396(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1397(.a(s_121), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1398(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1399(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1400(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2003(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2004(.a(gate287inter0), .b(s_208), .O(gate287inter1));
  and2  gate2005(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2006(.a(s_208), .O(gate287inter3));
  inv1  gate2007(.a(s_209), .O(gate287inter4));
  nand2 gate2008(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2009(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2010(.a(G663), .O(gate287inter7));
  inv1  gate2011(.a(G815), .O(gate287inter8));
  nand2 gate2012(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2013(.a(s_209), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2014(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2015(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2016(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate799(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate800(.a(gate288inter0), .b(s_36), .O(gate288inter1));
  and2  gate801(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate802(.a(s_36), .O(gate288inter3));
  inv1  gate803(.a(s_37), .O(gate288inter4));
  nand2 gate804(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate805(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate806(.a(G791), .O(gate288inter7));
  inv1  gate807(.a(G815), .O(gate288inter8));
  nand2 gate808(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate809(.a(s_37), .b(gate288inter3), .O(gate288inter10));
  nor2  gate810(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate811(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate812(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate743(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate744(.a(gate290inter0), .b(s_28), .O(gate290inter1));
  and2  gate745(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate746(.a(s_28), .O(gate290inter3));
  inv1  gate747(.a(s_29), .O(gate290inter4));
  nand2 gate748(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate749(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate750(.a(G820), .O(gate290inter7));
  inv1  gate751(.a(G821), .O(gate290inter8));
  nand2 gate752(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate753(.a(s_29), .b(gate290inter3), .O(gate290inter10));
  nor2  gate754(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate755(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate756(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1163(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1164(.a(gate293inter0), .b(s_88), .O(gate293inter1));
  and2  gate1165(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1166(.a(s_88), .O(gate293inter3));
  inv1  gate1167(.a(s_89), .O(gate293inter4));
  nand2 gate1168(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1169(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1170(.a(G828), .O(gate293inter7));
  inv1  gate1171(.a(G829), .O(gate293inter8));
  nand2 gate1172(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1173(.a(s_89), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1174(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1175(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1176(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1905(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1906(.a(gate294inter0), .b(s_194), .O(gate294inter1));
  and2  gate1907(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1908(.a(s_194), .O(gate294inter3));
  inv1  gate1909(.a(s_195), .O(gate294inter4));
  nand2 gate1910(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1911(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1912(.a(G832), .O(gate294inter7));
  inv1  gate1913(.a(G833), .O(gate294inter8));
  nand2 gate1914(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1915(.a(s_195), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1916(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1917(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1918(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate785(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate786(.a(gate296inter0), .b(s_34), .O(gate296inter1));
  and2  gate787(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate788(.a(s_34), .O(gate296inter3));
  inv1  gate789(.a(s_35), .O(gate296inter4));
  nand2 gate790(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate791(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate792(.a(G826), .O(gate296inter7));
  inv1  gate793(.a(G827), .O(gate296inter8));
  nand2 gate794(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate795(.a(s_35), .b(gate296inter3), .O(gate296inter10));
  nor2  gate796(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate797(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate798(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate771(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate772(.a(gate390inter0), .b(s_32), .O(gate390inter1));
  and2  gate773(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate774(.a(s_32), .O(gate390inter3));
  inv1  gate775(.a(s_33), .O(gate390inter4));
  nand2 gate776(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate777(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate778(.a(G4), .O(gate390inter7));
  inv1  gate779(.a(G1045), .O(gate390inter8));
  nand2 gate780(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate781(.a(s_33), .b(gate390inter3), .O(gate390inter10));
  nor2  gate782(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate783(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate784(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1667(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1668(.a(gate391inter0), .b(s_160), .O(gate391inter1));
  and2  gate1669(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1670(.a(s_160), .O(gate391inter3));
  inv1  gate1671(.a(s_161), .O(gate391inter4));
  nand2 gate1672(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1673(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1674(.a(G5), .O(gate391inter7));
  inv1  gate1675(.a(G1048), .O(gate391inter8));
  nand2 gate1676(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1677(.a(s_161), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1678(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1679(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1680(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate869(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate870(.a(gate392inter0), .b(s_46), .O(gate392inter1));
  and2  gate871(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate872(.a(s_46), .O(gate392inter3));
  inv1  gate873(.a(s_47), .O(gate392inter4));
  nand2 gate874(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate875(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate876(.a(G6), .O(gate392inter7));
  inv1  gate877(.a(G1051), .O(gate392inter8));
  nand2 gate878(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate879(.a(s_47), .b(gate392inter3), .O(gate392inter10));
  nor2  gate880(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate881(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate882(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1527(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1528(.a(gate394inter0), .b(s_140), .O(gate394inter1));
  and2  gate1529(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1530(.a(s_140), .O(gate394inter3));
  inv1  gate1531(.a(s_141), .O(gate394inter4));
  nand2 gate1532(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1533(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1534(.a(G8), .O(gate394inter7));
  inv1  gate1535(.a(G1057), .O(gate394inter8));
  nand2 gate1536(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1537(.a(s_141), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1538(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1539(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1540(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1639(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1640(.a(gate396inter0), .b(s_156), .O(gate396inter1));
  and2  gate1641(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1642(.a(s_156), .O(gate396inter3));
  inv1  gate1643(.a(s_157), .O(gate396inter4));
  nand2 gate1644(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1645(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1646(.a(G10), .O(gate396inter7));
  inv1  gate1647(.a(G1063), .O(gate396inter8));
  nand2 gate1648(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1649(.a(s_157), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1650(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1651(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1652(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1079(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1080(.a(gate400inter0), .b(s_76), .O(gate400inter1));
  and2  gate1081(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1082(.a(s_76), .O(gate400inter3));
  inv1  gate1083(.a(s_77), .O(gate400inter4));
  nand2 gate1084(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1085(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1086(.a(G14), .O(gate400inter7));
  inv1  gate1087(.a(G1075), .O(gate400inter8));
  nand2 gate1088(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1089(.a(s_77), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1090(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1091(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1092(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1107(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1108(.a(gate406inter0), .b(s_80), .O(gate406inter1));
  and2  gate1109(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1110(.a(s_80), .O(gate406inter3));
  inv1  gate1111(.a(s_81), .O(gate406inter4));
  nand2 gate1112(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1113(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1114(.a(G20), .O(gate406inter7));
  inv1  gate1115(.a(G1093), .O(gate406inter8));
  nand2 gate1116(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1117(.a(s_81), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1118(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1119(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1120(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate547(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate548(.a(gate408inter0), .b(s_0), .O(gate408inter1));
  and2  gate549(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate550(.a(s_0), .O(gate408inter3));
  inv1  gate551(.a(s_1), .O(gate408inter4));
  nand2 gate552(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate553(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate554(.a(G22), .O(gate408inter7));
  inv1  gate555(.a(G1099), .O(gate408inter8));
  nand2 gate556(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate557(.a(s_1), .b(gate408inter3), .O(gate408inter10));
  nor2  gate558(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate559(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate560(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate897(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate898(.a(gate413inter0), .b(s_50), .O(gate413inter1));
  and2  gate899(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate900(.a(s_50), .O(gate413inter3));
  inv1  gate901(.a(s_51), .O(gate413inter4));
  nand2 gate902(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate903(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate904(.a(G27), .O(gate413inter7));
  inv1  gate905(.a(G1114), .O(gate413inter8));
  nand2 gate906(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate907(.a(s_51), .b(gate413inter3), .O(gate413inter10));
  nor2  gate908(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate909(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate910(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate631(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate632(.a(gate416inter0), .b(s_12), .O(gate416inter1));
  and2  gate633(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate634(.a(s_12), .O(gate416inter3));
  inv1  gate635(.a(s_13), .O(gate416inter4));
  nand2 gate636(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate637(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate638(.a(G30), .O(gate416inter7));
  inv1  gate639(.a(G1123), .O(gate416inter8));
  nand2 gate640(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate641(.a(s_13), .b(gate416inter3), .O(gate416inter10));
  nor2  gate642(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate643(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate644(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1821(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1822(.a(gate419inter0), .b(s_182), .O(gate419inter1));
  and2  gate1823(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1824(.a(s_182), .O(gate419inter3));
  inv1  gate1825(.a(s_183), .O(gate419inter4));
  nand2 gate1826(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1827(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1828(.a(G1), .O(gate419inter7));
  inv1  gate1829(.a(G1132), .O(gate419inter8));
  nand2 gate1830(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1831(.a(s_183), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1832(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1833(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1834(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2577(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2578(.a(gate430inter0), .b(s_290), .O(gate430inter1));
  and2  gate2579(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2580(.a(s_290), .O(gate430inter3));
  inv1  gate2581(.a(s_291), .O(gate430inter4));
  nand2 gate2582(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2583(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2584(.a(G1051), .O(gate430inter7));
  inv1  gate2585(.a(G1147), .O(gate430inter8));
  nand2 gate2586(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2587(.a(s_291), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2588(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2589(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2590(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2129(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2130(.a(gate434inter0), .b(s_226), .O(gate434inter1));
  and2  gate2131(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2132(.a(s_226), .O(gate434inter3));
  inv1  gate2133(.a(s_227), .O(gate434inter4));
  nand2 gate2134(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2135(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2136(.a(G1057), .O(gate434inter7));
  inv1  gate2137(.a(G1153), .O(gate434inter8));
  nand2 gate2138(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2139(.a(s_227), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2140(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2141(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2142(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1597(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1598(.a(gate437inter0), .b(s_150), .O(gate437inter1));
  and2  gate1599(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1600(.a(s_150), .O(gate437inter3));
  inv1  gate1601(.a(s_151), .O(gate437inter4));
  nand2 gate1602(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1603(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1604(.a(G10), .O(gate437inter7));
  inv1  gate1605(.a(G1159), .O(gate437inter8));
  nand2 gate1606(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1607(.a(s_151), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1608(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1609(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1610(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2409(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2410(.a(gate439inter0), .b(s_266), .O(gate439inter1));
  and2  gate2411(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2412(.a(s_266), .O(gate439inter3));
  inv1  gate2413(.a(s_267), .O(gate439inter4));
  nand2 gate2414(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2415(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2416(.a(G11), .O(gate439inter7));
  inv1  gate2417(.a(G1162), .O(gate439inter8));
  nand2 gate2418(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2419(.a(s_267), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2420(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2421(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2422(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate603(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate604(.a(gate441inter0), .b(s_8), .O(gate441inter1));
  and2  gate605(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate606(.a(s_8), .O(gate441inter3));
  inv1  gate607(.a(s_9), .O(gate441inter4));
  nand2 gate608(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate609(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate610(.a(G12), .O(gate441inter7));
  inv1  gate611(.a(G1165), .O(gate441inter8));
  nand2 gate612(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate613(.a(s_9), .b(gate441inter3), .O(gate441inter10));
  nor2  gate614(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate615(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate616(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2647(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2648(.a(gate443inter0), .b(s_300), .O(gate443inter1));
  and2  gate2649(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2650(.a(s_300), .O(gate443inter3));
  inv1  gate2651(.a(s_301), .O(gate443inter4));
  nand2 gate2652(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2653(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2654(.a(G13), .O(gate443inter7));
  inv1  gate2655(.a(G1168), .O(gate443inter8));
  nand2 gate2656(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2657(.a(s_301), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2658(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2659(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2660(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2255(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2256(.a(gate444inter0), .b(s_244), .O(gate444inter1));
  and2  gate2257(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2258(.a(s_244), .O(gate444inter3));
  inv1  gate2259(.a(s_245), .O(gate444inter4));
  nand2 gate2260(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2261(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2262(.a(G1072), .O(gate444inter7));
  inv1  gate2263(.a(G1168), .O(gate444inter8));
  nand2 gate2264(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2265(.a(s_245), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2266(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2267(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2268(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1485(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1486(.a(gate445inter0), .b(s_134), .O(gate445inter1));
  and2  gate1487(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1488(.a(s_134), .O(gate445inter3));
  inv1  gate1489(.a(s_135), .O(gate445inter4));
  nand2 gate1490(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1491(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1492(.a(G14), .O(gate445inter7));
  inv1  gate1493(.a(G1171), .O(gate445inter8));
  nand2 gate1494(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1495(.a(s_135), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1496(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1497(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1498(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate2059(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2060(.a(gate446inter0), .b(s_216), .O(gate446inter1));
  and2  gate2061(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2062(.a(s_216), .O(gate446inter3));
  inv1  gate2063(.a(s_217), .O(gate446inter4));
  nand2 gate2064(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2065(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2066(.a(G1075), .O(gate446inter7));
  inv1  gate2067(.a(G1171), .O(gate446inter8));
  nand2 gate2068(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2069(.a(s_217), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2070(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2071(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2072(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1331(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1332(.a(gate447inter0), .b(s_112), .O(gate447inter1));
  and2  gate1333(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1334(.a(s_112), .O(gate447inter3));
  inv1  gate1335(.a(s_113), .O(gate447inter4));
  nand2 gate1336(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1337(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1338(.a(G15), .O(gate447inter7));
  inv1  gate1339(.a(G1174), .O(gate447inter8));
  nand2 gate1340(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1341(.a(s_113), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1342(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1343(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1344(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1751(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1752(.a(gate448inter0), .b(s_172), .O(gate448inter1));
  and2  gate1753(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1754(.a(s_172), .O(gate448inter3));
  inv1  gate1755(.a(s_173), .O(gate448inter4));
  nand2 gate1756(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1757(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1758(.a(G1078), .O(gate448inter7));
  inv1  gate1759(.a(G1174), .O(gate448inter8));
  nand2 gate1760(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1761(.a(s_173), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1762(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1763(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1764(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2283(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2284(.a(gate450inter0), .b(s_248), .O(gate450inter1));
  and2  gate2285(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2286(.a(s_248), .O(gate450inter3));
  inv1  gate2287(.a(s_249), .O(gate450inter4));
  nand2 gate2288(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2289(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2290(.a(G1081), .O(gate450inter7));
  inv1  gate2291(.a(G1177), .O(gate450inter8));
  nand2 gate2292(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2293(.a(s_249), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2294(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2295(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2296(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2017(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2018(.a(gate451inter0), .b(s_210), .O(gate451inter1));
  and2  gate2019(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2020(.a(s_210), .O(gate451inter3));
  inv1  gate2021(.a(s_211), .O(gate451inter4));
  nand2 gate2022(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2023(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2024(.a(G17), .O(gate451inter7));
  inv1  gate2025(.a(G1180), .O(gate451inter8));
  nand2 gate2026(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2027(.a(s_211), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2028(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2029(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2030(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1135(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1136(.a(gate452inter0), .b(s_84), .O(gate452inter1));
  and2  gate1137(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1138(.a(s_84), .O(gate452inter3));
  inv1  gate1139(.a(s_85), .O(gate452inter4));
  nand2 gate1140(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1141(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1142(.a(G1084), .O(gate452inter7));
  inv1  gate1143(.a(G1180), .O(gate452inter8));
  nand2 gate1144(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1145(.a(s_85), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1146(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1147(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1148(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate1513(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1514(.a(gate453inter0), .b(s_138), .O(gate453inter1));
  and2  gate1515(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1516(.a(s_138), .O(gate453inter3));
  inv1  gate1517(.a(s_139), .O(gate453inter4));
  nand2 gate1518(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1519(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1520(.a(G18), .O(gate453inter7));
  inv1  gate1521(.a(G1183), .O(gate453inter8));
  nand2 gate1522(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1523(.a(s_139), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1524(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1525(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1526(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1695(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1696(.a(gate454inter0), .b(s_164), .O(gate454inter1));
  and2  gate1697(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1698(.a(s_164), .O(gate454inter3));
  inv1  gate1699(.a(s_165), .O(gate454inter4));
  nand2 gate1700(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1701(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1702(.a(G1087), .O(gate454inter7));
  inv1  gate1703(.a(G1183), .O(gate454inter8));
  nand2 gate1704(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1705(.a(s_165), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1706(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1707(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1708(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1863(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1864(.a(gate456inter0), .b(s_188), .O(gate456inter1));
  and2  gate1865(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1866(.a(s_188), .O(gate456inter3));
  inv1  gate1867(.a(s_189), .O(gate456inter4));
  nand2 gate1868(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1869(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1870(.a(G1090), .O(gate456inter7));
  inv1  gate1871(.a(G1186), .O(gate456inter8));
  nand2 gate1872(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1873(.a(s_189), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1874(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1875(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1876(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate967(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate968(.a(gate457inter0), .b(s_60), .O(gate457inter1));
  and2  gate969(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate970(.a(s_60), .O(gate457inter3));
  inv1  gate971(.a(s_61), .O(gate457inter4));
  nand2 gate972(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate973(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate974(.a(G20), .O(gate457inter7));
  inv1  gate975(.a(G1189), .O(gate457inter8));
  nand2 gate976(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate977(.a(s_61), .b(gate457inter3), .O(gate457inter10));
  nor2  gate978(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate979(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate980(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1359(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1360(.a(gate459inter0), .b(s_116), .O(gate459inter1));
  and2  gate1361(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1362(.a(s_116), .O(gate459inter3));
  inv1  gate1363(.a(s_117), .O(gate459inter4));
  nand2 gate1364(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1365(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1366(.a(G21), .O(gate459inter7));
  inv1  gate1367(.a(G1192), .O(gate459inter8));
  nand2 gate1368(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1369(.a(s_117), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1370(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1371(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1372(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate925(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate926(.a(gate462inter0), .b(s_54), .O(gate462inter1));
  and2  gate927(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate928(.a(s_54), .O(gate462inter3));
  inv1  gate929(.a(s_55), .O(gate462inter4));
  nand2 gate930(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate931(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate932(.a(G1099), .O(gate462inter7));
  inv1  gate933(.a(G1195), .O(gate462inter8));
  nand2 gate934(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate935(.a(s_55), .b(gate462inter3), .O(gate462inter10));
  nor2  gate936(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate937(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate938(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1429(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1430(.a(gate465inter0), .b(s_126), .O(gate465inter1));
  and2  gate1431(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1432(.a(s_126), .O(gate465inter3));
  inv1  gate1433(.a(s_127), .O(gate465inter4));
  nand2 gate1434(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1435(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1436(.a(G24), .O(gate465inter7));
  inv1  gate1437(.a(G1201), .O(gate465inter8));
  nand2 gate1438(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1439(.a(s_127), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1440(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1441(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1442(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate701(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate702(.a(gate467inter0), .b(s_22), .O(gate467inter1));
  and2  gate703(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate704(.a(s_22), .O(gate467inter3));
  inv1  gate705(.a(s_23), .O(gate467inter4));
  nand2 gate706(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate707(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate708(.a(G25), .O(gate467inter7));
  inv1  gate709(.a(G1204), .O(gate467inter8));
  nand2 gate710(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate711(.a(s_23), .b(gate467inter3), .O(gate467inter10));
  nor2  gate712(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate713(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate714(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate2437(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2438(.a(gate468inter0), .b(s_270), .O(gate468inter1));
  and2  gate2439(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2440(.a(s_270), .O(gate468inter3));
  inv1  gate2441(.a(s_271), .O(gate468inter4));
  nand2 gate2442(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2443(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2444(.a(G1108), .O(gate468inter7));
  inv1  gate2445(.a(G1204), .O(gate468inter8));
  nand2 gate2446(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2447(.a(s_271), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2448(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2449(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2450(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2297(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2298(.a(gate470inter0), .b(s_250), .O(gate470inter1));
  and2  gate2299(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2300(.a(s_250), .O(gate470inter3));
  inv1  gate2301(.a(s_251), .O(gate470inter4));
  nand2 gate2302(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2303(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2304(.a(G1111), .O(gate470inter7));
  inv1  gate2305(.a(G1207), .O(gate470inter8));
  nand2 gate2306(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2307(.a(s_251), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2308(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2309(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2310(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate715(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate716(.a(gate471inter0), .b(s_24), .O(gate471inter1));
  and2  gate717(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate718(.a(s_24), .O(gate471inter3));
  inv1  gate719(.a(s_25), .O(gate471inter4));
  nand2 gate720(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate721(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate722(.a(G27), .O(gate471inter7));
  inv1  gate723(.a(G1210), .O(gate471inter8));
  nand2 gate724(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate725(.a(s_25), .b(gate471inter3), .O(gate471inter10));
  nor2  gate726(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate727(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate728(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2395(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2396(.a(gate472inter0), .b(s_264), .O(gate472inter1));
  and2  gate2397(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2398(.a(s_264), .O(gate472inter3));
  inv1  gate2399(.a(s_265), .O(gate472inter4));
  nand2 gate2400(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2401(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2402(.a(G1114), .O(gate472inter7));
  inv1  gate2403(.a(G1210), .O(gate472inter8));
  nand2 gate2404(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2405(.a(s_265), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2406(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2407(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2408(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2633(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2634(.a(gate475inter0), .b(s_298), .O(gate475inter1));
  and2  gate2635(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2636(.a(s_298), .O(gate475inter3));
  inv1  gate2637(.a(s_299), .O(gate475inter4));
  nand2 gate2638(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2639(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2640(.a(G29), .O(gate475inter7));
  inv1  gate2641(.a(G1216), .O(gate475inter8));
  nand2 gate2642(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2643(.a(s_299), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2644(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2645(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2646(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2591(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2592(.a(gate478inter0), .b(s_292), .O(gate478inter1));
  and2  gate2593(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2594(.a(s_292), .O(gate478inter3));
  inv1  gate2595(.a(s_293), .O(gate478inter4));
  nand2 gate2596(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2597(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2598(.a(G1123), .O(gate478inter7));
  inv1  gate2599(.a(G1219), .O(gate478inter8));
  nand2 gate2600(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2601(.a(s_293), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2602(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2603(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2604(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1261(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1262(.a(gate479inter0), .b(s_102), .O(gate479inter1));
  and2  gate1263(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1264(.a(s_102), .O(gate479inter3));
  inv1  gate1265(.a(s_103), .O(gate479inter4));
  nand2 gate1266(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1267(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1268(.a(G31), .O(gate479inter7));
  inv1  gate1269(.a(G1222), .O(gate479inter8));
  nand2 gate1270(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1271(.a(s_103), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1272(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1273(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1274(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1947(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1948(.a(gate482inter0), .b(s_200), .O(gate482inter1));
  and2  gate1949(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1950(.a(s_200), .O(gate482inter3));
  inv1  gate1951(.a(s_201), .O(gate482inter4));
  nand2 gate1952(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1953(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1954(.a(G1129), .O(gate482inter7));
  inv1  gate1955(.a(G1225), .O(gate482inter8));
  nand2 gate1956(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1957(.a(s_201), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1958(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1959(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1960(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1849(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1850(.a(gate486inter0), .b(s_186), .O(gate486inter1));
  and2  gate1851(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1852(.a(s_186), .O(gate486inter3));
  inv1  gate1853(.a(s_187), .O(gate486inter4));
  nand2 gate1854(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1855(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1856(.a(G1234), .O(gate486inter7));
  inv1  gate1857(.a(G1235), .O(gate486inter8));
  nand2 gate1858(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1859(.a(s_187), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1860(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1861(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1862(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate981(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate982(.a(gate489inter0), .b(s_62), .O(gate489inter1));
  and2  gate983(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate984(.a(s_62), .O(gate489inter3));
  inv1  gate985(.a(s_63), .O(gate489inter4));
  nand2 gate986(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate987(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate988(.a(G1240), .O(gate489inter7));
  inv1  gate989(.a(G1241), .O(gate489inter8));
  nand2 gate990(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate991(.a(s_63), .b(gate489inter3), .O(gate489inter10));
  nor2  gate992(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate993(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate994(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1709(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1710(.a(gate496inter0), .b(s_166), .O(gate496inter1));
  and2  gate1711(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1712(.a(s_166), .O(gate496inter3));
  inv1  gate1713(.a(s_167), .O(gate496inter4));
  nand2 gate1714(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1715(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1716(.a(G1254), .O(gate496inter7));
  inv1  gate1717(.a(G1255), .O(gate496inter8));
  nand2 gate1718(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1719(.a(s_167), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1720(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1721(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1722(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1065(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1066(.a(gate499inter0), .b(s_74), .O(gate499inter1));
  and2  gate1067(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1068(.a(s_74), .O(gate499inter3));
  inv1  gate1069(.a(s_75), .O(gate499inter4));
  nand2 gate1070(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1071(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1072(.a(G1260), .O(gate499inter7));
  inv1  gate1073(.a(G1261), .O(gate499inter8));
  nand2 gate1074(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1075(.a(s_75), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1076(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1077(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1078(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate841(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate842(.a(gate503inter0), .b(s_42), .O(gate503inter1));
  and2  gate843(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate844(.a(s_42), .O(gate503inter3));
  inv1  gate845(.a(s_43), .O(gate503inter4));
  nand2 gate846(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate847(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate848(.a(G1268), .O(gate503inter7));
  inv1  gate849(.a(G1269), .O(gate503inter8));
  nand2 gate850(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate851(.a(s_43), .b(gate503inter3), .O(gate503inter10));
  nor2  gate852(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate853(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate854(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1289(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1290(.a(gate504inter0), .b(s_106), .O(gate504inter1));
  and2  gate1291(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1292(.a(s_106), .O(gate504inter3));
  inv1  gate1293(.a(s_107), .O(gate504inter4));
  nand2 gate1294(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1295(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1296(.a(G1270), .O(gate504inter7));
  inv1  gate1297(.a(G1271), .O(gate504inter8));
  nand2 gate1298(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1299(.a(s_107), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1300(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1301(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1302(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1457(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1458(.a(gate505inter0), .b(s_130), .O(gate505inter1));
  and2  gate1459(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1460(.a(s_130), .O(gate505inter3));
  inv1  gate1461(.a(s_131), .O(gate505inter4));
  nand2 gate1462(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1463(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1464(.a(G1272), .O(gate505inter7));
  inv1  gate1465(.a(G1273), .O(gate505inter8));
  nand2 gate1466(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1467(.a(s_131), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1468(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1469(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1470(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule