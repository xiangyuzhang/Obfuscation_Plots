module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1149(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1150(.a(gate28inter0), .b(s_86), .O(gate28inter1));
  and2  gate1151(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1152(.a(s_86), .O(gate28inter3));
  inv1  gate1153(.a(s_87), .O(gate28inter4));
  nand2 gate1154(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1155(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1156(.a(G10), .O(gate28inter7));
  inv1  gate1157(.a(G14), .O(gate28inter8));
  nand2 gate1158(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1159(.a(s_87), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1160(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1161(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1162(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate911(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate912(.a(gate41inter0), .b(s_52), .O(gate41inter1));
  and2  gate913(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate914(.a(s_52), .O(gate41inter3));
  inv1  gate915(.a(s_53), .O(gate41inter4));
  nand2 gate916(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate917(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate918(.a(G1), .O(gate41inter7));
  inv1  gate919(.a(G266), .O(gate41inter8));
  nand2 gate920(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate921(.a(s_53), .b(gate41inter3), .O(gate41inter10));
  nor2  gate922(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate923(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate924(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate925(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate926(.a(gate44inter0), .b(s_54), .O(gate44inter1));
  and2  gate927(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate928(.a(s_54), .O(gate44inter3));
  inv1  gate929(.a(s_55), .O(gate44inter4));
  nand2 gate930(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate931(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate932(.a(G4), .O(gate44inter7));
  inv1  gate933(.a(G269), .O(gate44inter8));
  nand2 gate934(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate935(.a(s_55), .b(gate44inter3), .O(gate44inter10));
  nor2  gate936(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate937(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate938(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate939(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate940(.a(gate45inter0), .b(s_56), .O(gate45inter1));
  and2  gate941(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate942(.a(s_56), .O(gate45inter3));
  inv1  gate943(.a(s_57), .O(gate45inter4));
  nand2 gate944(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate945(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate946(.a(G5), .O(gate45inter7));
  inv1  gate947(.a(G272), .O(gate45inter8));
  nand2 gate948(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate949(.a(s_57), .b(gate45inter3), .O(gate45inter10));
  nor2  gate950(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate951(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate952(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1121(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1122(.a(gate48inter0), .b(s_82), .O(gate48inter1));
  and2  gate1123(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1124(.a(s_82), .O(gate48inter3));
  inv1  gate1125(.a(s_83), .O(gate48inter4));
  nand2 gate1126(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1127(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1128(.a(G8), .O(gate48inter7));
  inv1  gate1129(.a(G275), .O(gate48inter8));
  nand2 gate1130(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1131(.a(s_83), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1132(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1133(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1134(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1079(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1080(.a(gate52inter0), .b(s_76), .O(gate52inter1));
  and2  gate1081(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1082(.a(s_76), .O(gate52inter3));
  inv1  gate1083(.a(s_77), .O(gate52inter4));
  nand2 gate1084(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1085(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1086(.a(G12), .O(gate52inter7));
  inv1  gate1087(.a(G281), .O(gate52inter8));
  nand2 gate1088(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1089(.a(s_77), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1090(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1091(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1092(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate757(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate758(.a(gate55inter0), .b(s_30), .O(gate55inter1));
  and2  gate759(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate760(.a(s_30), .O(gate55inter3));
  inv1  gate761(.a(s_31), .O(gate55inter4));
  nand2 gate762(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate763(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate764(.a(G15), .O(gate55inter7));
  inv1  gate765(.a(G287), .O(gate55inter8));
  nand2 gate766(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate767(.a(s_31), .b(gate55inter3), .O(gate55inter10));
  nor2  gate768(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate769(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate770(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate981(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate982(.a(gate66inter0), .b(s_62), .O(gate66inter1));
  and2  gate983(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate984(.a(s_62), .O(gate66inter3));
  inv1  gate985(.a(s_63), .O(gate66inter4));
  nand2 gate986(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate987(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate988(.a(G26), .O(gate66inter7));
  inv1  gate989(.a(G302), .O(gate66inter8));
  nand2 gate990(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate991(.a(s_63), .b(gate66inter3), .O(gate66inter10));
  nor2  gate992(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate993(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate994(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate995(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate996(.a(gate86inter0), .b(s_64), .O(gate86inter1));
  and2  gate997(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate998(.a(s_64), .O(gate86inter3));
  inv1  gate999(.a(s_65), .O(gate86inter4));
  nand2 gate1000(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1001(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1002(.a(G8), .O(gate86inter7));
  inv1  gate1003(.a(G332), .O(gate86inter8));
  nand2 gate1004(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1005(.a(s_65), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1006(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1007(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1008(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate869(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate870(.a(gate109inter0), .b(s_46), .O(gate109inter1));
  and2  gate871(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate872(.a(s_46), .O(gate109inter3));
  inv1  gate873(.a(s_47), .O(gate109inter4));
  nand2 gate874(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate875(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate876(.a(G370), .O(gate109inter7));
  inv1  gate877(.a(G371), .O(gate109inter8));
  nand2 gate878(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate879(.a(s_47), .b(gate109inter3), .O(gate109inter10));
  nor2  gate880(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate881(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate882(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate617(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate618(.a(gate119inter0), .b(s_10), .O(gate119inter1));
  and2  gate619(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate620(.a(s_10), .O(gate119inter3));
  inv1  gate621(.a(s_11), .O(gate119inter4));
  nand2 gate622(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate623(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate624(.a(G390), .O(gate119inter7));
  inv1  gate625(.a(G391), .O(gate119inter8));
  nand2 gate626(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate627(.a(s_11), .b(gate119inter3), .O(gate119inter10));
  nor2  gate628(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate629(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate630(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate561(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate562(.a(gate136inter0), .b(s_2), .O(gate136inter1));
  and2  gate563(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate564(.a(s_2), .O(gate136inter3));
  inv1  gate565(.a(s_3), .O(gate136inter4));
  nand2 gate566(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate567(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate568(.a(G424), .O(gate136inter7));
  inv1  gate569(.a(G425), .O(gate136inter8));
  nand2 gate570(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate571(.a(s_3), .b(gate136inter3), .O(gate136inter10));
  nor2  gate572(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate573(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate574(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1009(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1010(.a(gate148inter0), .b(s_66), .O(gate148inter1));
  and2  gate1011(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1012(.a(s_66), .O(gate148inter3));
  inv1  gate1013(.a(s_67), .O(gate148inter4));
  nand2 gate1014(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1015(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1016(.a(G492), .O(gate148inter7));
  inv1  gate1017(.a(G495), .O(gate148inter8));
  nand2 gate1018(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1019(.a(s_67), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1020(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1021(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1022(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate575(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate576(.a(gate149inter0), .b(s_4), .O(gate149inter1));
  and2  gate577(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate578(.a(s_4), .O(gate149inter3));
  inv1  gate579(.a(s_5), .O(gate149inter4));
  nand2 gate580(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate581(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate582(.a(G498), .O(gate149inter7));
  inv1  gate583(.a(G501), .O(gate149inter8));
  nand2 gate584(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate585(.a(s_5), .b(gate149inter3), .O(gate149inter10));
  nor2  gate586(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate587(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate588(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate659(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate660(.a(gate158inter0), .b(s_16), .O(gate158inter1));
  and2  gate661(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate662(.a(s_16), .O(gate158inter3));
  inv1  gate663(.a(s_17), .O(gate158inter4));
  nand2 gate664(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate665(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate666(.a(G441), .O(gate158inter7));
  inv1  gate667(.a(G528), .O(gate158inter8));
  nand2 gate668(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate669(.a(s_17), .b(gate158inter3), .O(gate158inter10));
  nor2  gate670(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate671(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate672(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate743(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate744(.a(gate161inter0), .b(s_28), .O(gate161inter1));
  and2  gate745(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate746(.a(s_28), .O(gate161inter3));
  inv1  gate747(.a(s_29), .O(gate161inter4));
  nand2 gate748(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate749(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate750(.a(G450), .O(gate161inter7));
  inv1  gate751(.a(G534), .O(gate161inter8));
  nand2 gate752(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate753(.a(s_29), .b(gate161inter3), .O(gate161inter10));
  nor2  gate754(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate755(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate756(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate953(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate954(.a(gate162inter0), .b(s_58), .O(gate162inter1));
  and2  gate955(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate956(.a(s_58), .O(gate162inter3));
  inv1  gate957(.a(s_59), .O(gate162inter4));
  nand2 gate958(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate959(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate960(.a(G453), .O(gate162inter7));
  inv1  gate961(.a(G534), .O(gate162inter8));
  nand2 gate962(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate963(.a(s_59), .b(gate162inter3), .O(gate162inter10));
  nor2  gate964(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate965(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate966(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1219(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1220(.a(gate169inter0), .b(s_96), .O(gate169inter1));
  and2  gate1221(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1222(.a(s_96), .O(gate169inter3));
  inv1  gate1223(.a(s_97), .O(gate169inter4));
  nand2 gate1224(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1225(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1226(.a(G474), .O(gate169inter7));
  inv1  gate1227(.a(G546), .O(gate169inter8));
  nand2 gate1228(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1229(.a(s_97), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1230(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1231(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1232(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate729(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate730(.a(gate172inter0), .b(s_26), .O(gate172inter1));
  and2  gate731(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate732(.a(s_26), .O(gate172inter3));
  inv1  gate733(.a(s_27), .O(gate172inter4));
  nand2 gate734(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate735(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate736(.a(G483), .O(gate172inter7));
  inv1  gate737(.a(G549), .O(gate172inter8));
  nand2 gate738(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate739(.a(s_27), .b(gate172inter3), .O(gate172inter10));
  nor2  gate740(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate741(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate742(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1093(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1094(.a(gate186inter0), .b(s_78), .O(gate186inter1));
  and2  gate1095(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1096(.a(s_78), .O(gate186inter3));
  inv1  gate1097(.a(s_79), .O(gate186inter4));
  nand2 gate1098(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1099(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1100(.a(G572), .O(gate186inter7));
  inv1  gate1101(.a(G573), .O(gate186inter8));
  nand2 gate1102(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1103(.a(s_79), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1104(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1105(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1106(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1247(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1248(.a(gate195inter0), .b(s_100), .O(gate195inter1));
  and2  gate1249(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1250(.a(s_100), .O(gate195inter3));
  inv1  gate1251(.a(s_101), .O(gate195inter4));
  nand2 gate1252(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1253(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1254(.a(G590), .O(gate195inter7));
  inv1  gate1255(.a(G591), .O(gate195inter8));
  nand2 gate1256(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1257(.a(s_101), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1258(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1259(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1260(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate547(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate548(.a(gate203inter0), .b(s_0), .O(gate203inter1));
  and2  gate549(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate550(.a(s_0), .O(gate203inter3));
  inv1  gate551(.a(s_1), .O(gate203inter4));
  nand2 gate552(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate553(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate554(.a(G602), .O(gate203inter7));
  inv1  gate555(.a(G612), .O(gate203inter8));
  nand2 gate556(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate557(.a(s_1), .b(gate203inter3), .O(gate203inter10));
  nor2  gate558(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate559(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate560(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1023(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1024(.a(gate209inter0), .b(s_68), .O(gate209inter1));
  and2  gate1025(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1026(.a(s_68), .O(gate209inter3));
  inv1  gate1027(.a(s_69), .O(gate209inter4));
  nand2 gate1028(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1029(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1030(.a(G602), .O(gate209inter7));
  inv1  gate1031(.a(G666), .O(gate209inter8));
  nand2 gate1032(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1033(.a(s_69), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1034(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1035(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1036(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1135(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1136(.a(gate220inter0), .b(s_84), .O(gate220inter1));
  and2  gate1137(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1138(.a(s_84), .O(gate220inter3));
  inv1  gate1139(.a(s_85), .O(gate220inter4));
  nand2 gate1140(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1141(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1142(.a(G637), .O(gate220inter7));
  inv1  gate1143(.a(G681), .O(gate220inter8));
  nand2 gate1144(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1145(.a(s_85), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1146(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1147(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1148(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate883(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate884(.a(gate230inter0), .b(s_48), .O(gate230inter1));
  and2  gate885(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate886(.a(s_48), .O(gate230inter3));
  inv1  gate887(.a(s_49), .O(gate230inter4));
  nand2 gate888(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate889(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate890(.a(G700), .O(gate230inter7));
  inv1  gate891(.a(G701), .O(gate230inter8));
  nand2 gate892(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate893(.a(s_49), .b(gate230inter3), .O(gate230inter10));
  nor2  gate894(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate895(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate896(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1065(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1066(.a(gate231inter0), .b(s_74), .O(gate231inter1));
  and2  gate1067(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1068(.a(s_74), .O(gate231inter3));
  inv1  gate1069(.a(s_75), .O(gate231inter4));
  nand2 gate1070(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1071(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1072(.a(G702), .O(gate231inter7));
  inv1  gate1073(.a(G703), .O(gate231inter8));
  nand2 gate1074(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1075(.a(s_75), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1076(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1077(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1078(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate813(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate814(.a(gate237inter0), .b(s_38), .O(gate237inter1));
  and2  gate815(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate816(.a(s_38), .O(gate237inter3));
  inv1  gate817(.a(s_39), .O(gate237inter4));
  nand2 gate818(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate819(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate820(.a(G254), .O(gate237inter7));
  inv1  gate821(.a(G706), .O(gate237inter8));
  nand2 gate822(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate823(.a(s_39), .b(gate237inter3), .O(gate237inter10));
  nor2  gate824(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate825(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate826(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate841(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate842(.a(gate239inter0), .b(s_42), .O(gate239inter1));
  and2  gate843(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate844(.a(s_42), .O(gate239inter3));
  inv1  gate845(.a(s_43), .O(gate239inter4));
  nand2 gate846(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate847(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate848(.a(G260), .O(gate239inter7));
  inv1  gate849(.a(G712), .O(gate239inter8));
  nand2 gate850(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate851(.a(s_43), .b(gate239inter3), .O(gate239inter10));
  nor2  gate852(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate853(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate854(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1107(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1108(.a(gate245inter0), .b(s_80), .O(gate245inter1));
  and2  gate1109(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1110(.a(s_80), .O(gate245inter3));
  inv1  gate1111(.a(s_81), .O(gate245inter4));
  nand2 gate1112(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1113(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1114(.a(G248), .O(gate245inter7));
  inv1  gate1115(.a(G736), .O(gate245inter8));
  nand2 gate1116(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1117(.a(s_81), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1118(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1119(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1120(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1163(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1164(.a(gate253inter0), .b(s_88), .O(gate253inter1));
  and2  gate1165(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1166(.a(s_88), .O(gate253inter3));
  inv1  gate1167(.a(s_89), .O(gate253inter4));
  nand2 gate1168(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1169(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1170(.a(G260), .O(gate253inter7));
  inv1  gate1171(.a(G748), .O(gate253inter8));
  nand2 gate1172(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1173(.a(s_89), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1174(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1175(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1176(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1051(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1052(.a(gate256inter0), .b(s_72), .O(gate256inter1));
  and2  gate1053(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1054(.a(s_72), .O(gate256inter3));
  inv1  gate1055(.a(s_73), .O(gate256inter4));
  nand2 gate1056(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1057(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1058(.a(G715), .O(gate256inter7));
  inv1  gate1059(.a(G751), .O(gate256inter8));
  nand2 gate1060(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1061(.a(s_73), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1062(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1063(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1064(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate645(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate646(.a(gate262inter0), .b(s_14), .O(gate262inter1));
  and2  gate647(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate648(.a(s_14), .O(gate262inter3));
  inv1  gate649(.a(s_15), .O(gate262inter4));
  nand2 gate650(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate651(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate652(.a(G764), .O(gate262inter7));
  inv1  gate653(.a(G765), .O(gate262inter8));
  nand2 gate654(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate655(.a(s_15), .b(gate262inter3), .O(gate262inter10));
  nor2  gate656(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate657(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate658(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate799(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate800(.a(gate273inter0), .b(s_36), .O(gate273inter1));
  and2  gate801(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate802(.a(s_36), .O(gate273inter3));
  inv1  gate803(.a(s_37), .O(gate273inter4));
  nand2 gate804(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate805(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate806(.a(G642), .O(gate273inter7));
  inv1  gate807(.a(G794), .O(gate273inter8));
  nand2 gate808(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate809(.a(s_37), .b(gate273inter3), .O(gate273inter10));
  nor2  gate810(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate811(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate812(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate827(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate828(.a(gate276inter0), .b(s_40), .O(gate276inter1));
  and2  gate829(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate830(.a(s_40), .O(gate276inter3));
  inv1  gate831(.a(s_41), .O(gate276inter4));
  nand2 gate832(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate833(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate834(.a(G773), .O(gate276inter7));
  inv1  gate835(.a(G797), .O(gate276inter8));
  nand2 gate836(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate837(.a(s_41), .b(gate276inter3), .O(gate276inter10));
  nor2  gate838(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate839(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate840(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate715(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate716(.a(gate280inter0), .b(s_24), .O(gate280inter1));
  and2  gate717(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate718(.a(s_24), .O(gate280inter3));
  inv1  gate719(.a(s_25), .O(gate280inter4));
  nand2 gate720(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate721(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate722(.a(G779), .O(gate280inter7));
  inv1  gate723(.a(G803), .O(gate280inter8));
  nand2 gate724(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate725(.a(s_25), .b(gate280inter3), .O(gate280inter10));
  nor2  gate726(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate727(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate728(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate771(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate772(.a(gate281inter0), .b(s_32), .O(gate281inter1));
  and2  gate773(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate774(.a(s_32), .O(gate281inter3));
  inv1  gate775(.a(s_33), .O(gate281inter4));
  nand2 gate776(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate777(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate778(.a(G654), .O(gate281inter7));
  inv1  gate779(.a(G806), .O(gate281inter8));
  nand2 gate780(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate781(.a(s_33), .b(gate281inter3), .O(gate281inter10));
  nor2  gate782(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate783(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate784(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1177(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1178(.a(gate288inter0), .b(s_90), .O(gate288inter1));
  and2  gate1179(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1180(.a(s_90), .O(gate288inter3));
  inv1  gate1181(.a(s_91), .O(gate288inter4));
  nand2 gate1182(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1183(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1184(.a(G791), .O(gate288inter7));
  inv1  gate1185(.a(G815), .O(gate288inter8));
  nand2 gate1186(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1187(.a(s_91), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1188(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1189(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1190(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate603(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate604(.a(gate296inter0), .b(s_8), .O(gate296inter1));
  and2  gate605(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate606(.a(s_8), .O(gate296inter3));
  inv1  gate607(.a(s_9), .O(gate296inter4));
  nand2 gate608(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate609(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate610(.a(G826), .O(gate296inter7));
  inv1  gate611(.a(G827), .O(gate296inter8));
  nand2 gate612(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate613(.a(s_9), .b(gate296inter3), .O(gate296inter10));
  nor2  gate614(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate615(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate616(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate589(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate590(.a(gate394inter0), .b(s_6), .O(gate394inter1));
  and2  gate591(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate592(.a(s_6), .O(gate394inter3));
  inv1  gate593(.a(s_7), .O(gate394inter4));
  nand2 gate594(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate595(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate596(.a(G8), .O(gate394inter7));
  inv1  gate597(.a(G1057), .O(gate394inter8));
  nand2 gate598(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate599(.a(s_7), .b(gate394inter3), .O(gate394inter10));
  nor2  gate600(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate601(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate602(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1205(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1206(.a(gate396inter0), .b(s_94), .O(gate396inter1));
  and2  gate1207(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1208(.a(s_94), .O(gate396inter3));
  inv1  gate1209(.a(s_95), .O(gate396inter4));
  nand2 gate1210(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1211(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1212(.a(G10), .O(gate396inter7));
  inv1  gate1213(.a(G1063), .O(gate396inter8));
  nand2 gate1214(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1215(.a(s_95), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1216(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1217(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1218(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate701(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate702(.a(gate415inter0), .b(s_22), .O(gate415inter1));
  and2  gate703(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate704(.a(s_22), .O(gate415inter3));
  inv1  gate705(.a(s_23), .O(gate415inter4));
  nand2 gate706(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate707(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate708(.a(G29), .O(gate415inter7));
  inv1  gate709(.a(G1120), .O(gate415inter8));
  nand2 gate710(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate711(.a(s_23), .b(gate415inter3), .O(gate415inter10));
  nor2  gate712(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate713(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate714(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1191(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1192(.a(gate416inter0), .b(s_92), .O(gate416inter1));
  and2  gate1193(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1194(.a(s_92), .O(gate416inter3));
  inv1  gate1195(.a(s_93), .O(gate416inter4));
  nand2 gate1196(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1197(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1198(.a(G30), .O(gate416inter7));
  inv1  gate1199(.a(G1123), .O(gate416inter8));
  nand2 gate1200(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1201(.a(s_93), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1202(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1203(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1204(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate687(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate688(.a(gate424inter0), .b(s_20), .O(gate424inter1));
  and2  gate689(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate690(.a(s_20), .O(gate424inter3));
  inv1  gate691(.a(s_21), .O(gate424inter4));
  nand2 gate692(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate693(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate694(.a(G1042), .O(gate424inter7));
  inv1  gate695(.a(G1138), .O(gate424inter8));
  nand2 gate696(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate697(.a(s_21), .b(gate424inter3), .O(gate424inter10));
  nor2  gate698(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate699(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate700(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate673(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate674(.a(gate429inter0), .b(s_18), .O(gate429inter1));
  and2  gate675(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate676(.a(s_18), .O(gate429inter3));
  inv1  gate677(.a(s_19), .O(gate429inter4));
  nand2 gate678(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate679(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate680(.a(G6), .O(gate429inter7));
  inv1  gate681(.a(G1147), .O(gate429inter8));
  nand2 gate682(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate683(.a(s_19), .b(gate429inter3), .O(gate429inter10));
  nor2  gate684(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate685(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate686(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate631(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate632(.a(gate446inter0), .b(s_12), .O(gate446inter1));
  and2  gate633(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate634(.a(s_12), .O(gate446inter3));
  inv1  gate635(.a(s_13), .O(gate446inter4));
  nand2 gate636(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate637(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate638(.a(G1075), .O(gate446inter7));
  inv1  gate639(.a(G1171), .O(gate446inter8));
  nand2 gate640(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate641(.a(s_13), .b(gate446inter3), .O(gate446inter10));
  nor2  gate642(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate643(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate644(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1233(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1234(.a(gate447inter0), .b(s_98), .O(gate447inter1));
  and2  gate1235(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1236(.a(s_98), .O(gate447inter3));
  inv1  gate1237(.a(s_99), .O(gate447inter4));
  nand2 gate1238(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1239(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1240(.a(G15), .O(gate447inter7));
  inv1  gate1241(.a(G1174), .O(gate447inter8));
  nand2 gate1242(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1243(.a(s_99), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1244(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1245(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1246(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate785(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate786(.a(gate449inter0), .b(s_34), .O(gate449inter1));
  and2  gate787(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate788(.a(s_34), .O(gate449inter3));
  inv1  gate789(.a(s_35), .O(gate449inter4));
  nand2 gate790(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate791(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate792(.a(G16), .O(gate449inter7));
  inv1  gate793(.a(G1177), .O(gate449inter8));
  nand2 gate794(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate795(.a(s_35), .b(gate449inter3), .O(gate449inter10));
  nor2  gate796(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate797(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate798(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate855(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate856(.a(gate463inter0), .b(s_44), .O(gate463inter1));
  and2  gate857(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate858(.a(s_44), .O(gate463inter3));
  inv1  gate859(.a(s_45), .O(gate463inter4));
  nand2 gate860(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate861(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate862(.a(G23), .O(gate463inter7));
  inv1  gate863(.a(G1198), .O(gate463inter8));
  nand2 gate864(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate865(.a(s_45), .b(gate463inter3), .O(gate463inter10));
  nor2  gate866(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate867(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate868(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate897(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate898(.a(gate476inter0), .b(s_50), .O(gate476inter1));
  and2  gate899(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate900(.a(s_50), .O(gate476inter3));
  inv1  gate901(.a(s_51), .O(gate476inter4));
  nand2 gate902(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate903(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate904(.a(G1120), .O(gate476inter7));
  inv1  gate905(.a(G1216), .O(gate476inter8));
  nand2 gate906(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate907(.a(s_51), .b(gate476inter3), .O(gate476inter10));
  nor2  gate908(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate909(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate910(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1037(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1038(.a(gate499inter0), .b(s_70), .O(gate499inter1));
  and2  gate1039(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1040(.a(s_70), .O(gate499inter3));
  inv1  gate1041(.a(s_71), .O(gate499inter4));
  nand2 gate1042(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1043(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1044(.a(G1260), .O(gate499inter7));
  inv1  gate1045(.a(G1261), .O(gate499inter8));
  nand2 gate1046(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1047(.a(s_71), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1048(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1049(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1050(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate967(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate968(.a(gate506inter0), .b(s_60), .O(gate506inter1));
  and2  gate969(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate970(.a(s_60), .O(gate506inter3));
  inv1  gate971(.a(s_61), .O(gate506inter4));
  nand2 gate972(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate973(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate974(.a(G1274), .O(gate506inter7));
  inv1  gate975(.a(G1275), .O(gate506inter8));
  nand2 gate976(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate977(.a(s_61), .b(gate506inter3), .O(gate506inter10));
  nor2  gate978(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate979(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate980(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule