module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1877(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1878(.a(gate19inter0), .b(s_190), .O(gate19inter1));
  and2  gate1879(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1880(.a(s_190), .O(gate19inter3));
  inv1  gate1881(.a(s_191), .O(gate19inter4));
  nand2 gate1882(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1883(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1884(.a(G21), .O(gate19inter7));
  inv1  gate1885(.a(G22), .O(gate19inter8));
  nand2 gate1886(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1887(.a(s_191), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1888(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1889(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1890(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1765(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1766(.a(gate21inter0), .b(s_174), .O(gate21inter1));
  and2  gate1767(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1768(.a(s_174), .O(gate21inter3));
  inv1  gate1769(.a(s_175), .O(gate21inter4));
  nand2 gate1770(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1771(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1772(.a(G25), .O(gate21inter7));
  inv1  gate1773(.a(G26), .O(gate21inter8));
  nand2 gate1774(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1775(.a(s_175), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1776(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1777(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1778(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1639(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1640(.a(gate24inter0), .b(s_156), .O(gate24inter1));
  and2  gate1641(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1642(.a(s_156), .O(gate24inter3));
  inv1  gate1643(.a(s_157), .O(gate24inter4));
  nand2 gate1644(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1645(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1646(.a(G31), .O(gate24inter7));
  inv1  gate1647(.a(G32), .O(gate24inter8));
  nand2 gate1648(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1649(.a(s_157), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1650(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1651(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1652(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1051(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1052(.a(gate28inter0), .b(s_72), .O(gate28inter1));
  and2  gate1053(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1054(.a(s_72), .O(gate28inter3));
  inv1  gate1055(.a(s_73), .O(gate28inter4));
  nand2 gate1056(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1057(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1058(.a(G10), .O(gate28inter7));
  inv1  gate1059(.a(G14), .O(gate28inter8));
  nand2 gate1060(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1061(.a(s_73), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1062(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1063(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1064(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1107(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1108(.a(gate37inter0), .b(s_80), .O(gate37inter1));
  and2  gate1109(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1110(.a(s_80), .O(gate37inter3));
  inv1  gate1111(.a(s_81), .O(gate37inter4));
  nand2 gate1112(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1113(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1114(.a(G19), .O(gate37inter7));
  inv1  gate1115(.a(G23), .O(gate37inter8));
  nand2 gate1116(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1117(.a(s_81), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1118(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1119(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1120(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1093(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1094(.a(gate38inter0), .b(s_78), .O(gate38inter1));
  and2  gate1095(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1096(.a(s_78), .O(gate38inter3));
  inv1  gate1097(.a(s_79), .O(gate38inter4));
  nand2 gate1098(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1099(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1100(.a(G27), .O(gate38inter7));
  inv1  gate1101(.a(G31), .O(gate38inter8));
  nand2 gate1102(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1103(.a(s_79), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1104(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1105(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1106(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate729(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate730(.a(gate41inter0), .b(s_26), .O(gate41inter1));
  and2  gate731(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate732(.a(s_26), .O(gate41inter3));
  inv1  gate733(.a(s_27), .O(gate41inter4));
  nand2 gate734(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate735(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate736(.a(G1), .O(gate41inter7));
  inv1  gate737(.a(G266), .O(gate41inter8));
  nand2 gate738(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate739(.a(s_27), .b(gate41inter3), .O(gate41inter10));
  nor2  gate740(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate741(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate742(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate687(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate688(.a(gate44inter0), .b(s_20), .O(gate44inter1));
  and2  gate689(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate690(.a(s_20), .O(gate44inter3));
  inv1  gate691(.a(s_21), .O(gate44inter4));
  nand2 gate692(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate693(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate694(.a(G4), .O(gate44inter7));
  inv1  gate695(.a(G269), .O(gate44inter8));
  nand2 gate696(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate697(.a(s_21), .b(gate44inter3), .O(gate44inter10));
  nor2  gate698(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate699(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate700(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate841(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate842(.a(gate50inter0), .b(s_42), .O(gate50inter1));
  and2  gate843(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate844(.a(s_42), .O(gate50inter3));
  inv1  gate845(.a(s_43), .O(gate50inter4));
  nand2 gate846(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate847(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate848(.a(G10), .O(gate50inter7));
  inv1  gate849(.a(G278), .O(gate50inter8));
  nand2 gate850(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate851(.a(s_43), .b(gate50inter3), .O(gate50inter10));
  nor2  gate852(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate853(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate854(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2171(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2172(.a(gate51inter0), .b(s_232), .O(gate51inter1));
  and2  gate2173(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2174(.a(s_232), .O(gate51inter3));
  inv1  gate2175(.a(s_233), .O(gate51inter4));
  nand2 gate2176(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2177(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2178(.a(G11), .O(gate51inter7));
  inv1  gate2179(.a(G281), .O(gate51inter8));
  nand2 gate2180(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2181(.a(s_233), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2182(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2183(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2184(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1527(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1528(.a(gate54inter0), .b(s_140), .O(gate54inter1));
  and2  gate1529(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1530(.a(s_140), .O(gate54inter3));
  inv1  gate1531(.a(s_141), .O(gate54inter4));
  nand2 gate1532(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1533(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1534(.a(G14), .O(gate54inter7));
  inv1  gate1535(.a(G284), .O(gate54inter8));
  nand2 gate1536(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1537(.a(s_141), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1538(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1539(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1540(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1401(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1402(.a(gate60inter0), .b(s_122), .O(gate60inter1));
  and2  gate1403(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1404(.a(s_122), .O(gate60inter3));
  inv1  gate1405(.a(s_123), .O(gate60inter4));
  nand2 gate1406(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1407(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1408(.a(G20), .O(gate60inter7));
  inv1  gate1409(.a(G293), .O(gate60inter8));
  nand2 gate1410(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1411(.a(s_123), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1412(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1413(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1414(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate673(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate674(.a(gate66inter0), .b(s_18), .O(gate66inter1));
  and2  gate675(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate676(.a(s_18), .O(gate66inter3));
  inv1  gate677(.a(s_19), .O(gate66inter4));
  nand2 gate678(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate679(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate680(.a(G26), .O(gate66inter7));
  inv1  gate681(.a(G302), .O(gate66inter8));
  nand2 gate682(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate683(.a(s_19), .b(gate66inter3), .O(gate66inter10));
  nor2  gate684(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate685(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate686(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1891(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1892(.a(gate70inter0), .b(s_192), .O(gate70inter1));
  and2  gate1893(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1894(.a(s_192), .O(gate70inter3));
  inv1  gate1895(.a(s_193), .O(gate70inter4));
  nand2 gate1896(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1897(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1898(.a(G30), .O(gate70inter7));
  inv1  gate1899(.a(G308), .O(gate70inter8));
  nand2 gate1900(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1901(.a(s_193), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1902(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1903(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1904(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate603(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate604(.a(gate74inter0), .b(s_8), .O(gate74inter1));
  and2  gate605(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate606(.a(s_8), .O(gate74inter3));
  inv1  gate607(.a(s_9), .O(gate74inter4));
  nand2 gate608(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate609(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate610(.a(G5), .O(gate74inter7));
  inv1  gate611(.a(G314), .O(gate74inter8));
  nand2 gate612(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate613(.a(s_9), .b(gate74inter3), .O(gate74inter10));
  nor2  gate614(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate615(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate616(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate883(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate884(.a(gate76inter0), .b(s_48), .O(gate76inter1));
  and2  gate885(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate886(.a(s_48), .O(gate76inter3));
  inv1  gate887(.a(s_49), .O(gate76inter4));
  nand2 gate888(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate889(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate890(.a(G13), .O(gate76inter7));
  inv1  gate891(.a(G317), .O(gate76inter8));
  nand2 gate892(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate893(.a(s_49), .b(gate76inter3), .O(gate76inter10));
  nor2  gate894(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate895(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate896(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2115(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2116(.a(gate81inter0), .b(s_224), .O(gate81inter1));
  and2  gate2117(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2118(.a(s_224), .O(gate81inter3));
  inv1  gate2119(.a(s_225), .O(gate81inter4));
  nand2 gate2120(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2121(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2122(.a(G3), .O(gate81inter7));
  inv1  gate2123(.a(G326), .O(gate81inter8));
  nand2 gate2124(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2125(.a(s_225), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2126(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2127(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2128(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate743(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate744(.a(gate83inter0), .b(s_28), .O(gate83inter1));
  and2  gate745(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate746(.a(s_28), .O(gate83inter3));
  inv1  gate747(.a(s_29), .O(gate83inter4));
  nand2 gate748(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate749(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate750(.a(G11), .O(gate83inter7));
  inv1  gate751(.a(G329), .O(gate83inter8));
  nand2 gate752(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate753(.a(s_29), .b(gate83inter3), .O(gate83inter10));
  nor2  gate754(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate755(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate756(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate869(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate870(.a(gate105inter0), .b(s_46), .O(gate105inter1));
  and2  gate871(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate872(.a(s_46), .O(gate105inter3));
  inv1  gate873(.a(s_47), .O(gate105inter4));
  nand2 gate874(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate875(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate876(.a(G362), .O(gate105inter7));
  inv1  gate877(.a(G363), .O(gate105inter8));
  nand2 gate878(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate879(.a(s_47), .b(gate105inter3), .O(gate105inter10));
  nor2  gate880(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate881(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate882(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1681(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1682(.a(gate106inter0), .b(s_162), .O(gate106inter1));
  and2  gate1683(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1684(.a(s_162), .O(gate106inter3));
  inv1  gate1685(.a(s_163), .O(gate106inter4));
  nand2 gate1686(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1687(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1688(.a(G364), .O(gate106inter7));
  inv1  gate1689(.a(G365), .O(gate106inter8));
  nand2 gate1690(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1691(.a(s_163), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1692(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1693(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1694(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate967(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate968(.a(gate112inter0), .b(s_60), .O(gate112inter1));
  and2  gate969(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate970(.a(s_60), .O(gate112inter3));
  inv1  gate971(.a(s_61), .O(gate112inter4));
  nand2 gate972(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate973(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate974(.a(G376), .O(gate112inter7));
  inv1  gate975(.a(G377), .O(gate112inter8));
  nand2 gate976(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate977(.a(s_61), .b(gate112inter3), .O(gate112inter10));
  nor2  gate978(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate979(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate980(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1443(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1444(.a(gate125inter0), .b(s_128), .O(gate125inter1));
  and2  gate1445(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1446(.a(s_128), .O(gate125inter3));
  inv1  gate1447(.a(s_129), .O(gate125inter4));
  nand2 gate1448(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1449(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1450(.a(G402), .O(gate125inter7));
  inv1  gate1451(.a(G403), .O(gate125inter8));
  nand2 gate1452(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1453(.a(s_129), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1454(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1455(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1456(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1695(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1696(.a(gate126inter0), .b(s_164), .O(gate126inter1));
  and2  gate1697(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1698(.a(s_164), .O(gate126inter3));
  inv1  gate1699(.a(s_165), .O(gate126inter4));
  nand2 gate1700(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1701(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1702(.a(G404), .O(gate126inter7));
  inv1  gate1703(.a(G405), .O(gate126inter8));
  nand2 gate1704(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1705(.a(s_165), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1706(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1707(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1708(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1485(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1486(.a(gate132inter0), .b(s_134), .O(gate132inter1));
  and2  gate1487(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1488(.a(s_134), .O(gate132inter3));
  inv1  gate1489(.a(s_135), .O(gate132inter4));
  nand2 gate1490(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1491(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1492(.a(G416), .O(gate132inter7));
  inv1  gate1493(.a(G417), .O(gate132inter8));
  nand2 gate1494(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1495(.a(s_135), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1496(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1497(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1498(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1261(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1262(.a(gate135inter0), .b(s_102), .O(gate135inter1));
  and2  gate1263(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1264(.a(s_102), .O(gate135inter3));
  inv1  gate1265(.a(s_103), .O(gate135inter4));
  nand2 gate1266(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1267(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1268(.a(G422), .O(gate135inter7));
  inv1  gate1269(.a(G423), .O(gate135inter8));
  nand2 gate1270(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1271(.a(s_103), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1272(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1273(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1274(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate995(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate996(.a(gate136inter0), .b(s_64), .O(gate136inter1));
  and2  gate997(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate998(.a(s_64), .O(gate136inter3));
  inv1  gate999(.a(s_65), .O(gate136inter4));
  nand2 gate1000(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1001(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1002(.a(G424), .O(gate136inter7));
  inv1  gate1003(.a(G425), .O(gate136inter8));
  nand2 gate1004(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1005(.a(s_65), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1006(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1007(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1008(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1709(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1710(.a(gate144inter0), .b(s_166), .O(gate144inter1));
  and2  gate1711(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1712(.a(s_166), .O(gate144inter3));
  inv1  gate1713(.a(s_167), .O(gate144inter4));
  nand2 gate1714(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1715(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1716(.a(G468), .O(gate144inter7));
  inv1  gate1717(.a(G471), .O(gate144inter8));
  nand2 gate1718(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1719(.a(s_167), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1720(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1721(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1722(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate911(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate912(.a(gate145inter0), .b(s_52), .O(gate145inter1));
  and2  gate913(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate914(.a(s_52), .O(gate145inter3));
  inv1  gate915(.a(s_53), .O(gate145inter4));
  nand2 gate916(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate917(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate918(.a(G474), .O(gate145inter7));
  inv1  gate919(.a(G477), .O(gate145inter8));
  nand2 gate920(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate921(.a(s_53), .b(gate145inter3), .O(gate145inter10));
  nor2  gate922(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate923(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate924(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1149(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1150(.a(gate147inter0), .b(s_86), .O(gate147inter1));
  and2  gate1151(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1152(.a(s_86), .O(gate147inter3));
  inv1  gate1153(.a(s_87), .O(gate147inter4));
  nand2 gate1154(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1155(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1156(.a(G486), .O(gate147inter7));
  inv1  gate1157(.a(G489), .O(gate147inter8));
  nand2 gate1158(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1159(.a(s_87), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1160(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1161(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1162(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1723(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1724(.a(gate148inter0), .b(s_168), .O(gate148inter1));
  and2  gate1725(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1726(.a(s_168), .O(gate148inter3));
  inv1  gate1727(.a(s_169), .O(gate148inter4));
  nand2 gate1728(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1729(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1730(.a(G492), .O(gate148inter7));
  inv1  gate1731(.a(G495), .O(gate148inter8));
  nand2 gate1732(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1733(.a(s_169), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1734(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1735(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1736(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2199(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2200(.a(gate150inter0), .b(s_236), .O(gate150inter1));
  and2  gate2201(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2202(.a(s_236), .O(gate150inter3));
  inv1  gate2203(.a(s_237), .O(gate150inter4));
  nand2 gate2204(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2205(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2206(.a(G504), .O(gate150inter7));
  inv1  gate2207(.a(G507), .O(gate150inter8));
  nand2 gate2208(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2209(.a(s_237), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2210(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2211(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2212(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1303(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1304(.a(gate153inter0), .b(s_108), .O(gate153inter1));
  and2  gate1305(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1306(.a(s_108), .O(gate153inter3));
  inv1  gate1307(.a(s_109), .O(gate153inter4));
  nand2 gate1308(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1309(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1310(.a(G426), .O(gate153inter7));
  inv1  gate1311(.a(G522), .O(gate153inter8));
  nand2 gate1312(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1313(.a(s_109), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1314(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1315(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1316(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2143(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2144(.a(gate154inter0), .b(s_228), .O(gate154inter1));
  and2  gate2145(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2146(.a(s_228), .O(gate154inter3));
  inv1  gate2147(.a(s_229), .O(gate154inter4));
  nand2 gate2148(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2149(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2150(.a(G429), .O(gate154inter7));
  inv1  gate2151(.a(G522), .O(gate154inter8));
  nand2 gate2152(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2153(.a(s_229), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2154(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2155(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2156(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1863(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1864(.a(gate155inter0), .b(s_188), .O(gate155inter1));
  and2  gate1865(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1866(.a(s_188), .O(gate155inter3));
  inv1  gate1867(.a(s_189), .O(gate155inter4));
  nand2 gate1868(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1869(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1870(.a(G432), .O(gate155inter7));
  inv1  gate1871(.a(G525), .O(gate155inter8));
  nand2 gate1872(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1873(.a(s_189), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1874(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1875(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1876(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2101(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2102(.a(gate161inter0), .b(s_222), .O(gate161inter1));
  and2  gate2103(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2104(.a(s_222), .O(gate161inter3));
  inv1  gate2105(.a(s_223), .O(gate161inter4));
  nand2 gate2106(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2107(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2108(.a(G450), .O(gate161inter7));
  inv1  gate2109(.a(G534), .O(gate161inter8));
  nand2 gate2110(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2111(.a(s_223), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2112(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2113(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2114(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1191(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1192(.a(gate162inter0), .b(s_92), .O(gate162inter1));
  and2  gate1193(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1194(.a(s_92), .O(gate162inter3));
  inv1  gate1195(.a(s_93), .O(gate162inter4));
  nand2 gate1196(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1197(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1198(.a(G453), .O(gate162inter7));
  inv1  gate1199(.a(G534), .O(gate162inter8));
  nand2 gate1200(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1201(.a(s_93), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1202(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1203(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1204(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate1205(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1206(.a(gate163inter0), .b(s_94), .O(gate163inter1));
  and2  gate1207(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1208(.a(s_94), .O(gate163inter3));
  inv1  gate1209(.a(s_95), .O(gate163inter4));
  nand2 gate1210(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1211(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1212(.a(G456), .O(gate163inter7));
  inv1  gate1213(.a(G537), .O(gate163inter8));
  nand2 gate1214(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1215(.a(s_95), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1216(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1217(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1218(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1079(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1080(.a(gate165inter0), .b(s_76), .O(gate165inter1));
  and2  gate1081(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1082(.a(s_76), .O(gate165inter3));
  inv1  gate1083(.a(s_77), .O(gate165inter4));
  nand2 gate1084(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1085(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1086(.a(G462), .O(gate165inter7));
  inv1  gate1087(.a(G540), .O(gate165inter8));
  nand2 gate1088(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1089(.a(s_77), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1090(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1091(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1092(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate981(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate982(.a(gate166inter0), .b(s_62), .O(gate166inter1));
  and2  gate983(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate984(.a(s_62), .O(gate166inter3));
  inv1  gate985(.a(s_63), .O(gate166inter4));
  nand2 gate986(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate987(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate988(.a(G465), .O(gate166inter7));
  inv1  gate989(.a(G540), .O(gate166inter8));
  nand2 gate990(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate991(.a(s_63), .b(gate166inter3), .O(gate166inter10));
  nor2  gate992(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate993(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate994(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1905(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1906(.a(gate167inter0), .b(s_194), .O(gate167inter1));
  and2  gate1907(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1908(.a(s_194), .O(gate167inter3));
  inv1  gate1909(.a(s_195), .O(gate167inter4));
  nand2 gate1910(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1911(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1912(.a(G468), .O(gate167inter7));
  inv1  gate1913(.a(G543), .O(gate167inter8));
  nand2 gate1914(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1915(.a(s_195), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1916(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1917(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1918(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate715(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate716(.a(gate168inter0), .b(s_24), .O(gate168inter1));
  and2  gate717(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate718(.a(s_24), .O(gate168inter3));
  inv1  gate719(.a(s_25), .O(gate168inter4));
  nand2 gate720(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate721(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate722(.a(G471), .O(gate168inter7));
  inv1  gate723(.a(G543), .O(gate168inter8));
  nand2 gate724(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate725(.a(s_25), .b(gate168inter3), .O(gate168inter10));
  nor2  gate726(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate727(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate728(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1373(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1374(.a(gate171inter0), .b(s_118), .O(gate171inter1));
  and2  gate1375(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1376(.a(s_118), .O(gate171inter3));
  inv1  gate1377(.a(s_119), .O(gate171inter4));
  nand2 gate1378(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1379(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1380(.a(G480), .O(gate171inter7));
  inv1  gate1381(.a(G549), .O(gate171inter8));
  nand2 gate1382(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1383(.a(s_119), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1384(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1385(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1386(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1023(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1024(.a(gate177inter0), .b(s_68), .O(gate177inter1));
  and2  gate1025(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1026(.a(s_68), .O(gate177inter3));
  inv1  gate1027(.a(s_69), .O(gate177inter4));
  nand2 gate1028(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1029(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1030(.a(G498), .O(gate177inter7));
  inv1  gate1031(.a(G558), .O(gate177inter8));
  nand2 gate1032(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1033(.a(s_69), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1034(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1035(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1036(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1555(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1556(.a(gate178inter0), .b(s_144), .O(gate178inter1));
  and2  gate1557(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1558(.a(s_144), .O(gate178inter3));
  inv1  gate1559(.a(s_145), .O(gate178inter4));
  nand2 gate1560(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1561(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1562(.a(G501), .O(gate178inter7));
  inv1  gate1563(.a(G558), .O(gate178inter8));
  nand2 gate1564(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1565(.a(s_145), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1566(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1567(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1568(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate631(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate632(.a(gate180inter0), .b(s_12), .O(gate180inter1));
  and2  gate633(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate634(.a(s_12), .O(gate180inter3));
  inv1  gate635(.a(s_13), .O(gate180inter4));
  nand2 gate636(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate637(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate638(.a(G507), .O(gate180inter7));
  inv1  gate639(.a(G561), .O(gate180inter8));
  nand2 gate640(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate641(.a(s_13), .b(gate180inter3), .O(gate180inter10));
  nor2  gate642(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate643(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate644(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate617(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate618(.a(gate183inter0), .b(s_10), .O(gate183inter1));
  and2  gate619(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate620(.a(s_10), .O(gate183inter3));
  inv1  gate621(.a(s_11), .O(gate183inter4));
  nand2 gate622(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate623(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate624(.a(G516), .O(gate183inter7));
  inv1  gate625(.a(G567), .O(gate183inter8));
  nand2 gate626(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate627(.a(s_11), .b(gate183inter3), .O(gate183inter10));
  nor2  gate628(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate629(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate630(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate589(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate590(.a(gate185inter0), .b(s_6), .O(gate185inter1));
  and2  gate591(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate592(.a(s_6), .O(gate185inter3));
  inv1  gate593(.a(s_7), .O(gate185inter4));
  nand2 gate594(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate595(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate596(.a(G570), .O(gate185inter7));
  inv1  gate597(.a(G571), .O(gate185inter8));
  nand2 gate598(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate599(.a(s_7), .b(gate185inter3), .O(gate185inter10));
  nor2  gate600(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate601(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate602(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate561(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate562(.a(gate188inter0), .b(s_2), .O(gate188inter1));
  and2  gate563(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate564(.a(s_2), .O(gate188inter3));
  inv1  gate565(.a(s_3), .O(gate188inter4));
  nand2 gate566(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate567(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate568(.a(G576), .O(gate188inter7));
  inv1  gate569(.a(G577), .O(gate188inter8));
  nand2 gate570(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate571(.a(s_3), .b(gate188inter3), .O(gate188inter10));
  nor2  gate572(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate573(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate574(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1751(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1752(.a(gate194inter0), .b(s_172), .O(gate194inter1));
  and2  gate1753(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1754(.a(s_172), .O(gate194inter3));
  inv1  gate1755(.a(s_173), .O(gate194inter4));
  nand2 gate1756(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1757(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1758(.a(G588), .O(gate194inter7));
  inv1  gate1759(.a(G589), .O(gate194inter8));
  nand2 gate1760(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1761(.a(s_173), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1762(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1763(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1764(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate799(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate800(.a(gate199inter0), .b(s_36), .O(gate199inter1));
  and2  gate801(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate802(.a(s_36), .O(gate199inter3));
  inv1  gate803(.a(s_37), .O(gate199inter4));
  nand2 gate804(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate805(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate806(.a(G598), .O(gate199inter7));
  inv1  gate807(.a(G599), .O(gate199inter8));
  nand2 gate808(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate809(.a(s_37), .b(gate199inter3), .O(gate199inter10));
  nor2  gate810(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate811(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate812(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1835(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1836(.a(gate200inter0), .b(s_184), .O(gate200inter1));
  and2  gate1837(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1838(.a(s_184), .O(gate200inter3));
  inv1  gate1839(.a(s_185), .O(gate200inter4));
  nand2 gate1840(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1841(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1842(.a(G600), .O(gate200inter7));
  inv1  gate1843(.a(G601), .O(gate200inter8));
  nand2 gate1844(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1845(.a(s_185), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1846(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1847(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1848(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1457(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1458(.a(gate201inter0), .b(s_130), .O(gate201inter1));
  and2  gate1459(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1460(.a(s_130), .O(gate201inter3));
  inv1  gate1461(.a(s_131), .O(gate201inter4));
  nand2 gate1462(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1463(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1464(.a(G602), .O(gate201inter7));
  inv1  gate1465(.a(G607), .O(gate201inter8));
  nand2 gate1466(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1467(.a(s_131), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1468(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1469(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1470(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1289(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1290(.a(gate202inter0), .b(s_106), .O(gate202inter1));
  and2  gate1291(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1292(.a(s_106), .O(gate202inter3));
  inv1  gate1293(.a(s_107), .O(gate202inter4));
  nand2 gate1294(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1295(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1296(.a(G612), .O(gate202inter7));
  inv1  gate1297(.a(G617), .O(gate202inter8));
  nand2 gate1298(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1299(.a(s_107), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1300(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1301(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1302(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1947(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1948(.a(gate203inter0), .b(s_200), .O(gate203inter1));
  and2  gate1949(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1950(.a(s_200), .O(gate203inter3));
  inv1  gate1951(.a(s_201), .O(gate203inter4));
  nand2 gate1952(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1953(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1954(.a(G602), .O(gate203inter7));
  inv1  gate1955(.a(G612), .O(gate203inter8));
  nand2 gate1956(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1957(.a(s_201), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1958(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1959(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1960(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1989(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1990(.a(gate208inter0), .b(s_206), .O(gate208inter1));
  and2  gate1991(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1992(.a(s_206), .O(gate208inter3));
  inv1  gate1993(.a(s_207), .O(gate208inter4));
  nand2 gate1994(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1995(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1996(.a(G627), .O(gate208inter7));
  inv1  gate1997(.a(G637), .O(gate208inter8));
  nand2 gate1998(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1999(.a(s_207), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2000(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2001(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2002(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1779(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1780(.a(gate210inter0), .b(s_176), .O(gate210inter1));
  and2  gate1781(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1782(.a(s_176), .O(gate210inter3));
  inv1  gate1783(.a(s_177), .O(gate210inter4));
  nand2 gate1784(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1785(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1786(.a(G607), .O(gate210inter7));
  inv1  gate1787(.a(G666), .O(gate210inter8));
  nand2 gate1788(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1789(.a(s_177), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1790(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1791(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1792(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1653(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1654(.a(gate211inter0), .b(s_158), .O(gate211inter1));
  and2  gate1655(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1656(.a(s_158), .O(gate211inter3));
  inv1  gate1657(.a(s_159), .O(gate211inter4));
  nand2 gate1658(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1659(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1660(.a(G612), .O(gate211inter7));
  inv1  gate1661(.a(G669), .O(gate211inter8));
  nand2 gate1662(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1663(.a(s_159), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1664(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1665(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1666(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2045(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2046(.a(gate212inter0), .b(s_214), .O(gate212inter1));
  and2  gate2047(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2048(.a(s_214), .O(gate212inter3));
  inv1  gate2049(.a(s_215), .O(gate212inter4));
  nand2 gate2050(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2051(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2052(.a(G617), .O(gate212inter7));
  inv1  gate2053(.a(G669), .O(gate212inter8));
  nand2 gate2054(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2055(.a(s_215), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2056(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2057(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2058(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1177(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1178(.a(gate218inter0), .b(s_90), .O(gate218inter1));
  and2  gate1179(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1180(.a(s_90), .O(gate218inter3));
  inv1  gate1181(.a(s_91), .O(gate218inter4));
  nand2 gate1182(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1183(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1184(.a(G627), .O(gate218inter7));
  inv1  gate1185(.a(G678), .O(gate218inter8));
  nand2 gate1186(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1187(.a(s_91), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1188(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1189(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1190(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate547(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate548(.a(gate222inter0), .b(s_0), .O(gate222inter1));
  and2  gate549(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate550(.a(s_0), .O(gate222inter3));
  inv1  gate551(.a(s_1), .O(gate222inter4));
  nand2 gate552(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate553(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate554(.a(G632), .O(gate222inter7));
  inv1  gate555(.a(G684), .O(gate222inter8));
  nand2 gate556(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate557(.a(s_1), .b(gate222inter3), .O(gate222inter10));
  nor2  gate558(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate559(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate560(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1513(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1514(.a(gate239inter0), .b(s_138), .O(gate239inter1));
  and2  gate1515(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1516(.a(s_138), .O(gate239inter3));
  inv1  gate1517(.a(s_139), .O(gate239inter4));
  nand2 gate1518(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1519(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1520(.a(G260), .O(gate239inter7));
  inv1  gate1521(.a(G712), .O(gate239inter8));
  nand2 gate1522(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1523(.a(s_139), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1524(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1525(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1526(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate925(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate926(.a(gate240inter0), .b(s_54), .O(gate240inter1));
  and2  gate927(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate928(.a(s_54), .O(gate240inter3));
  inv1  gate929(.a(s_55), .O(gate240inter4));
  nand2 gate930(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate931(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate932(.a(G263), .O(gate240inter7));
  inv1  gate933(.a(G715), .O(gate240inter8));
  nand2 gate934(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate935(.a(s_55), .b(gate240inter3), .O(gate240inter10));
  nor2  gate936(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate937(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate938(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1471(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1472(.a(gate241inter0), .b(s_132), .O(gate241inter1));
  and2  gate1473(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1474(.a(s_132), .O(gate241inter3));
  inv1  gate1475(.a(s_133), .O(gate241inter4));
  nand2 gate1476(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1477(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1478(.a(G242), .O(gate241inter7));
  inv1  gate1479(.a(G730), .O(gate241inter8));
  nand2 gate1480(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1481(.a(s_133), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1482(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1483(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1484(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1597(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1598(.a(gate256inter0), .b(s_150), .O(gate256inter1));
  and2  gate1599(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1600(.a(s_150), .O(gate256inter3));
  inv1  gate1601(.a(s_151), .O(gate256inter4));
  nand2 gate1602(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1603(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1604(.a(G715), .O(gate256inter7));
  inv1  gate1605(.a(G751), .O(gate256inter8));
  nand2 gate1606(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1607(.a(s_151), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1608(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1609(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1610(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1569(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1570(.a(gate258inter0), .b(s_146), .O(gate258inter1));
  and2  gate1571(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1572(.a(s_146), .O(gate258inter3));
  inv1  gate1573(.a(s_147), .O(gate258inter4));
  nand2 gate1574(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1575(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1576(.a(G756), .O(gate258inter7));
  inv1  gate1577(.a(G757), .O(gate258inter8));
  nand2 gate1578(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1579(.a(s_147), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1580(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1581(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1582(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1009(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1010(.a(gate259inter0), .b(s_66), .O(gate259inter1));
  and2  gate1011(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1012(.a(s_66), .O(gate259inter3));
  inv1  gate1013(.a(s_67), .O(gate259inter4));
  nand2 gate1014(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1015(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1016(.a(G758), .O(gate259inter7));
  inv1  gate1017(.a(G759), .O(gate259inter8));
  nand2 gate1018(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1019(.a(s_67), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1020(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1021(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1022(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1317(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1318(.a(gate262inter0), .b(s_110), .O(gate262inter1));
  and2  gate1319(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1320(.a(s_110), .O(gate262inter3));
  inv1  gate1321(.a(s_111), .O(gate262inter4));
  nand2 gate1322(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1323(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1324(.a(G764), .O(gate262inter7));
  inv1  gate1325(.a(G765), .O(gate262inter8));
  nand2 gate1326(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1327(.a(s_111), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1328(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1329(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1330(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1135(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1136(.a(gate263inter0), .b(s_84), .O(gate263inter1));
  and2  gate1137(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1138(.a(s_84), .O(gate263inter3));
  inv1  gate1139(.a(s_85), .O(gate263inter4));
  nand2 gate1140(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1141(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1142(.a(G766), .O(gate263inter7));
  inv1  gate1143(.a(G767), .O(gate263inter8));
  nand2 gate1144(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1145(.a(s_85), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1146(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1147(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1148(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2087(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2088(.a(gate270inter0), .b(s_220), .O(gate270inter1));
  and2  gate2089(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2090(.a(s_220), .O(gate270inter3));
  inv1  gate2091(.a(s_221), .O(gate270inter4));
  nand2 gate2092(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2093(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2094(.a(G657), .O(gate270inter7));
  inv1  gate2095(.a(G785), .O(gate270inter8));
  nand2 gate2096(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2097(.a(s_221), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2098(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2099(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2100(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2017(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2018(.a(gate272inter0), .b(s_210), .O(gate272inter1));
  and2  gate2019(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2020(.a(s_210), .O(gate272inter3));
  inv1  gate2021(.a(s_211), .O(gate272inter4));
  nand2 gate2022(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2023(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2024(.a(G663), .O(gate272inter7));
  inv1  gate2025(.a(G791), .O(gate272inter8));
  nand2 gate2026(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2027(.a(s_211), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2028(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2029(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2030(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1667(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1668(.a(gate282inter0), .b(s_160), .O(gate282inter1));
  and2  gate1669(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1670(.a(s_160), .O(gate282inter3));
  inv1  gate1671(.a(s_161), .O(gate282inter4));
  nand2 gate1672(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1673(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1674(.a(G782), .O(gate282inter7));
  inv1  gate1675(.a(G806), .O(gate282inter8));
  nand2 gate1676(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1677(.a(s_161), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1678(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1679(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1680(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1737(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1738(.a(gate284inter0), .b(s_170), .O(gate284inter1));
  and2  gate1739(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1740(.a(s_170), .O(gate284inter3));
  inv1  gate1741(.a(s_171), .O(gate284inter4));
  nand2 gate1742(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1743(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1744(.a(G785), .O(gate284inter7));
  inv1  gate1745(.a(G809), .O(gate284inter8));
  nand2 gate1746(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1747(.a(s_171), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1748(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1749(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1750(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate953(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate954(.a(gate286inter0), .b(s_58), .O(gate286inter1));
  and2  gate955(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate956(.a(s_58), .O(gate286inter3));
  inv1  gate957(.a(s_59), .O(gate286inter4));
  nand2 gate958(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate959(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate960(.a(G788), .O(gate286inter7));
  inv1  gate961(.a(G812), .O(gate286inter8));
  nand2 gate962(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate963(.a(s_59), .b(gate286inter3), .O(gate286inter10));
  nor2  gate964(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate965(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate966(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate897(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate898(.a(gate288inter0), .b(s_50), .O(gate288inter1));
  and2  gate899(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate900(.a(s_50), .O(gate288inter3));
  inv1  gate901(.a(s_51), .O(gate288inter4));
  nand2 gate902(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate903(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate904(.a(G791), .O(gate288inter7));
  inv1  gate905(.a(G815), .O(gate288inter8));
  nand2 gate906(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate907(.a(s_51), .b(gate288inter3), .O(gate288inter10));
  nor2  gate908(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate909(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate910(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1219(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1220(.a(gate291inter0), .b(s_96), .O(gate291inter1));
  and2  gate1221(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1222(.a(s_96), .O(gate291inter3));
  inv1  gate1223(.a(s_97), .O(gate291inter4));
  nand2 gate1224(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1225(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1226(.a(G822), .O(gate291inter7));
  inv1  gate1227(.a(G823), .O(gate291inter8));
  nand2 gate1228(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1229(.a(s_97), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1230(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1231(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1232(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate645(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate646(.a(gate292inter0), .b(s_14), .O(gate292inter1));
  and2  gate647(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate648(.a(s_14), .O(gate292inter3));
  inv1  gate649(.a(s_15), .O(gate292inter4));
  nand2 gate650(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate651(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate652(.a(G824), .O(gate292inter7));
  inv1  gate653(.a(G825), .O(gate292inter8));
  nand2 gate654(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate655(.a(s_15), .b(gate292inter3), .O(gate292inter10));
  nor2  gate656(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate657(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate658(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1247(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1248(.a(gate293inter0), .b(s_100), .O(gate293inter1));
  and2  gate1249(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1250(.a(s_100), .O(gate293inter3));
  inv1  gate1251(.a(s_101), .O(gate293inter4));
  nand2 gate1252(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1253(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1254(.a(G828), .O(gate293inter7));
  inv1  gate1255(.a(G829), .O(gate293inter8));
  nand2 gate1256(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1257(.a(s_101), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1258(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1259(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1260(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate701(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate702(.a(gate392inter0), .b(s_22), .O(gate392inter1));
  and2  gate703(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate704(.a(s_22), .O(gate392inter3));
  inv1  gate705(.a(s_23), .O(gate392inter4));
  nand2 gate706(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate707(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate708(.a(G6), .O(gate392inter7));
  inv1  gate709(.a(G1051), .O(gate392inter8));
  nand2 gate710(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate711(.a(s_23), .b(gate392inter3), .O(gate392inter10));
  nor2  gate712(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate713(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate714(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1849(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1850(.a(gate394inter0), .b(s_186), .O(gate394inter1));
  and2  gate1851(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1852(.a(s_186), .O(gate394inter3));
  inv1  gate1853(.a(s_187), .O(gate394inter4));
  nand2 gate1854(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1855(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1856(.a(G8), .O(gate394inter7));
  inv1  gate1857(.a(G1057), .O(gate394inter8));
  nand2 gate1858(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1859(.a(s_187), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1860(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1861(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1862(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1933(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1934(.a(gate395inter0), .b(s_198), .O(gate395inter1));
  and2  gate1935(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1936(.a(s_198), .O(gate395inter3));
  inv1  gate1937(.a(s_199), .O(gate395inter4));
  nand2 gate1938(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1939(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1940(.a(G9), .O(gate395inter7));
  inv1  gate1941(.a(G1060), .O(gate395inter8));
  nand2 gate1942(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1943(.a(s_199), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1944(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1945(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1946(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1065(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1066(.a(gate399inter0), .b(s_74), .O(gate399inter1));
  and2  gate1067(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1068(.a(s_74), .O(gate399inter3));
  inv1  gate1069(.a(s_75), .O(gate399inter4));
  nand2 gate1070(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1071(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1072(.a(G13), .O(gate399inter7));
  inv1  gate1073(.a(G1072), .O(gate399inter8));
  nand2 gate1074(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1075(.a(s_75), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1076(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1077(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1078(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1625(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1626(.a(gate401inter0), .b(s_154), .O(gate401inter1));
  and2  gate1627(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1628(.a(s_154), .O(gate401inter3));
  inv1  gate1629(.a(s_155), .O(gate401inter4));
  nand2 gate1630(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1631(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1632(.a(G15), .O(gate401inter7));
  inv1  gate1633(.a(G1078), .O(gate401inter8));
  nand2 gate1634(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1635(.a(s_155), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1636(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1637(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1638(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1541(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1542(.a(gate404inter0), .b(s_142), .O(gate404inter1));
  and2  gate1543(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1544(.a(s_142), .O(gate404inter3));
  inv1  gate1545(.a(s_143), .O(gate404inter4));
  nand2 gate1546(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1547(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1548(.a(G18), .O(gate404inter7));
  inv1  gate1549(.a(G1087), .O(gate404inter8));
  nand2 gate1550(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1551(.a(s_143), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1552(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1553(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1554(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2003(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2004(.a(gate408inter0), .b(s_208), .O(gate408inter1));
  and2  gate2005(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2006(.a(s_208), .O(gate408inter3));
  inv1  gate2007(.a(s_209), .O(gate408inter4));
  nand2 gate2008(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2009(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2010(.a(G22), .O(gate408inter7));
  inv1  gate2011(.a(G1099), .O(gate408inter8));
  nand2 gate2012(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2013(.a(s_209), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2014(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2015(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2016(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1359(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1360(.a(gate410inter0), .b(s_116), .O(gate410inter1));
  and2  gate1361(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1362(.a(s_116), .O(gate410inter3));
  inv1  gate1363(.a(s_117), .O(gate410inter4));
  nand2 gate1364(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1365(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1366(.a(G24), .O(gate410inter7));
  inv1  gate1367(.a(G1105), .O(gate410inter8));
  nand2 gate1368(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1369(.a(s_117), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1370(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1371(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1372(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate2213(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2214(.a(gate411inter0), .b(s_238), .O(gate411inter1));
  and2  gate2215(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2216(.a(s_238), .O(gate411inter3));
  inv1  gate2217(.a(s_239), .O(gate411inter4));
  nand2 gate2218(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2219(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2220(.a(G25), .O(gate411inter7));
  inv1  gate2221(.a(G1108), .O(gate411inter8));
  nand2 gate2222(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2223(.a(s_239), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2224(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2225(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2226(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate771(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate772(.a(gate414inter0), .b(s_32), .O(gate414inter1));
  and2  gate773(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate774(.a(s_32), .O(gate414inter3));
  inv1  gate775(.a(s_33), .O(gate414inter4));
  nand2 gate776(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate777(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate778(.a(G28), .O(gate414inter7));
  inv1  gate779(.a(G1117), .O(gate414inter8));
  nand2 gate780(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate781(.a(s_33), .b(gate414inter3), .O(gate414inter10));
  nor2  gate782(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate783(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate784(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1499(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1500(.a(gate417inter0), .b(s_136), .O(gate417inter1));
  and2  gate1501(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1502(.a(s_136), .O(gate417inter3));
  inv1  gate1503(.a(s_137), .O(gate417inter4));
  nand2 gate1504(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1505(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1506(.a(G31), .O(gate417inter7));
  inv1  gate1507(.a(G1126), .O(gate417inter8));
  nand2 gate1508(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1509(.a(s_137), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1510(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1511(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1512(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2073(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2074(.a(gate420inter0), .b(s_218), .O(gate420inter1));
  and2  gate2075(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2076(.a(s_218), .O(gate420inter3));
  inv1  gate2077(.a(s_219), .O(gate420inter4));
  nand2 gate2078(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2079(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2080(.a(G1036), .O(gate420inter7));
  inv1  gate2081(.a(G1132), .O(gate420inter8));
  nand2 gate2082(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2083(.a(s_219), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2084(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2085(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2086(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate855(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate856(.a(gate424inter0), .b(s_44), .O(gate424inter1));
  and2  gate857(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate858(.a(s_44), .O(gate424inter3));
  inv1  gate859(.a(s_45), .O(gate424inter4));
  nand2 gate860(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate861(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate862(.a(G1042), .O(gate424inter7));
  inv1  gate863(.a(G1138), .O(gate424inter8));
  nand2 gate864(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate865(.a(s_45), .b(gate424inter3), .O(gate424inter10));
  nor2  gate866(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate867(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate868(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1611(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1612(.a(gate428inter0), .b(s_152), .O(gate428inter1));
  and2  gate1613(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1614(.a(s_152), .O(gate428inter3));
  inv1  gate1615(.a(s_153), .O(gate428inter4));
  nand2 gate1616(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1617(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1618(.a(G1048), .O(gate428inter7));
  inv1  gate1619(.a(G1144), .O(gate428inter8));
  nand2 gate1620(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1621(.a(s_153), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1622(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1623(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1624(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate757(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate758(.a(gate430inter0), .b(s_30), .O(gate430inter1));
  and2  gate759(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate760(.a(s_30), .O(gate430inter3));
  inv1  gate761(.a(s_31), .O(gate430inter4));
  nand2 gate762(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate763(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate764(.a(G1051), .O(gate430inter7));
  inv1  gate765(.a(G1147), .O(gate430inter8));
  nand2 gate766(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate767(.a(s_31), .b(gate430inter3), .O(gate430inter10));
  nor2  gate768(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate769(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate770(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate827(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate828(.a(gate435inter0), .b(s_40), .O(gate435inter1));
  and2  gate829(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate830(.a(s_40), .O(gate435inter3));
  inv1  gate831(.a(s_41), .O(gate435inter4));
  nand2 gate832(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate833(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate834(.a(G9), .O(gate435inter7));
  inv1  gate835(.a(G1156), .O(gate435inter8));
  nand2 gate836(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate837(.a(s_41), .b(gate435inter3), .O(gate435inter10));
  nor2  gate838(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate839(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate840(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate813(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate814(.a(gate436inter0), .b(s_38), .O(gate436inter1));
  and2  gate815(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate816(.a(s_38), .O(gate436inter3));
  inv1  gate817(.a(s_39), .O(gate436inter4));
  nand2 gate818(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate819(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate820(.a(G1060), .O(gate436inter7));
  inv1  gate821(.a(G1156), .O(gate436inter8));
  nand2 gate822(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate823(.a(s_39), .b(gate436inter3), .O(gate436inter10));
  nor2  gate824(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate825(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate826(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1331(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1332(.a(gate437inter0), .b(s_112), .O(gate437inter1));
  and2  gate1333(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1334(.a(s_112), .O(gate437inter3));
  inv1  gate1335(.a(s_113), .O(gate437inter4));
  nand2 gate1336(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1337(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1338(.a(G10), .O(gate437inter7));
  inv1  gate1339(.a(G1159), .O(gate437inter8));
  nand2 gate1340(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1341(.a(s_113), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1342(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1343(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1344(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1163(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1164(.a(gate440inter0), .b(s_88), .O(gate440inter1));
  and2  gate1165(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1166(.a(s_88), .O(gate440inter3));
  inv1  gate1167(.a(s_89), .O(gate440inter4));
  nand2 gate1168(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1169(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1170(.a(G1066), .O(gate440inter7));
  inv1  gate1171(.a(G1162), .O(gate440inter8));
  nand2 gate1172(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1173(.a(s_89), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1174(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1175(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1176(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1583(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1584(.a(gate445inter0), .b(s_148), .O(gate445inter1));
  and2  gate1585(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1586(.a(s_148), .O(gate445inter3));
  inv1  gate1587(.a(s_149), .O(gate445inter4));
  nand2 gate1588(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1589(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1590(.a(G14), .O(gate445inter7));
  inv1  gate1591(.a(G1171), .O(gate445inter8));
  nand2 gate1592(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1593(.a(s_149), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1594(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1595(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1596(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1037(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1038(.a(gate447inter0), .b(s_70), .O(gate447inter1));
  and2  gate1039(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1040(.a(s_70), .O(gate447inter3));
  inv1  gate1041(.a(s_71), .O(gate447inter4));
  nand2 gate1042(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1043(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1044(.a(G15), .O(gate447inter7));
  inv1  gate1045(.a(G1174), .O(gate447inter8));
  nand2 gate1046(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1047(.a(s_71), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1048(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1049(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1050(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2129(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2130(.a(gate454inter0), .b(s_226), .O(gate454inter1));
  and2  gate2131(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2132(.a(s_226), .O(gate454inter3));
  inv1  gate2133(.a(s_227), .O(gate454inter4));
  nand2 gate2134(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2135(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2136(.a(G1087), .O(gate454inter7));
  inv1  gate2137(.a(G1183), .O(gate454inter8));
  nand2 gate2138(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2139(.a(s_227), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2140(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2141(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2142(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate2157(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2158(.a(gate455inter0), .b(s_230), .O(gate455inter1));
  and2  gate2159(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2160(.a(s_230), .O(gate455inter3));
  inv1  gate2161(.a(s_231), .O(gate455inter4));
  nand2 gate2162(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2163(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2164(.a(G19), .O(gate455inter7));
  inv1  gate2165(.a(G1186), .O(gate455inter8));
  nand2 gate2166(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2167(.a(s_231), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2168(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2169(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2170(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate2059(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2060(.a(gate456inter0), .b(s_216), .O(gate456inter1));
  and2  gate2061(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2062(.a(s_216), .O(gate456inter3));
  inv1  gate2063(.a(s_217), .O(gate456inter4));
  nand2 gate2064(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2065(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2066(.a(G1090), .O(gate456inter7));
  inv1  gate2067(.a(G1186), .O(gate456inter8));
  nand2 gate2068(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2069(.a(s_217), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2070(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2071(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2072(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1275(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1276(.a(gate458inter0), .b(s_104), .O(gate458inter1));
  and2  gate1277(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1278(.a(s_104), .O(gate458inter3));
  inv1  gate1279(.a(s_105), .O(gate458inter4));
  nand2 gate1280(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1281(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1282(.a(G1093), .O(gate458inter7));
  inv1  gate1283(.a(G1189), .O(gate458inter8));
  nand2 gate1284(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1285(.a(s_105), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1286(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1287(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1288(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate785(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate786(.a(gate460inter0), .b(s_34), .O(gate460inter1));
  and2  gate787(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate788(.a(s_34), .O(gate460inter3));
  inv1  gate789(.a(s_35), .O(gate460inter4));
  nand2 gate790(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate791(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate792(.a(G1096), .O(gate460inter7));
  inv1  gate793(.a(G1192), .O(gate460inter8));
  nand2 gate794(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate795(.a(s_35), .b(gate460inter3), .O(gate460inter10));
  nor2  gate796(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate797(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate798(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate1919(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1920(.a(gate461inter0), .b(s_196), .O(gate461inter1));
  and2  gate1921(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1922(.a(s_196), .O(gate461inter3));
  inv1  gate1923(.a(s_197), .O(gate461inter4));
  nand2 gate1924(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1925(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1926(.a(G22), .O(gate461inter7));
  inv1  gate1927(.a(G1195), .O(gate461inter8));
  nand2 gate1928(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1929(.a(s_197), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1930(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1931(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1932(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate1121(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1122(.a(gate462inter0), .b(s_82), .O(gate462inter1));
  and2  gate1123(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1124(.a(s_82), .O(gate462inter3));
  inv1  gate1125(.a(s_83), .O(gate462inter4));
  nand2 gate1126(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1127(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1128(.a(G1099), .O(gate462inter7));
  inv1  gate1129(.a(G1195), .O(gate462inter8));
  nand2 gate1130(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1131(.a(s_83), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1132(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1133(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1134(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1793(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1794(.a(gate463inter0), .b(s_178), .O(gate463inter1));
  and2  gate1795(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1796(.a(s_178), .O(gate463inter3));
  inv1  gate1797(.a(s_179), .O(gate463inter4));
  nand2 gate1798(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1799(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1800(.a(G23), .O(gate463inter7));
  inv1  gate1801(.a(G1198), .O(gate463inter8));
  nand2 gate1802(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1803(.a(s_179), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1804(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1805(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1806(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2031(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2032(.a(gate465inter0), .b(s_212), .O(gate465inter1));
  and2  gate2033(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2034(.a(s_212), .O(gate465inter3));
  inv1  gate2035(.a(s_213), .O(gate465inter4));
  nand2 gate2036(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2037(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2038(.a(G24), .O(gate465inter7));
  inv1  gate2039(.a(G1201), .O(gate465inter8));
  nand2 gate2040(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2041(.a(s_213), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2042(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2043(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2044(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate939(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate940(.a(gate467inter0), .b(s_56), .O(gate467inter1));
  and2  gate941(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate942(.a(s_56), .O(gate467inter3));
  inv1  gate943(.a(s_57), .O(gate467inter4));
  nand2 gate944(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate945(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate946(.a(G25), .O(gate467inter7));
  inv1  gate947(.a(G1204), .O(gate467inter8));
  nand2 gate948(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate949(.a(s_57), .b(gate467inter3), .O(gate467inter10));
  nor2  gate950(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate951(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate952(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1429(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1430(.a(gate468inter0), .b(s_126), .O(gate468inter1));
  and2  gate1431(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1432(.a(s_126), .O(gate468inter3));
  inv1  gate1433(.a(s_127), .O(gate468inter4));
  nand2 gate1434(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1435(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1436(.a(G1108), .O(gate468inter7));
  inv1  gate1437(.a(G1204), .O(gate468inter8));
  nand2 gate1438(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1439(.a(s_127), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1440(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1441(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1442(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2227(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2228(.a(gate471inter0), .b(s_240), .O(gate471inter1));
  and2  gate2229(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2230(.a(s_240), .O(gate471inter3));
  inv1  gate2231(.a(s_241), .O(gate471inter4));
  nand2 gate2232(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2233(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2234(.a(G27), .O(gate471inter7));
  inv1  gate2235(.a(G1210), .O(gate471inter8));
  nand2 gate2236(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2237(.a(s_241), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2238(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2239(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2240(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate659(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate660(.a(gate475inter0), .b(s_16), .O(gate475inter1));
  and2  gate661(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate662(.a(s_16), .O(gate475inter3));
  inv1  gate663(.a(s_17), .O(gate475inter4));
  nand2 gate664(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate665(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate666(.a(G29), .O(gate475inter7));
  inv1  gate667(.a(G1216), .O(gate475inter8));
  nand2 gate668(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate669(.a(s_17), .b(gate475inter3), .O(gate475inter10));
  nor2  gate670(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate671(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate672(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1807(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1808(.a(gate479inter0), .b(s_180), .O(gate479inter1));
  and2  gate1809(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1810(.a(s_180), .O(gate479inter3));
  inv1  gate1811(.a(s_181), .O(gate479inter4));
  nand2 gate1812(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1813(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1814(.a(G31), .O(gate479inter7));
  inv1  gate1815(.a(G1222), .O(gate479inter8));
  nand2 gate1816(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1817(.a(s_181), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1818(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1819(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1820(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1387(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1388(.a(gate480inter0), .b(s_120), .O(gate480inter1));
  and2  gate1389(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1390(.a(s_120), .O(gate480inter3));
  inv1  gate1391(.a(s_121), .O(gate480inter4));
  nand2 gate1392(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1393(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1394(.a(G1126), .O(gate480inter7));
  inv1  gate1395(.a(G1222), .O(gate480inter8));
  nand2 gate1396(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1397(.a(s_121), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1398(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1399(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1400(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1415(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1416(.a(gate482inter0), .b(s_124), .O(gate482inter1));
  and2  gate1417(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1418(.a(s_124), .O(gate482inter3));
  inv1  gate1419(.a(s_125), .O(gate482inter4));
  nand2 gate1420(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1421(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1422(.a(G1129), .O(gate482inter7));
  inv1  gate1423(.a(G1225), .O(gate482inter8));
  nand2 gate1424(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1425(.a(s_125), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1426(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1427(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1428(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1345(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1346(.a(gate485inter0), .b(s_114), .O(gate485inter1));
  and2  gate1347(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1348(.a(s_114), .O(gate485inter3));
  inv1  gate1349(.a(s_115), .O(gate485inter4));
  nand2 gate1350(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1351(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1352(.a(G1232), .O(gate485inter7));
  inv1  gate1353(.a(G1233), .O(gate485inter8));
  nand2 gate1354(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1355(.a(s_115), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1356(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1357(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1358(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1233(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1234(.a(gate489inter0), .b(s_98), .O(gate489inter1));
  and2  gate1235(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1236(.a(s_98), .O(gate489inter3));
  inv1  gate1237(.a(s_99), .O(gate489inter4));
  nand2 gate1238(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1239(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1240(.a(G1240), .O(gate489inter7));
  inv1  gate1241(.a(G1241), .O(gate489inter8));
  nand2 gate1242(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1243(.a(s_99), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1244(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1245(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1246(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1961(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1962(.a(gate493inter0), .b(s_202), .O(gate493inter1));
  and2  gate1963(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1964(.a(s_202), .O(gate493inter3));
  inv1  gate1965(.a(s_203), .O(gate493inter4));
  nand2 gate1966(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1967(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1968(.a(G1248), .O(gate493inter7));
  inv1  gate1969(.a(G1249), .O(gate493inter8));
  nand2 gate1970(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1971(.a(s_203), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1972(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1973(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1974(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1975(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1976(.a(gate500inter0), .b(s_204), .O(gate500inter1));
  and2  gate1977(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1978(.a(s_204), .O(gate500inter3));
  inv1  gate1979(.a(s_205), .O(gate500inter4));
  nand2 gate1980(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1981(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1982(.a(G1262), .O(gate500inter7));
  inv1  gate1983(.a(G1263), .O(gate500inter8));
  nand2 gate1984(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1985(.a(s_205), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1986(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1987(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1988(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1821(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1822(.a(gate502inter0), .b(s_182), .O(gate502inter1));
  and2  gate1823(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1824(.a(s_182), .O(gate502inter3));
  inv1  gate1825(.a(s_183), .O(gate502inter4));
  nand2 gate1826(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1827(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1828(.a(G1266), .O(gate502inter7));
  inv1  gate1829(.a(G1267), .O(gate502inter8));
  nand2 gate1830(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1831(.a(s_183), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1832(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1833(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1834(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2185(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2186(.a(gate509inter0), .b(s_234), .O(gate509inter1));
  and2  gate2187(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2188(.a(s_234), .O(gate509inter3));
  inv1  gate2189(.a(s_235), .O(gate509inter4));
  nand2 gate2190(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2191(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2192(.a(G1280), .O(gate509inter7));
  inv1  gate2193(.a(G1281), .O(gate509inter8));
  nand2 gate2194(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2195(.a(s_235), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2196(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2197(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2198(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate575(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate576(.a(gate513inter0), .b(s_4), .O(gate513inter1));
  and2  gate577(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate578(.a(s_4), .O(gate513inter3));
  inv1  gate579(.a(s_5), .O(gate513inter4));
  nand2 gate580(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate581(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate582(.a(G1288), .O(gate513inter7));
  inv1  gate583(.a(G1289), .O(gate513inter8));
  nand2 gate584(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate585(.a(s_5), .b(gate513inter3), .O(gate513inter10));
  nor2  gate586(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate587(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate588(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule