module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate679(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate680(.a(gate3inter0), .b(s_68), .O(gate3inter1));
  and2  gate681(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate682(.a(s_68), .O(gate3inter3));
  inv1  gate683(.a(s_69), .O(gate3inter4));
  nand2 gate684(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate685(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate686(.a(N17), .O(gate3inter7));
  inv1  gate687(.a(N21), .O(gate3inter8));
  nand2 gate688(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate689(.a(s_69), .b(gate3inter3), .O(gate3inter10));
  nor2  gate690(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate691(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate692(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );

  xor2  gate343(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate344(.a(gate16inter0), .b(s_20), .O(gate16inter1));
  and2  gate345(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate346(.a(s_20), .O(gate16inter3));
  inv1  gate347(.a(s_21), .O(gate16inter4));
  nand2 gate348(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate349(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate350(.a(N121), .O(gate16inter7));
  inv1  gate351(.a(N125), .O(gate16inter8));
  nand2 gate352(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate353(.a(s_21), .b(gate16inter3), .O(gate16inter10));
  nor2  gate354(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate355(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate356(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate567(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate568(.a(gate25inter0), .b(s_52), .O(gate25inter1));
  and2  gate569(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate570(.a(s_52), .O(gate25inter3));
  inv1  gate571(.a(s_53), .O(gate25inter4));
  nand2 gate572(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate573(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate574(.a(N1), .O(gate25inter7));
  inv1  gate575(.a(N17), .O(gate25inter8));
  nand2 gate576(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate577(.a(s_53), .b(gate25inter3), .O(gate25inter10));
  nor2  gate578(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate579(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate580(.a(gate25inter12), .b(gate25inter1), .O(N274));
xor2 gate26( .a(N33), .b(N49), .O(N275) );

  xor2  gate539(.a(N21), .b(N5), .O(gate27inter0));
  nand2 gate540(.a(gate27inter0), .b(s_48), .O(gate27inter1));
  and2  gate541(.a(N21), .b(N5), .O(gate27inter2));
  inv1  gate542(.a(s_48), .O(gate27inter3));
  inv1  gate543(.a(s_49), .O(gate27inter4));
  nand2 gate544(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate545(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate546(.a(N5), .O(gate27inter7));
  inv1  gate547(.a(N21), .O(gate27inter8));
  nand2 gate548(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate549(.a(s_49), .b(gate27inter3), .O(gate27inter10));
  nor2  gate550(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate551(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate552(.a(gate27inter12), .b(gate27inter1), .O(N276));

  xor2  gate609(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate610(.a(gate28inter0), .b(s_58), .O(gate28inter1));
  and2  gate611(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate612(.a(s_58), .O(gate28inter3));
  inv1  gate613(.a(s_59), .O(gate28inter4));
  nand2 gate614(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate615(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate616(.a(N37), .O(gate28inter7));
  inv1  gate617(.a(N53), .O(gate28inter8));
  nand2 gate618(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate619(.a(s_59), .b(gate28inter3), .O(gate28inter10));
  nor2  gate620(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate621(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate622(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate329(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate330(.a(gate30inter0), .b(s_18), .O(gate30inter1));
  and2  gate331(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate332(.a(s_18), .O(gate30inter3));
  inv1  gate333(.a(s_19), .O(gate30inter4));
  nand2 gate334(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate335(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate336(.a(N41), .O(gate30inter7));
  inv1  gate337(.a(N57), .O(gate30inter8));
  nand2 gate338(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate339(.a(s_19), .b(gate30inter3), .O(gate30inter10));
  nor2  gate340(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate341(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate342(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );

  xor2  gate399(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate400(.a(gate34inter0), .b(s_28), .O(gate34inter1));
  and2  gate401(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate402(.a(s_28), .O(gate34inter3));
  inv1  gate403(.a(s_29), .O(gate34inter4));
  nand2 gate404(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate405(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate406(.a(N97), .O(gate34inter7));
  inv1  gate407(.a(N113), .O(gate34inter8));
  nand2 gate408(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate409(.a(s_29), .b(gate34inter3), .O(gate34inter10));
  nor2  gate410(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate411(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate412(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );

  xor2  gate693(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate694(.a(gate37inter0), .b(s_70), .O(gate37inter1));
  and2  gate695(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate696(.a(s_70), .O(gate37inter3));
  inv1  gate697(.a(s_71), .O(gate37inter4));
  nand2 gate698(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate699(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate700(.a(N73), .O(gate37inter7));
  inv1  gate701(.a(N89), .O(gate37inter8));
  nand2 gate702(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate703(.a(s_71), .b(gate37inter3), .O(gate37inter10));
  nor2  gate704(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate705(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate706(.a(gate37inter12), .b(gate37inter1), .O(N286));
xor2 gate38( .a(N105), .b(N121), .O(N287) );

  xor2  gate455(.a(N93), .b(N77), .O(gate39inter0));
  nand2 gate456(.a(gate39inter0), .b(s_36), .O(gate39inter1));
  and2  gate457(.a(N93), .b(N77), .O(gate39inter2));
  inv1  gate458(.a(s_36), .O(gate39inter3));
  inv1  gate459(.a(s_37), .O(gate39inter4));
  nand2 gate460(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate461(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate462(.a(N77), .O(gate39inter7));
  inv1  gate463(.a(N93), .O(gate39inter8));
  nand2 gate464(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate465(.a(s_37), .b(gate39inter3), .O(gate39inter10));
  nor2  gate466(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate467(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate468(.a(gate39inter12), .b(gate39inter1), .O(N288));
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );

  xor2  gate511(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate512(.a(gate43inter0), .b(s_44), .O(gate43inter1));
  and2  gate513(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate514(.a(s_44), .O(gate43inter3));
  inv1  gate515(.a(s_45), .O(gate43inter4));
  nand2 gate516(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate517(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate518(.a(N254), .O(gate43inter7));
  inv1  gate519(.a(N255), .O(gate43inter8));
  nand2 gate520(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate521(.a(s_45), .b(gate43inter3), .O(gate43inter10));
  nor2  gate522(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate523(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate524(.a(gate43inter12), .b(gate43inter1), .O(N296));
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );

  xor2  gate203(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate204(.a(gate46inter0), .b(s_0), .O(gate46inter1));
  and2  gate205(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate206(.a(s_0), .O(gate46inter3));
  inv1  gate207(.a(s_1), .O(gate46inter4));
  nand2 gate208(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate209(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate210(.a(N260), .O(gate46inter7));
  inv1  gate211(.a(N261), .O(gate46inter8));
  nand2 gate212(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate213(.a(s_1), .b(gate46inter3), .O(gate46inter10));
  nor2  gate214(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate215(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate216(.a(gate46inter12), .b(gate46inter1), .O(N305));
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate231(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate232(.a(gate50inter0), .b(s_4), .O(gate50inter1));
  and2  gate233(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate234(.a(s_4), .O(gate50inter3));
  inv1  gate235(.a(s_5), .O(gate50inter4));
  nand2 gate236(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate237(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate238(.a(N276), .O(gate50inter7));
  inv1  gate239(.a(N277), .O(gate50inter8));
  nand2 gate240(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate241(.a(s_5), .b(gate50inter3), .O(gate50inter10));
  nor2  gate242(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate243(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate244(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate357(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate358(.a(gate55inter0), .b(s_22), .O(gate55inter1));
  and2  gate359(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate360(.a(s_22), .O(gate55inter3));
  inv1  gate361(.a(s_23), .O(gate55inter4));
  nand2 gate362(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate363(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate364(.a(N286), .O(gate55inter7));
  inv1  gate365(.a(N287), .O(gate55inter8));
  nand2 gate366(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate367(.a(s_23), .b(gate55inter3), .O(gate55inter10));
  nor2  gate368(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate369(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate370(.a(gate55inter12), .b(gate55inter1), .O(N320));

  xor2  gate273(.a(N289), .b(N288), .O(gate56inter0));
  nand2 gate274(.a(gate56inter0), .b(s_10), .O(gate56inter1));
  and2  gate275(.a(N289), .b(N288), .O(gate56inter2));
  inv1  gate276(.a(s_10), .O(gate56inter3));
  inv1  gate277(.a(s_11), .O(gate56inter4));
  nand2 gate278(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate279(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate280(.a(N288), .O(gate56inter7));
  inv1  gate281(.a(N289), .O(gate56inter8));
  nand2 gate282(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate283(.a(s_11), .b(gate56inter3), .O(gate56inter10));
  nor2  gate284(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate285(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate286(.a(gate56inter12), .b(gate56inter1), .O(N321));

  xor2  gate315(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate316(.a(gate57inter0), .b(s_16), .O(gate57inter1));
  and2  gate317(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate318(.a(s_16), .O(gate57inter3));
  inv1  gate319(.a(s_17), .O(gate57inter4));
  nand2 gate320(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate321(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate322(.a(N290), .O(gate57inter7));
  inv1  gate323(.a(N293), .O(gate57inter8));
  nand2 gate324(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate325(.a(s_17), .b(gate57inter3), .O(gate57inter10));
  nor2  gate326(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate327(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate328(.a(gate57inter12), .b(gate57inter1), .O(N338));
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );

  xor2  gate553(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate554(.a(gate63inter0), .b(s_50), .O(gate63inter1));
  and2  gate555(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate556(.a(s_50), .O(gate63inter3));
  inv1  gate557(.a(s_51), .O(gate63inter4));
  nand2 gate558(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate559(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate560(.a(N302), .O(gate63inter7));
  inv1  gate561(.a(N308), .O(gate63inter8));
  nand2 gate562(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate563(.a(s_51), .b(gate63inter3), .O(gate63inter10));
  nor2  gate564(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate565(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate566(.a(gate63inter12), .b(gate63inter1), .O(N344));

  xor2  gate385(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate386(.a(gate64inter0), .b(s_26), .O(gate64inter1));
  and2  gate387(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate388(.a(s_26), .O(gate64inter3));
  inv1  gate389(.a(s_27), .O(gate64inter4));
  nand2 gate390(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate391(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate392(.a(N305), .O(gate64inter7));
  inv1  gate393(.a(N311), .O(gate64inter8));
  nand2 gate394(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate395(.a(s_27), .b(gate64inter3), .O(gate64inter10));
  nor2  gate396(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate397(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate398(.a(gate64inter12), .b(gate64inter1), .O(N345));

  xor2  gate287(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate288(.a(gate65inter0), .b(s_12), .O(gate65inter1));
  and2  gate289(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate290(.a(s_12), .O(gate65inter3));
  inv1  gate291(.a(s_13), .O(gate65inter4));
  nand2 gate292(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate293(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate294(.a(N266), .O(gate65inter7));
  inv1  gate295(.a(N342), .O(gate65inter8));
  nand2 gate296(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate297(.a(s_13), .b(gate65inter3), .O(gate65inter10));
  nor2  gate298(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate299(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate300(.a(gate65inter12), .b(gate65inter1), .O(N346));
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate245(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate246(.a(gate70inter0), .b(s_6), .O(gate70inter1));
  and2  gate247(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate248(.a(s_6), .O(gate70inter3));
  inv1  gate249(.a(s_7), .O(gate70inter4));
  nand2 gate250(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate251(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate252(.a(N271), .O(gate70inter7));
  inv1  gate253(.a(N339), .O(gate70inter8));
  nand2 gate254(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate255(.a(s_7), .b(gate70inter3), .O(gate70inter10));
  nor2  gate256(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate257(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate258(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );

  xor2  gate217(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate218(.a(gate73inter0), .b(s_2), .O(gate73inter1));
  and2  gate219(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate220(.a(s_2), .O(gate73inter3));
  inv1  gate221(.a(s_3), .O(gate73inter4));
  nand2 gate222(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate223(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate224(.a(N314), .O(gate73inter7));
  inv1  gate225(.a(N346), .O(gate73inter8));
  nand2 gate226(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate227(.a(s_3), .b(gate73inter3), .O(gate73inter10));
  nor2  gate228(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate229(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate230(.a(gate73inter12), .b(gate73inter1), .O(N354));

  xor2  gate441(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate442(.a(gate74inter0), .b(s_34), .O(gate74inter1));
  and2  gate443(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate444(.a(s_34), .O(gate74inter3));
  inv1  gate445(.a(s_35), .O(gate74inter4));
  nand2 gate446(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate447(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate448(.a(N315), .O(gate74inter7));
  inv1  gate449(.a(N347), .O(gate74inter8));
  nand2 gate450(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate451(.a(s_35), .b(gate74inter3), .O(gate74inter10));
  nor2  gate452(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate453(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate454(.a(gate74inter12), .b(gate74inter1), .O(N367));

  xor2  gate637(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate638(.a(gate75inter0), .b(s_62), .O(gate75inter1));
  and2  gate639(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate640(.a(s_62), .O(gate75inter3));
  inv1  gate641(.a(s_63), .O(gate75inter4));
  nand2 gate642(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate643(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate644(.a(N316), .O(gate75inter7));
  inv1  gate645(.a(N348), .O(gate75inter8));
  nand2 gate646(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate647(.a(s_63), .b(gate75inter3), .O(gate75inter10));
  nor2  gate648(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate649(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate650(.a(gate75inter12), .b(gate75inter1), .O(N380));

  xor2  gate371(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate372(.a(gate76inter0), .b(s_24), .O(gate76inter1));
  and2  gate373(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate374(.a(s_24), .O(gate76inter3));
  inv1  gate375(.a(s_25), .O(gate76inter4));
  nand2 gate376(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate377(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate378(.a(N317), .O(gate76inter7));
  inv1  gate379(.a(N349), .O(gate76inter8));
  nand2 gate380(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate381(.a(s_25), .b(gate76inter3), .O(gate76inter10));
  nor2  gate382(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate383(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate384(.a(gate76inter12), .b(gate76inter1), .O(N393));

  xor2  gate525(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate526(.a(gate77inter0), .b(s_46), .O(gate77inter1));
  and2  gate527(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate528(.a(s_46), .O(gate77inter3));
  inv1  gate529(.a(s_47), .O(gate77inter4));
  nand2 gate530(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate531(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate532(.a(N318), .O(gate77inter7));
  inv1  gate533(.a(N350), .O(gate77inter8));
  nand2 gate534(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate535(.a(s_47), .b(gate77inter3), .O(gate77inter10));
  nor2  gate536(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate537(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate538(.a(gate77inter12), .b(gate77inter1), .O(N406));
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );

  xor2  gate483(.a(N692), .b(N1), .O(gate171inter0));
  nand2 gate484(.a(gate171inter0), .b(s_40), .O(gate171inter1));
  and2  gate485(.a(N692), .b(N1), .O(gate171inter2));
  inv1  gate486(.a(s_40), .O(gate171inter3));
  inv1  gate487(.a(s_41), .O(gate171inter4));
  nand2 gate488(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate489(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate490(.a(N1), .O(gate171inter7));
  inv1  gate491(.a(N692), .O(gate171inter8));
  nand2 gate492(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate493(.a(s_41), .b(gate171inter3), .O(gate171inter10));
  nor2  gate494(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate495(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate496(.a(gate171inter12), .b(gate171inter1), .O(N724));

  xor2  gate301(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate302(.a(gate172inter0), .b(s_14), .O(gate172inter1));
  and2  gate303(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate304(.a(s_14), .O(gate172inter3));
  inv1  gate305(.a(s_15), .O(gate172inter4));
  nand2 gate306(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate307(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate308(.a(N5), .O(gate172inter7));
  inv1  gate309(.a(N693), .O(gate172inter8));
  nand2 gate310(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate311(.a(s_15), .b(gate172inter3), .O(gate172inter10));
  nor2  gate312(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate313(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate314(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );

  xor2  gate651(.a(N695), .b(N13), .O(gate174inter0));
  nand2 gate652(.a(gate174inter0), .b(s_64), .O(gate174inter1));
  and2  gate653(.a(N695), .b(N13), .O(gate174inter2));
  inv1  gate654(.a(s_64), .O(gate174inter3));
  inv1  gate655(.a(s_65), .O(gate174inter4));
  nand2 gate656(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate657(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate658(.a(N13), .O(gate174inter7));
  inv1  gate659(.a(N695), .O(gate174inter8));
  nand2 gate660(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate661(.a(s_65), .b(gate174inter3), .O(gate174inter10));
  nor2  gate662(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate663(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate664(.a(gate174inter12), .b(gate174inter1), .O(N727));
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate665(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate666(.a(gate176inter0), .b(s_66), .O(gate176inter1));
  and2  gate667(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate668(.a(s_66), .O(gate176inter3));
  inv1  gate669(.a(s_67), .O(gate176inter4));
  nand2 gate670(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate671(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate672(.a(N21), .O(gate176inter7));
  inv1  gate673(.a(N697), .O(gate176inter8));
  nand2 gate674(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate675(.a(s_67), .b(gate176inter3), .O(gate176inter10));
  nor2  gate676(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate677(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate678(.a(gate176inter12), .b(gate176inter1), .O(N729));

  xor2  gate581(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate582(.a(gate177inter0), .b(s_54), .O(gate177inter1));
  and2  gate583(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate584(.a(s_54), .O(gate177inter3));
  inv1  gate585(.a(s_55), .O(gate177inter4));
  nand2 gate586(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate587(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate588(.a(N25), .O(gate177inter7));
  inv1  gate589(.a(N698), .O(gate177inter8));
  nand2 gate590(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate591(.a(s_55), .b(gate177inter3), .O(gate177inter10));
  nor2  gate592(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate593(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate594(.a(gate177inter12), .b(gate177inter1), .O(N730));
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );

  xor2  gate469(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate470(.a(gate182inter0), .b(s_38), .O(gate182inter1));
  and2  gate471(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate472(.a(s_38), .O(gate182inter3));
  inv1  gate473(.a(s_39), .O(gate182inter4));
  nand2 gate474(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate475(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate476(.a(N45), .O(gate182inter7));
  inv1  gate477(.a(N703), .O(gate182inter8));
  nand2 gate478(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate479(.a(s_39), .b(gate182inter3), .O(gate182inter10));
  nor2  gate480(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate481(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate482(.a(gate182inter12), .b(gate182inter1), .O(N735));

  xor2  gate259(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate260(.a(gate183inter0), .b(s_8), .O(gate183inter1));
  and2  gate261(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate262(.a(s_8), .O(gate183inter3));
  inv1  gate263(.a(s_9), .O(gate183inter4));
  nand2 gate264(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate265(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate266(.a(N49), .O(gate183inter7));
  inv1  gate267(.a(N704), .O(gate183inter8));
  nand2 gate268(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate269(.a(s_9), .b(gate183inter3), .O(gate183inter10));
  nor2  gate270(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate271(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate272(.a(gate183inter12), .b(gate183inter1), .O(N736));

  xor2  gate413(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate414(.a(gate184inter0), .b(s_30), .O(gate184inter1));
  and2  gate415(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate416(.a(s_30), .O(gate184inter3));
  inv1  gate417(.a(s_31), .O(gate184inter4));
  nand2 gate418(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate419(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate420(.a(N53), .O(gate184inter7));
  inv1  gate421(.a(N705), .O(gate184inter8));
  nand2 gate422(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate423(.a(s_31), .b(gate184inter3), .O(gate184inter10));
  nor2  gate424(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate425(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate426(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );

  xor2  gate497(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate498(.a(gate189inter0), .b(s_42), .O(gate189inter1));
  and2  gate499(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate500(.a(s_42), .O(gate189inter3));
  inv1  gate501(.a(s_43), .O(gate189inter4));
  nand2 gate502(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate503(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate504(.a(N73), .O(gate189inter7));
  inv1  gate505(.a(N710), .O(gate189inter8));
  nand2 gate506(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate507(.a(s_43), .b(gate189inter3), .O(gate189inter10));
  nor2  gate508(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate509(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate510(.a(gate189inter12), .b(gate189inter1), .O(N742));

  xor2  gate427(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate428(.a(gate190inter0), .b(s_32), .O(gate190inter1));
  and2  gate429(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate430(.a(s_32), .O(gate190inter3));
  inv1  gate431(.a(s_33), .O(gate190inter4));
  nand2 gate432(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate433(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate434(.a(N77), .O(gate190inter7));
  inv1  gate435(.a(N711), .O(gate190inter8));
  nand2 gate436(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate437(.a(s_33), .b(gate190inter3), .O(gate190inter10));
  nor2  gate438(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate439(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate440(.a(gate190inter12), .b(gate190inter1), .O(N743));
xor2 gate191( .a(N81), .b(N712), .O(N744) );

  xor2  gate595(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate596(.a(gate192inter0), .b(s_56), .O(gate192inter1));
  and2  gate597(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate598(.a(s_56), .O(gate192inter3));
  inv1  gate599(.a(s_57), .O(gate192inter4));
  nand2 gate600(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate601(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate602(.a(N85), .O(gate192inter7));
  inv1  gate603(.a(N713), .O(gate192inter8));
  nand2 gate604(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate605(.a(s_57), .b(gate192inter3), .O(gate192inter10));
  nor2  gate606(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate607(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate608(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );

  xor2  gate623(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate624(.a(gate195inter0), .b(s_60), .O(gate195inter1));
  and2  gate625(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate626(.a(s_60), .O(gate195inter3));
  inv1  gate627(.a(s_61), .O(gate195inter4));
  nand2 gate628(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate629(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate630(.a(N97), .O(gate195inter7));
  inv1  gate631(.a(N716), .O(gate195inter8));
  nand2 gate632(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate633(.a(s_61), .b(gate195inter3), .O(gate195inter10));
  nor2  gate634(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate635(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate636(.a(gate195inter12), .b(gate195inter1), .O(N748));
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule