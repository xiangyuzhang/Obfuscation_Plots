module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2409(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2410(.a(gate12inter0), .b(s_266), .O(gate12inter1));
  and2  gate2411(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2412(.a(s_266), .O(gate12inter3));
  inv1  gate2413(.a(s_267), .O(gate12inter4));
  nand2 gate2414(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2415(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2416(.a(G7), .O(gate12inter7));
  inv1  gate2417(.a(G8), .O(gate12inter8));
  nand2 gate2418(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2419(.a(s_267), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2420(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2421(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2422(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2255(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2256(.a(gate14inter0), .b(s_244), .O(gate14inter1));
  and2  gate2257(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2258(.a(s_244), .O(gate14inter3));
  inv1  gate2259(.a(s_245), .O(gate14inter4));
  nand2 gate2260(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2261(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2262(.a(G11), .O(gate14inter7));
  inv1  gate2263(.a(G12), .O(gate14inter8));
  nand2 gate2264(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2265(.a(s_245), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2266(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2267(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2268(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2381(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2382(.a(gate16inter0), .b(s_262), .O(gate16inter1));
  and2  gate2383(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2384(.a(s_262), .O(gate16inter3));
  inv1  gate2385(.a(s_263), .O(gate16inter4));
  nand2 gate2386(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2387(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2388(.a(G15), .O(gate16inter7));
  inv1  gate2389(.a(G16), .O(gate16inter8));
  nand2 gate2390(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2391(.a(s_263), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2392(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2393(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2394(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate925(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate926(.a(gate17inter0), .b(s_54), .O(gate17inter1));
  and2  gate927(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate928(.a(s_54), .O(gate17inter3));
  inv1  gate929(.a(s_55), .O(gate17inter4));
  nand2 gate930(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate931(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate932(.a(G17), .O(gate17inter7));
  inv1  gate933(.a(G18), .O(gate17inter8));
  nand2 gate934(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate935(.a(s_55), .b(gate17inter3), .O(gate17inter10));
  nor2  gate936(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate937(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate938(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2787(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2788(.a(gate26inter0), .b(s_320), .O(gate26inter1));
  and2  gate2789(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2790(.a(s_320), .O(gate26inter3));
  inv1  gate2791(.a(s_321), .O(gate26inter4));
  nand2 gate2792(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2793(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2794(.a(G9), .O(gate26inter7));
  inv1  gate2795(.a(G13), .O(gate26inter8));
  nand2 gate2796(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2797(.a(s_321), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2798(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2799(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2800(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate2157(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2158(.a(gate27inter0), .b(s_230), .O(gate27inter1));
  and2  gate2159(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2160(.a(s_230), .O(gate27inter3));
  inv1  gate2161(.a(s_231), .O(gate27inter4));
  nand2 gate2162(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2163(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2164(.a(G2), .O(gate27inter7));
  inv1  gate2165(.a(G6), .O(gate27inter8));
  nand2 gate2166(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2167(.a(s_231), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2168(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2169(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2170(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate2479(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2480(.a(gate28inter0), .b(s_276), .O(gate28inter1));
  and2  gate2481(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2482(.a(s_276), .O(gate28inter3));
  inv1  gate2483(.a(s_277), .O(gate28inter4));
  nand2 gate2484(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2485(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2486(.a(G10), .O(gate28inter7));
  inv1  gate2487(.a(G14), .O(gate28inter8));
  nand2 gate2488(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2489(.a(s_277), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2490(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2491(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2492(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2885(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2886(.a(gate33inter0), .b(s_334), .O(gate33inter1));
  and2  gate2887(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2888(.a(s_334), .O(gate33inter3));
  inv1  gate2889(.a(s_335), .O(gate33inter4));
  nand2 gate2890(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2891(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2892(.a(G17), .O(gate33inter7));
  inv1  gate2893(.a(G21), .O(gate33inter8));
  nand2 gate2894(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2895(.a(s_335), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2896(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2897(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2898(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2227(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2228(.a(gate34inter0), .b(s_240), .O(gate34inter1));
  and2  gate2229(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2230(.a(s_240), .O(gate34inter3));
  inv1  gate2231(.a(s_241), .O(gate34inter4));
  nand2 gate2232(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2233(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2234(.a(G25), .O(gate34inter7));
  inv1  gate2235(.a(G29), .O(gate34inter8));
  nand2 gate2236(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2237(.a(s_241), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2238(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2239(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2240(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate2759(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2760(.a(gate35inter0), .b(s_316), .O(gate35inter1));
  and2  gate2761(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2762(.a(s_316), .O(gate35inter3));
  inv1  gate2763(.a(s_317), .O(gate35inter4));
  nand2 gate2764(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2765(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2766(.a(G18), .O(gate35inter7));
  inv1  gate2767(.a(G22), .O(gate35inter8));
  nand2 gate2768(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2769(.a(s_317), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2770(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2771(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2772(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1737(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1738(.a(gate36inter0), .b(s_170), .O(gate36inter1));
  and2  gate1739(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1740(.a(s_170), .O(gate36inter3));
  inv1  gate1741(.a(s_171), .O(gate36inter4));
  nand2 gate1742(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1743(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1744(.a(G26), .O(gate36inter7));
  inv1  gate1745(.a(G30), .O(gate36inter8));
  nand2 gate1746(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1747(.a(s_171), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1748(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1749(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1750(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1723(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1724(.a(gate38inter0), .b(s_168), .O(gate38inter1));
  and2  gate1725(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1726(.a(s_168), .O(gate38inter3));
  inv1  gate1727(.a(s_169), .O(gate38inter4));
  nand2 gate1728(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1729(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1730(.a(G27), .O(gate38inter7));
  inv1  gate1731(.a(G31), .O(gate38inter8));
  nand2 gate1732(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1733(.a(s_169), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1734(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1735(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1736(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1807(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1808(.a(gate39inter0), .b(s_180), .O(gate39inter1));
  and2  gate1809(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1810(.a(s_180), .O(gate39inter3));
  inv1  gate1811(.a(s_181), .O(gate39inter4));
  nand2 gate1812(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1813(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1814(.a(G20), .O(gate39inter7));
  inv1  gate1815(.a(G24), .O(gate39inter8));
  nand2 gate1816(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1817(.a(s_181), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1818(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1819(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1820(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2843(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2844(.a(gate42inter0), .b(s_328), .O(gate42inter1));
  and2  gate2845(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2846(.a(s_328), .O(gate42inter3));
  inv1  gate2847(.a(s_329), .O(gate42inter4));
  nand2 gate2848(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2849(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2850(.a(G2), .O(gate42inter7));
  inv1  gate2851(.a(G266), .O(gate42inter8));
  nand2 gate2852(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2853(.a(s_329), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2854(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2855(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2856(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate785(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate786(.a(gate44inter0), .b(s_34), .O(gate44inter1));
  and2  gate787(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate788(.a(s_34), .O(gate44inter3));
  inv1  gate789(.a(s_35), .O(gate44inter4));
  nand2 gate790(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate791(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate792(.a(G4), .O(gate44inter7));
  inv1  gate793(.a(G269), .O(gate44inter8));
  nand2 gate794(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate795(.a(s_35), .b(gate44inter3), .O(gate44inter10));
  nor2  gate796(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate797(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate798(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2549(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2550(.a(gate47inter0), .b(s_286), .O(gate47inter1));
  and2  gate2551(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2552(.a(s_286), .O(gate47inter3));
  inv1  gate2553(.a(s_287), .O(gate47inter4));
  nand2 gate2554(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2555(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2556(.a(G7), .O(gate47inter7));
  inv1  gate2557(.a(G275), .O(gate47inter8));
  nand2 gate2558(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2559(.a(s_287), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2560(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2561(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2562(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1359(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1360(.a(gate48inter0), .b(s_116), .O(gate48inter1));
  and2  gate1361(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1362(.a(s_116), .O(gate48inter3));
  inv1  gate1363(.a(s_117), .O(gate48inter4));
  nand2 gate1364(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1365(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1366(.a(G8), .O(gate48inter7));
  inv1  gate1367(.a(G275), .O(gate48inter8));
  nand2 gate1368(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1369(.a(s_117), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1370(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1371(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1372(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1793(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1794(.a(gate49inter0), .b(s_178), .O(gate49inter1));
  and2  gate1795(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1796(.a(s_178), .O(gate49inter3));
  inv1  gate1797(.a(s_179), .O(gate49inter4));
  nand2 gate1798(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1799(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1800(.a(G9), .O(gate49inter7));
  inv1  gate1801(.a(G278), .O(gate49inter8));
  nand2 gate1802(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1803(.a(s_179), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1804(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1805(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1806(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1849(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1850(.a(gate54inter0), .b(s_186), .O(gate54inter1));
  and2  gate1851(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1852(.a(s_186), .O(gate54inter3));
  inv1  gate1853(.a(s_187), .O(gate54inter4));
  nand2 gate1854(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1855(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1856(.a(G14), .O(gate54inter7));
  inv1  gate1857(.a(G284), .O(gate54inter8));
  nand2 gate1858(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1859(.a(s_187), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1860(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1861(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1862(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate2059(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2060(.a(gate55inter0), .b(s_216), .O(gate55inter1));
  and2  gate2061(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2062(.a(s_216), .O(gate55inter3));
  inv1  gate2063(.a(s_217), .O(gate55inter4));
  nand2 gate2064(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2065(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2066(.a(G15), .O(gate55inter7));
  inv1  gate2067(.a(G287), .O(gate55inter8));
  nand2 gate2068(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2069(.a(s_217), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2070(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2071(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2072(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1429(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1430(.a(gate56inter0), .b(s_126), .O(gate56inter1));
  and2  gate1431(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1432(.a(s_126), .O(gate56inter3));
  inv1  gate1433(.a(s_127), .O(gate56inter4));
  nand2 gate1434(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1435(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1436(.a(G16), .O(gate56inter7));
  inv1  gate1437(.a(G287), .O(gate56inter8));
  nand2 gate1438(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1439(.a(s_127), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1440(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1441(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1442(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2955(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2956(.a(gate60inter0), .b(s_344), .O(gate60inter1));
  and2  gate2957(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2958(.a(s_344), .O(gate60inter3));
  inv1  gate2959(.a(s_345), .O(gate60inter4));
  nand2 gate2960(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2961(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2962(.a(G20), .O(gate60inter7));
  inv1  gate2963(.a(G293), .O(gate60inter8));
  nand2 gate2964(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2965(.a(s_345), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2966(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2967(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2968(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2857(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2858(.a(gate62inter0), .b(s_330), .O(gate62inter1));
  and2  gate2859(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2860(.a(s_330), .O(gate62inter3));
  inv1  gate2861(.a(s_331), .O(gate62inter4));
  nand2 gate2862(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2863(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2864(.a(G22), .O(gate62inter7));
  inv1  gate2865(.a(G296), .O(gate62inter8));
  nand2 gate2866(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2867(.a(s_331), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2868(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2869(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2870(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2199(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2200(.a(gate63inter0), .b(s_236), .O(gate63inter1));
  and2  gate2201(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2202(.a(s_236), .O(gate63inter3));
  inv1  gate2203(.a(s_237), .O(gate63inter4));
  nand2 gate2204(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2205(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2206(.a(G23), .O(gate63inter7));
  inv1  gate2207(.a(G299), .O(gate63inter8));
  nand2 gate2208(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2209(.a(s_237), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2210(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2211(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2212(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2507(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2508(.a(gate67inter0), .b(s_280), .O(gate67inter1));
  and2  gate2509(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2510(.a(s_280), .O(gate67inter3));
  inv1  gate2511(.a(s_281), .O(gate67inter4));
  nand2 gate2512(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2513(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2514(.a(G27), .O(gate67inter7));
  inv1  gate2515(.a(G305), .O(gate67inter8));
  nand2 gate2516(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2517(.a(s_281), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2518(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2519(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2520(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1821(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1822(.a(gate69inter0), .b(s_182), .O(gate69inter1));
  and2  gate1823(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1824(.a(s_182), .O(gate69inter3));
  inv1  gate1825(.a(s_183), .O(gate69inter4));
  nand2 gate1826(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1827(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1828(.a(G29), .O(gate69inter7));
  inv1  gate1829(.a(G308), .O(gate69inter8));
  nand2 gate1830(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1831(.a(s_183), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1832(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1833(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1834(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate2101(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2102(.a(gate75inter0), .b(s_222), .O(gate75inter1));
  and2  gate2103(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2104(.a(s_222), .O(gate75inter3));
  inv1  gate2105(.a(s_223), .O(gate75inter4));
  nand2 gate2106(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2107(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2108(.a(G9), .O(gate75inter7));
  inv1  gate2109(.a(G317), .O(gate75inter8));
  nand2 gate2110(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2111(.a(s_223), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2112(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2113(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2114(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1485(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1486(.a(gate76inter0), .b(s_134), .O(gate76inter1));
  and2  gate1487(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1488(.a(s_134), .O(gate76inter3));
  inv1  gate1489(.a(s_135), .O(gate76inter4));
  nand2 gate1490(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1491(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1492(.a(G13), .O(gate76inter7));
  inv1  gate1493(.a(G317), .O(gate76inter8));
  nand2 gate1494(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1495(.a(s_135), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1496(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1497(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1498(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1065(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1066(.a(gate79inter0), .b(s_74), .O(gate79inter1));
  and2  gate1067(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1068(.a(s_74), .O(gate79inter3));
  inv1  gate1069(.a(s_75), .O(gate79inter4));
  nand2 gate1070(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1071(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1072(.a(G10), .O(gate79inter7));
  inv1  gate1073(.a(G323), .O(gate79inter8));
  nand2 gate1074(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1075(.a(s_75), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1076(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1077(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1078(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate855(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate856(.a(gate80inter0), .b(s_44), .O(gate80inter1));
  and2  gate857(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate858(.a(s_44), .O(gate80inter3));
  inv1  gate859(.a(s_45), .O(gate80inter4));
  nand2 gate860(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate861(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate862(.a(G14), .O(gate80inter7));
  inv1  gate863(.a(G323), .O(gate80inter8));
  nand2 gate864(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate865(.a(s_45), .b(gate80inter3), .O(gate80inter10));
  nor2  gate866(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate867(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate868(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate547(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate548(.a(gate81inter0), .b(s_0), .O(gate81inter1));
  and2  gate549(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate550(.a(s_0), .O(gate81inter3));
  inv1  gate551(.a(s_1), .O(gate81inter4));
  nand2 gate552(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate553(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate554(.a(G3), .O(gate81inter7));
  inv1  gate555(.a(G326), .O(gate81inter8));
  nand2 gate556(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate557(.a(s_1), .b(gate81inter3), .O(gate81inter10));
  nor2  gate558(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate559(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate560(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2633(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2634(.a(gate88inter0), .b(s_298), .O(gate88inter1));
  and2  gate2635(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2636(.a(s_298), .O(gate88inter3));
  inv1  gate2637(.a(s_299), .O(gate88inter4));
  nand2 gate2638(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2639(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2640(.a(G16), .O(gate88inter7));
  inv1  gate2641(.a(G335), .O(gate88inter8));
  nand2 gate2642(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2643(.a(s_299), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2644(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2645(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2646(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate631(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate632(.a(gate89inter0), .b(s_12), .O(gate89inter1));
  and2  gate633(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate634(.a(s_12), .O(gate89inter3));
  inv1  gate635(.a(s_13), .O(gate89inter4));
  nand2 gate636(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate637(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate638(.a(G17), .O(gate89inter7));
  inv1  gate639(.a(G338), .O(gate89inter8));
  nand2 gate640(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate641(.a(s_13), .b(gate89inter3), .O(gate89inter10));
  nor2  gate642(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate643(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate644(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1317(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1318(.a(gate90inter0), .b(s_110), .O(gate90inter1));
  and2  gate1319(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1320(.a(s_110), .O(gate90inter3));
  inv1  gate1321(.a(s_111), .O(gate90inter4));
  nand2 gate1322(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1323(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1324(.a(G21), .O(gate90inter7));
  inv1  gate1325(.a(G338), .O(gate90inter8));
  nand2 gate1326(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1327(.a(s_111), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1328(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1329(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1330(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate841(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate842(.a(gate91inter0), .b(s_42), .O(gate91inter1));
  and2  gate843(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate844(.a(s_42), .O(gate91inter3));
  inv1  gate845(.a(s_43), .O(gate91inter4));
  nand2 gate846(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate847(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate848(.a(G25), .O(gate91inter7));
  inv1  gate849(.a(G341), .O(gate91inter8));
  nand2 gate850(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate851(.a(s_43), .b(gate91inter3), .O(gate91inter10));
  nor2  gate852(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate853(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate854(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2717(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2718(.a(gate92inter0), .b(s_310), .O(gate92inter1));
  and2  gate2719(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2720(.a(s_310), .O(gate92inter3));
  inv1  gate2721(.a(s_311), .O(gate92inter4));
  nand2 gate2722(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2723(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2724(.a(G29), .O(gate92inter7));
  inv1  gate2725(.a(G341), .O(gate92inter8));
  nand2 gate2726(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2727(.a(s_311), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2728(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2729(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2730(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1597(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1598(.a(gate94inter0), .b(s_150), .O(gate94inter1));
  and2  gate1599(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1600(.a(s_150), .O(gate94inter3));
  inv1  gate1601(.a(s_151), .O(gate94inter4));
  nand2 gate1602(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1603(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1604(.a(G22), .O(gate94inter7));
  inv1  gate1605(.a(G344), .O(gate94inter8));
  nand2 gate1606(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1607(.a(s_151), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1608(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1609(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1610(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2395(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2396(.a(gate100inter0), .b(s_264), .O(gate100inter1));
  and2  gate2397(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2398(.a(s_264), .O(gate100inter3));
  inv1  gate2399(.a(s_265), .O(gate100inter4));
  nand2 gate2400(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2401(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2402(.a(G31), .O(gate100inter7));
  inv1  gate2403(.a(G353), .O(gate100inter8));
  nand2 gate2404(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2405(.a(s_265), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2406(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2407(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2408(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1261(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1262(.a(gate103inter0), .b(s_102), .O(gate103inter1));
  and2  gate1263(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1264(.a(s_102), .O(gate103inter3));
  inv1  gate1265(.a(s_103), .O(gate103inter4));
  nand2 gate1266(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1267(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1268(.a(G28), .O(gate103inter7));
  inv1  gate1269(.a(G359), .O(gate103inter8));
  nand2 gate1270(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1271(.a(s_103), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1272(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1273(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1274(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1835(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1836(.a(gate105inter0), .b(s_184), .O(gate105inter1));
  and2  gate1837(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1838(.a(s_184), .O(gate105inter3));
  inv1  gate1839(.a(s_185), .O(gate105inter4));
  nand2 gate1840(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1841(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1842(.a(G362), .O(gate105inter7));
  inv1  gate1843(.a(G363), .O(gate105inter8));
  nand2 gate1844(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1845(.a(s_185), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1846(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1847(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1848(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate995(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate996(.a(gate106inter0), .b(s_64), .O(gate106inter1));
  and2  gate997(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate998(.a(s_64), .O(gate106inter3));
  inv1  gate999(.a(s_65), .O(gate106inter4));
  nand2 gate1000(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1001(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1002(.a(G364), .O(gate106inter7));
  inv1  gate1003(.a(G365), .O(gate106inter8));
  nand2 gate1004(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1005(.a(s_65), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1006(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1007(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1008(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2997(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2998(.a(gate110inter0), .b(s_350), .O(gate110inter1));
  and2  gate2999(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate3000(.a(s_350), .O(gate110inter3));
  inv1  gate3001(.a(s_351), .O(gate110inter4));
  nand2 gate3002(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate3003(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate3004(.a(G372), .O(gate110inter7));
  inv1  gate3005(.a(G373), .O(gate110inter8));
  nand2 gate3006(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate3007(.a(s_351), .b(gate110inter3), .O(gate110inter10));
  nor2  gate3008(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate3009(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate3010(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2745(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2746(.a(gate112inter0), .b(s_314), .O(gate112inter1));
  and2  gate2747(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2748(.a(s_314), .O(gate112inter3));
  inv1  gate2749(.a(s_315), .O(gate112inter4));
  nand2 gate2750(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2751(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2752(.a(G376), .O(gate112inter7));
  inv1  gate2753(.a(G377), .O(gate112inter8));
  nand2 gate2754(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2755(.a(s_315), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2756(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2757(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2758(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1191(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1192(.a(gate113inter0), .b(s_92), .O(gate113inter1));
  and2  gate1193(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1194(.a(s_92), .O(gate113inter3));
  inv1  gate1195(.a(s_93), .O(gate113inter4));
  nand2 gate1196(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1197(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1198(.a(G378), .O(gate113inter7));
  inv1  gate1199(.a(G379), .O(gate113inter8));
  nand2 gate1200(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1201(.a(s_93), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1202(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1203(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1204(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1205(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1206(.a(gate115inter0), .b(s_94), .O(gate115inter1));
  and2  gate1207(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1208(.a(s_94), .O(gate115inter3));
  inv1  gate1209(.a(s_95), .O(gate115inter4));
  nand2 gate1210(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1211(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1212(.a(G382), .O(gate115inter7));
  inv1  gate1213(.a(G383), .O(gate115inter8));
  nand2 gate1214(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1215(.a(s_95), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1216(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1217(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1218(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2297(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2298(.a(gate120inter0), .b(s_250), .O(gate120inter1));
  and2  gate2299(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2300(.a(s_250), .O(gate120inter3));
  inv1  gate2301(.a(s_251), .O(gate120inter4));
  nand2 gate2302(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2303(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2304(.a(G392), .O(gate120inter7));
  inv1  gate2305(.a(G393), .O(gate120inter8));
  nand2 gate2306(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2307(.a(s_251), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2308(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2309(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2310(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1163(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1164(.a(gate122inter0), .b(s_88), .O(gate122inter1));
  and2  gate1165(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1166(.a(s_88), .O(gate122inter3));
  inv1  gate1167(.a(s_89), .O(gate122inter4));
  nand2 gate1168(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1169(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1170(.a(G396), .O(gate122inter7));
  inv1  gate1171(.a(G397), .O(gate122inter8));
  nand2 gate1172(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1173(.a(s_89), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1174(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1175(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1176(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1555(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1556(.a(gate123inter0), .b(s_144), .O(gate123inter1));
  and2  gate1557(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1558(.a(s_144), .O(gate123inter3));
  inv1  gate1559(.a(s_145), .O(gate123inter4));
  nand2 gate1560(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1561(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1562(.a(G398), .O(gate123inter7));
  inv1  gate1563(.a(G399), .O(gate123inter8));
  nand2 gate1564(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1565(.a(s_145), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1566(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1567(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1568(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate2871(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2872(.a(gate124inter0), .b(s_332), .O(gate124inter1));
  and2  gate2873(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2874(.a(s_332), .O(gate124inter3));
  inv1  gate2875(.a(s_333), .O(gate124inter4));
  nand2 gate2876(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2877(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2878(.a(G400), .O(gate124inter7));
  inv1  gate2879(.a(G401), .O(gate124inter8));
  nand2 gate2880(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2881(.a(s_333), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2882(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2883(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2884(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate2675(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2676(.a(gate125inter0), .b(s_304), .O(gate125inter1));
  and2  gate2677(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2678(.a(s_304), .O(gate125inter3));
  inv1  gate2679(.a(s_305), .O(gate125inter4));
  nand2 gate2680(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2681(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2682(.a(G402), .O(gate125inter7));
  inv1  gate2683(.a(G403), .O(gate125inter8));
  nand2 gate2684(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2685(.a(s_305), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2686(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2687(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2688(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1331(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1332(.a(gate126inter0), .b(s_112), .O(gate126inter1));
  and2  gate1333(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1334(.a(s_112), .O(gate126inter3));
  inv1  gate1335(.a(s_113), .O(gate126inter4));
  nand2 gate1336(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1337(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1338(.a(G404), .O(gate126inter7));
  inv1  gate1339(.a(G405), .O(gate126inter8));
  nand2 gate1340(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1341(.a(s_113), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1342(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1343(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1344(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate911(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate912(.a(gate129inter0), .b(s_52), .O(gate129inter1));
  and2  gate913(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate914(.a(s_52), .O(gate129inter3));
  inv1  gate915(.a(s_53), .O(gate129inter4));
  nand2 gate916(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate917(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate918(.a(G410), .O(gate129inter7));
  inv1  gate919(.a(G411), .O(gate129inter8));
  nand2 gate920(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate921(.a(s_53), .b(gate129inter3), .O(gate129inter10));
  nor2  gate922(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate923(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate924(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2605(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2606(.a(gate130inter0), .b(s_294), .O(gate130inter1));
  and2  gate2607(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2608(.a(s_294), .O(gate130inter3));
  inv1  gate2609(.a(s_295), .O(gate130inter4));
  nand2 gate2610(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2611(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2612(.a(G412), .O(gate130inter7));
  inv1  gate2613(.a(G413), .O(gate130inter8));
  nand2 gate2614(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2615(.a(s_295), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2616(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2617(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2618(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate799(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate800(.a(gate132inter0), .b(s_36), .O(gate132inter1));
  and2  gate801(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate802(.a(s_36), .O(gate132inter3));
  inv1  gate803(.a(s_37), .O(gate132inter4));
  nand2 gate804(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate805(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate806(.a(G416), .O(gate132inter7));
  inv1  gate807(.a(G417), .O(gate132inter8));
  nand2 gate808(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate809(.a(s_37), .b(gate132inter3), .O(gate132inter10));
  nor2  gate810(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate811(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate812(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate869(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate870(.a(gate134inter0), .b(s_46), .O(gate134inter1));
  and2  gate871(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate872(.a(s_46), .O(gate134inter3));
  inv1  gate873(.a(s_47), .O(gate134inter4));
  nand2 gate874(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate875(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate876(.a(G420), .O(gate134inter7));
  inv1  gate877(.a(G421), .O(gate134inter8));
  nand2 gate878(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate879(.a(s_47), .b(gate134inter3), .O(gate134inter10));
  nor2  gate880(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate881(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate882(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2269(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2270(.a(gate139inter0), .b(s_246), .O(gate139inter1));
  and2  gate2271(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2272(.a(s_246), .O(gate139inter3));
  inv1  gate2273(.a(s_247), .O(gate139inter4));
  nand2 gate2274(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2275(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2276(.a(G438), .O(gate139inter7));
  inv1  gate2277(.a(G441), .O(gate139inter8));
  nand2 gate2278(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2279(.a(s_247), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2280(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2281(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2282(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate939(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate940(.a(gate144inter0), .b(s_56), .O(gate144inter1));
  and2  gate941(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate942(.a(s_56), .O(gate144inter3));
  inv1  gate943(.a(s_57), .O(gate144inter4));
  nand2 gate944(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate945(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate946(.a(G468), .O(gate144inter7));
  inv1  gate947(.a(G471), .O(gate144inter8));
  nand2 gate948(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate949(.a(s_57), .b(gate144inter3), .O(gate144inter10));
  nor2  gate950(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate951(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate952(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2031(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2032(.a(gate151inter0), .b(s_212), .O(gate151inter1));
  and2  gate2033(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2034(.a(s_212), .O(gate151inter3));
  inv1  gate2035(.a(s_213), .O(gate151inter4));
  nand2 gate2036(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2037(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2038(.a(G510), .O(gate151inter7));
  inv1  gate2039(.a(G513), .O(gate151inter8));
  nand2 gate2040(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2041(.a(s_213), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2042(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2043(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2044(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2129(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2130(.a(gate154inter0), .b(s_226), .O(gate154inter1));
  and2  gate2131(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2132(.a(s_226), .O(gate154inter3));
  inv1  gate2133(.a(s_227), .O(gate154inter4));
  nand2 gate2134(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2135(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2136(.a(G429), .O(gate154inter7));
  inv1  gate2137(.a(G522), .O(gate154inter8));
  nand2 gate2138(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2139(.a(s_227), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2140(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2141(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2142(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1387(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1388(.a(gate155inter0), .b(s_120), .O(gate155inter1));
  and2  gate1389(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1390(.a(s_120), .O(gate155inter3));
  inv1  gate1391(.a(s_121), .O(gate155inter4));
  nand2 gate1392(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1393(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1394(.a(G432), .O(gate155inter7));
  inv1  gate1395(.a(G525), .O(gate155inter8));
  nand2 gate1396(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1397(.a(s_121), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1398(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1399(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1400(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate589(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate590(.a(gate157inter0), .b(s_6), .O(gate157inter1));
  and2  gate591(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate592(.a(s_6), .O(gate157inter3));
  inv1  gate593(.a(s_7), .O(gate157inter4));
  nand2 gate594(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate595(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate596(.a(G438), .O(gate157inter7));
  inv1  gate597(.a(G528), .O(gate157inter8));
  nand2 gate598(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate599(.a(s_7), .b(gate157inter3), .O(gate157inter10));
  nor2  gate600(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate601(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate602(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate771(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate772(.a(gate158inter0), .b(s_32), .O(gate158inter1));
  and2  gate773(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate774(.a(s_32), .O(gate158inter3));
  inv1  gate775(.a(s_33), .O(gate158inter4));
  nand2 gate776(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate777(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate778(.a(G441), .O(gate158inter7));
  inv1  gate779(.a(G528), .O(gate158inter8));
  nand2 gate780(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate781(.a(s_33), .b(gate158inter3), .O(gate158inter10));
  nor2  gate782(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate783(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate784(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1303(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1304(.a(gate160inter0), .b(s_108), .O(gate160inter1));
  and2  gate1305(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1306(.a(s_108), .O(gate160inter3));
  inv1  gate1307(.a(s_109), .O(gate160inter4));
  nand2 gate1308(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1309(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1310(.a(G447), .O(gate160inter7));
  inv1  gate1311(.a(G531), .O(gate160inter8));
  nand2 gate1312(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1313(.a(s_109), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1314(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1315(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1316(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1863(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1864(.a(gate162inter0), .b(s_188), .O(gate162inter1));
  and2  gate1865(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1866(.a(s_188), .O(gate162inter3));
  inv1  gate1867(.a(s_189), .O(gate162inter4));
  nand2 gate1868(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1869(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1870(.a(G453), .O(gate162inter7));
  inv1  gate1871(.a(G534), .O(gate162inter8));
  nand2 gate1872(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1873(.a(s_189), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1874(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1875(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1876(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate953(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate954(.a(gate168inter0), .b(s_58), .O(gate168inter1));
  and2  gate955(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate956(.a(s_58), .O(gate168inter3));
  inv1  gate957(.a(s_59), .O(gate168inter4));
  nand2 gate958(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate959(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate960(.a(G471), .O(gate168inter7));
  inv1  gate961(.a(G543), .O(gate168inter8));
  nand2 gate962(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate963(.a(s_59), .b(gate168inter3), .O(gate168inter10));
  nor2  gate964(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate965(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate966(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate813(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate814(.a(gate170inter0), .b(s_38), .O(gate170inter1));
  and2  gate815(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate816(.a(s_38), .O(gate170inter3));
  inv1  gate817(.a(s_39), .O(gate170inter4));
  nand2 gate818(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate819(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate820(.a(G477), .O(gate170inter7));
  inv1  gate821(.a(G546), .O(gate170inter8));
  nand2 gate822(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate823(.a(s_39), .b(gate170inter3), .O(gate170inter10));
  nor2  gate824(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate825(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate826(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2815(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2816(.a(gate174inter0), .b(s_324), .O(gate174inter1));
  and2  gate2817(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2818(.a(s_324), .O(gate174inter3));
  inv1  gate2819(.a(s_325), .O(gate174inter4));
  nand2 gate2820(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2821(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2822(.a(G489), .O(gate174inter7));
  inv1  gate2823(.a(G552), .O(gate174inter8));
  nand2 gate2824(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2825(.a(s_325), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2826(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2827(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2828(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1177(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1178(.a(gate177inter0), .b(s_90), .O(gate177inter1));
  and2  gate1179(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1180(.a(s_90), .O(gate177inter3));
  inv1  gate1181(.a(s_91), .O(gate177inter4));
  nand2 gate1182(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1183(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1184(.a(G498), .O(gate177inter7));
  inv1  gate1185(.a(G558), .O(gate177inter8));
  nand2 gate1186(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1187(.a(s_91), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1188(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1189(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1190(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2703(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2704(.a(gate179inter0), .b(s_308), .O(gate179inter1));
  and2  gate2705(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2706(.a(s_308), .O(gate179inter3));
  inv1  gate2707(.a(s_309), .O(gate179inter4));
  nand2 gate2708(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2709(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2710(.a(G504), .O(gate179inter7));
  inv1  gate2711(.a(G561), .O(gate179inter8));
  nand2 gate2712(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2713(.a(s_309), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2714(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2715(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2716(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1093(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1094(.a(gate180inter0), .b(s_78), .O(gate180inter1));
  and2  gate1095(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1096(.a(s_78), .O(gate180inter3));
  inv1  gate1097(.a(s_79), .O(gate180inter4));
  nand2 gate1098(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1099(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1100(.a(G507), .O(gate180inter7));
  inv1  gate1101(.a(G561), .O(gate180inter8));
  nand2 gate1102(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1103(.a(s_79), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1104(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1105(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1106(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1569(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1570(.a(gate181inter0), .b(s_146), .O(gate181inter1));
  and2  gate1571(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1572(.a(s_146), .O(gate181inter3));
  inv1  gate1573(.a(s_147), .O(gate181inter4));
  nand2 gate1574(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1575(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1576(.a(G510), .O(gate181inter7));
  inv1  gate1577(.a(G564), .O(gate181inter8));
  nand2 gate1578(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1579(.a(s_147), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1580(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1581(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1582(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2087(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2088(.a(gate182inter0), .b(s_220), .O(gate182inter1));
  and2  gate2089(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2090(.a(s_220), .O(gate182inter3));
  inv1  gate2091(.a(s_221), .O(gate182inter4));
  nand2 gate2092(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2093(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2094(.a(G513), .O(gate182inter7));
  inv1  gate2095(.a(G564), .O(gate182inter8));
  nand2 gate2096(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2097(.a(s_221), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2098(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2099(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2100(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2577(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2578(.a(gate184inter0), .b(s_290), .O(gate184inter1));
  and2  gate2579(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2580(.a(s_290), .O(gate184inter3));
  inv1  gate2581(.a(s_291), .O(gate184inter4));
  nand2 gate2582(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2583(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2584(.a(G519), .O(gate184inter7));
  inv1  gate2585(.a(G567), .O(gate184inter8));
  nand2 gate2586(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2587(.a(s_291), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2588(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2589(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2590(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1471(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1472(.a(gate185inter0), .b(s_132), .O(gate185inter1));
  and2  gate1473(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1474(.a(s_132), .O(gate185inter3));
  inv1  gate1475(.a(s_133), .O(gate185inter4));
  nand2 gate1476(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1477(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1478(.a(G570), .O(gate185inter7));
  inv1  gate1479(.a(G571), .O(gate185inter8));
  nand2 gate1480(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1481(.a(s_133), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1482(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1483(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1484(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate883(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate884(.a(gate186inter0), .b(s_48), .O(gate186inter1));
  and2  gate885(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate886(.a(s_48), .O(gate186inter3));
  inv1  gate887(.a(s_49), .O(gate186inter4));
  nand2 gate888(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate889(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate890(.a(G572), .O(gate186inter7));
  inv1  gate891(.a(G573), .O(gate186inter8));
  nand2 gate892(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate893(.a(s_49), .b(gate186inter3), .O(gate186inter10));
  nor2  gate894(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate895(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate896(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate743(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate744(.a(gate188inter0), .b(s_28), .O(gate188inter1));
  and2  gate745(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate746(.a(s_28), .O(gate188inter3));
  inv1  gate747(.a(s_29), .O(gate188inter4));
  nand2 gate748(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate749(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate750(.a(G576), .O(gate188inter7));
  inv1  gate751(.a(G577), .O(gate188inter8));
  nand2 gate752(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate753(.a(s_29), .b(gate188inter3), .O(gate188inter10));
  nor2  gate754(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate755(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate756(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1121(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1122(.a(gate190inter0), .b(s_82), .O(gate190inter1));
  and2  gate1123(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1124(.a(s_82), .O(gate190inter3));
  inv1  gate1125(.a(s_83), .O(gate190inter4));
  nand2 gate1126(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1127(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1128(.a(G580), .O(gate190inter7));
  inv1  gate1129(.a(G581), .O(gate190inter8));
  nand2 gate1130(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1131(.a(s_83), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1132(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1133(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1134(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2003(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2004(.a(gate191inter0), .b(s_208), .O(gate191inter1));
  and2  gate2005(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2006(.a(s_208), .O(gate191inter3));
  inv1  gate2007(.a(s_209), .O(gate191inter4));
  nand2 gate2008(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2009(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2010(.a(G582), .O(gate191inter7));
  inv1  gate2011(.a(G583), .O(gate191inter8));
  nand2 gate2012(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2013(.a(s_209), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2014(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2015(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2016(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1149(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1150(.a(gate194inter0), .b(s_86), .O(gate194inter1));
  and2  gate1151(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1152(.a(s_86), .O(gate194inter3));
  inv1  gate1153(.a(s_87), .O(gate194inter4));
  nand2 gate1154(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1155(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1156(.a(G588), .O(gate194inter7));
  inv1  gate1157(.a(G589), .O(gate194inter8));
  nand2 gate1158(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1159(.a(s_87), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1160(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1161(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1162(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate603(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate604(.a(gate196inter0), .b(s_8), .O(gate196inter1));
  and2  gate605(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate606(.a(s_8), .O(gate196inter3));
  inv1  gate607(.a(s_9), .O(gate196inter4));
  nand2 gate608(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate609(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate610(.a(G592), .O(gate196inter7));
  inv1  gate611(.a(G593), .O(gate196inter8));
  nand2 gate612(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate613(.a(s_9), .b(gate196inter3), .O(gate196inter10));
  nor2  gate614(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate615(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate616(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate2535(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2536(.a(gate197inter0), .b(s_284), .O(gate197inter1));
  and2  gate2537(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2538(.a(s_284), .O(gate197inter3));
  inv1  gate2539(.a(s_285), .O(gate197inter4));
  nand2 gate2540(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2541(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2542(.a(G594), .O(gate197inter7));
  inv1  gate2543(.a(G595), .O(gate197inter8));
  nand2 gate2544(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2545(.a(s_285), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2546(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2547(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2548(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate561(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate562(.a(gate199inter0), .b(s_2), .O(gate199inter1));
  and2  gate563(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate564(.a(s_2), .O(gate199inter3));
  inv1  gate565(.a(s_3), .O(gate199inter4));
  nand2 gate566(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate567(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate568(.a(G598), .O(gate199inter7));
  inv1  gate569(.a(G599), .O(gate199inter8));
  nand2 gate570(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate571(.a(s_3), .b(gate199inter3), .O(gate199inter10));
  nor2  gate572(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate573(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate574(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate2045(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2046(.a(gate200inter0), .b(s_214), .O(gate200inter1));
  and2  gate2047(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2048(.a(s_214), .O(gate200inter3));
  inv1  gate2049(.a(s_215), .O(gate200inter4));
  nand2 gate2050(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2051(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2052(.a(G600), .O(gate200inter7));
  inv1  gate2053(.a(G601), .O(gate200inter8));
  nand2 gate2054(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2055(.a(s_215), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2056(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2057(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2058(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1779(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1780(.a(gate202inter0), .b(s_176), .O(gate202inter1));
  and2  gate1781(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1782(.a(s_176), .O(gate202inter3));
  inv1  gate1783(.a(s_177), .O(gate202inter4));
  nand2 gate1784(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1785(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1786(.a(G612), .O(gate202inter7));
  inv1  gate1787(.a(G617), .O(gate202inter8));
  nand2 gate1788(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1789(.a(s_177), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1790(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1791(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1792(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2647(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2648(.a(gate204inter0), .b(s_300), .O(gate204inter1));
  and2  gate2649(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2650(.a(s_300), .O(gate204inter3));
  inv1  gate2651(.a(s_301), .O(gate204inter4));
  nand2 gate2652(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2653(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2654(.a(G607), .O(gate204inter7));
  inv1  gate2655(.a(G617), .O(gate204inter8));
  nand2 gate2656(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2657(.a(s_301), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2658(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2659(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2660(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1961(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1962(.a(gate207inter0), .b(s_202), .O(gate207inter1));
  and2  gate1963(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1964(.a(s_202), .O(gate207inter3));
  inv1  gate1965(.a(s_203), .O(gate207inter4));
  nand2 gate1966(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1967(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1968(.a(G622), .O(gate207inter7));
  inv1  gate1969(.a(G632), .O(gate207inter8));
  nand2 gate1970(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1971(.a(s_203), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1972(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1973(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1974(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate757(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate758(.a(gate211inter0), .b(s_30), .O(gate211inter1));
  and2  gate759(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate760(.a(s_30), .O(gate211inter3));
  inv1  gate761(.a(s_31), .O(gate211inter4));
  nand2 gate762(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate763(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate764(.a(G612), .O(gate211inter7));
  inv1  gate765(.a(G669), .O(gate211inter8));
  nand2 gate766(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate767(.a(s_31), .b(gate211inter3), .O(gate211inter10));
  nor2  gate768(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate769(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate770(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate897(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate898(.a(gate212inter0), .b(s_50), .O(gate212inter1));
  and2  gate899(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate900(.a(s_50), .O(gate212inter3));
  inv1  gate901(.a(s_51), .O(gate212inter4));
  nand2 gate902(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate903(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate904(.a(G617), .O(gate212inter7));
  inv1  gate905(.a(G669), .O(gate212inter8));
  nand2 gate906(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate907(.a(s_51), .b(gate212inter3), .O(gate212inter10));
  nor2  gate908(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate909(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate910(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate659(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate660(.a(gate213inter0), .b(s_16), .O(gate213inter1));
  and2  gate661(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate662(.a(s_16), .O(gate213inter3));
  inv1  gate663(.a(s_17), .O(gate213inter4));
  nand2 gate664(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate665(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate666(.a(G602), .O(gate213inter7));
  inv1  gate667(.a(G672), .O(gate213inter8));
  nand2 gate668(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate669(.a(s_17), .b(gate213inter3), .O(gate213inter10));
  nor2  gate670(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate671(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate672(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1457(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1458(.a(gate217inter0), .b(s_130), .O(gate217inter1));
  and2  gate1459(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1460(.a(s_130), .O(gate217inter3));
  inv1  gate1461(.a(s_131), .O(gate217inter4));
  nand2 gate1462(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1463(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1464(.a(G622), .O(gate217inter7));
  inv1  gate1465(.a(G678), .O(gate217inter8));
  nand2 gate1466(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1467(.a(s_131), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1468(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1469(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1470(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2969(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2970(.a(gate220inter0), .b(s_346), .O(gate220inter1));
  and2  gate2971(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2972(.a(s_346), .O(gate220inter3));
  inv1  gate2973(.a(s_347), .O(gate220inter4));
  nand2 gate2974(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2975(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2976(.a(G637), .O(gate220inter7));
  inv1  gate2977(.a(G681), .O(gate220inter8));
  nand2 gate2978(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2979(.a(s_347), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2980(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2981(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2982(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1583(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1584(.a(gate226inter0), .b(s_148), .O(gate226inter1));
  and2  gate1585(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1586(.a(s_148), .O(gate226inter3));
  inv1  gate1587(.a(s_149), .O(gate226inter4));
  nand2 gate1588(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1589(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1590(.a(G692), .O(gate226inter7));
  inv1  gate1591(.a(G693), .O(gate226inter8));
  nand2 gate1592(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1593(.a(s_149), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1594(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1595(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1596(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1219(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1220(.a(gate235inter0), .b(s_96), .O(gate235inter1));
  and2  gate1221(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1222(.a(s_96), .O(gate235inter3));
  inv1  gate1223(.a(s_97), .O(gate235inter4));
  nand2 gate1224(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1225(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1226(.a(G248), .O(gate235inter7));
  inv1  gate1227(.a(G724), .O(gate235inter8));
  nand2 gate1228(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1229(.a(s_97), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1230(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1231(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1232(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2465(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2466(.a(gate238inter0), .b(s_274), .O(gate238inter1));
  and2  gate2467(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2468(.a(s_274), .O(gate238inter3));
  inv1  gate2469(.a(s_275), .O(gate238inter4));
  nand2 gate2470(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2471(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2472(.a(G257), .O(gate238inter7));
  inv1  gate2473(.a(G709), .O(gate238inter8));
  nand2 gate2474(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2475(.a(s_275), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2476(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2477(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2478(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1499(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1500(.a(gate244inter0), .b(s_136), .O(gate244inter1));
  and2  gate1501(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1502(.a(s_136), .O(gate244inter3));
  inv1  gate1503(.a(s_137), .O(gate244inter4));
  nand2 gate1504(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1505(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1506(.a(G721), .O(gate244inter7));
  inv1  gate1507(.a(G733), .O(gate244inter8));
  nand2 gate1508(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1509(.a(s_137), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1510(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1511(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1512(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1527(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1528(.a(gate245inter0), .b(s_140), .O(gate245inter1));
  and2  gate1529(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1530(.a(s_140), .O(gate245inter3));
  inv1  gate1531(.a(s_141), .O(gate245inter4));
  nand2 gate1532(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1533(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1534(.a(G248), .O(gate245inter7));
  inv1  gate1535(.a(G736), .O(gate245inter8));
  nand2 gate1536(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1537(.a(s_141), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1538(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1539(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1540(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1891(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1892(.a(gate246inter0), .b(s_192), .O(gate246inter1));
  and2  gate1893(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1894(.a(s_192), .O(gate246inter3));
  inv1  gate1895(.a(s_193), .O(gate246inter4));
  nand2 gate1896(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1897(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1898(.a(G724), .O(gate246inter7));
  inv1  gate1899(.a(G736), .O(gate246inter8));
  nand2 gate1900(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1901(.a(s_193), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1902(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1903(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1904(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate981(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate982(.a(gate247inter0), .b(s_62), .O(gate247inter1));
  and2  gate983(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate984(.a(s_62), .O(gate247inter3));
  inv1  gate985(.a(s_63), .O(gate247inter4));
  nand2 gate986(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate987(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate988(.a(G251), .O(gate247inter7));
  inv1  gate989(.a(G739), .O(gate247inter8));
  nand2 gate990(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate991(.a(s_63), .b(gate247inter3), .O(gate247inter10));
  nor2  gate992(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate993(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate994(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2437(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2438(.a(gate250inter0), .b(s_270), .O(gate250inter1));
  and2  gate2439(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2440(.a(s_270), .O(gate250inter3));
  inv1  gate2441(.a(s_271), .O(gate250inter4));
  nand2 gate2442(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2443(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2444(.a(G706), .O(gate250inter7));
  inv1  gate2445(.a(G742), .O(gate250inter8));
  nand2 gate2446(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2447(.a(s_271), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2448(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2449(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2450(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1051(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1052(.a(gate256inter0), .b(s_72), .O(gate256inter1));
  and2  gate1053(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1054(.a(s_72), .O(gate256inter3));
  inv1  gate1055(.a(s_73), .O(gate256inter4));
  nand2 gate1056(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1057(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1058(.a(G715), .O(gate256inter7));
  inv1  gate1059(.a(G751), .O(gate256inter8));
  nand2 gate1060(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1061(.a(s_73), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1062(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1063(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1064(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate2283(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2284(.a(gate259inter0), .b(s_248), .O(gate259inter1));
  and2  gate2285(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2286(.a(s_248), .O(gate259inter3));
  inv1  gate2287(.a(s_249), .O(gate259inter4));
  nand2 gate2288(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2289(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2290(.a(G758), .O(gate259inter7));
  inv1  gate2291(.a(G759), .O(gate259inter8));
  nand2 gate2292(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2293(.a(s_249), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2294(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2295(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2296(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1037(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1038(.a(gate261inter0), .b(s_70), .O(gate261inter1));
  and2  gate1039(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1040(.a(s_70), .O(gate261inter3));
  inv1  gate1041(.a(s_71), .O(gate261inter4));
  nand2 gate1042(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1043(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1044(.a(G762), .O(gate261inter7));
  inv1  gate1045(.a(G763), .O(gate261inter8));
  nand2 gate1046(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1047(.a(s_71), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1048(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1049(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1050(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1009(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1010(.a(gate262inter0), .b(s_66), .O(gate262inter1));
  and2  gate1011(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1012(.a(s_66), .O(gate262inter3));
  inv1  gate1013(.a(s_67), .O(gate262inter4));
  nand2 gate1014(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1015(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1016(.a(G764), .O(gate262inter7));
  inv1  gate1017(.a(G765), .O(gate262inter8));
  nand2 gate1018(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1019(.a(s_67), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1020(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1021(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1022(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1513(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1514(.a(gate264inter0), .b(s_138), .O(gate264inter1));
  and2  gate1515(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1516(.a(s_138), .O(gate264inter3));
  inv1  gate1517(.a(s_139), .O(gate264inter4));
  nand2 gate1518(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1519(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1520(.a(G768), .O(gate264inter7));
  inv1  gate1521(.a(G769), .O(gate264inter8));
  nand2 gate1522(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1523(.a(s_139), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1524(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1525(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1526(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate673(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate674(.a(gate266inter0), .b(s_18), .O(gate266inter1));
  and2  gate675(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate676(.a(s_18), .O(gate266inter3));
  inv1  gate677(.a(s_19), .O(gate266inter4));
  nand2 gate678(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate679(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate680(.a(G645), .O(gate266inter7));
  inv1  gate681(.a(G773), .O(gate266inter8));
  nand2 gate682(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate683(.a(s_19), .b(gate266inter3), .O(gate266inter10));
  nor2  gate684(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate685(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate686(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2115(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2116(.a(gate269inter0), .b(s_224), .O(gate269inter1));
  and2  gate2117(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2118(.a(s_224), .O(gate269inter3));
  inv1  gate2119(.a(s_225), .O(gate269inter4));
  nand2 gate2120(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2121(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2122(.a(G654), .O(gate269inter7));
  inv1  gate2123(.a(G782), .O(gate269inter8));
  nand2 gate2124(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2125(.a(s_225), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2126(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2127(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2128(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2661(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2662(.a(gate271inter0), .b(s_302), .O(gate271inter1));
  and2  gate2663(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2664(.a(s_302), .O(gate271inter3));
  inv1  gate2665(.a(s_303), .O(gate271inter4));
  nand2 gate2666(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2667(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2668(.a(G660), .O(gate271inter7));
  inv1  gate2669(.a(G788), .O(gate271inter8));
  nand2 gate2670(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2671(.a(s_303), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2672(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2673(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2674(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2773(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2774(.a(gate273inter0), .b(s_318), .O(gate273inter1));
  and2  gate2775(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2776(.a(s_318), .O(gate273inter3));
  inv1  gate2777(.a(s_319), .O(gate273inter4));
  nand2 gate2778(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2779(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2780(.a(G642), .O(gate273inter7));
  inv1  gate2781(.a(G794), .O(gate273inter8));
  nand2 gate2782(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2783(.a(s_319), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2784(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2785(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2786(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2213(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2214(.a(gate274inter0), .b(s_238), .O(gate274inter1));
  and2  gate2215(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2216(.a(s_238), .O(gate274inter3));
  inv1  gate2217(.a(s_239), .O(gate274inter4));
  nand2 gate2218(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2219(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2220(.a(G770), .O(gate274inter7));
  inv1  gate2221(.a(G794), .O(gate274inter8));
  nand2 gate2222(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2223(.a(s_239), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2224(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2225(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2226(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1877(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1878(.a(gate275inter0), .b(s_190), .O(gate275inter1));
  and2  gate1879(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1880(.a(s_190), .O(gate275inter3));
  inv1  gate1881(.a(s_191), .O(gate275inter4));
  nand2 gate1882(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1883(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1884(.a(G645), .O(gate275inter7));
  inv1  gate1885(.a(G797), .O(gate275inter8));
  nand2 gate1886(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1887(.a(s_191), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1888(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1889(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1890(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate645(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate646(.a(gate276inter0), .b(s_14), .O(gate276inter1));
  and2  gate647(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate648(.a(s_14), .O(gate276inter3));
  inv1  gate649(.a(s_15), .O(gate276inter4));
  nand2 gate650(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate651(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate652(.a(G773), .O(gate276inter7));
  inv1  gate653(.a(G797), .O(gate276inter8));
  nand2 gate654(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate655(.a(s_15), .b(gate276inter3), .O(gate276inter10));
  nor2  gate656(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate657(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate658(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2521(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2522(.a(gate279inter0), .b(s_282), .O(gate279inter1));
  and2  gate2523(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2524(.a(s_282), .O(gate279inter3));
  inv1  gate2525(.a(s_283), .O(gate279inter4));
  nand2 gate2526(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2527(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2528(.a(G651), .O(gate279inter7));
  inv1  gate2529(.a(G803), .O(gate279inter8));
  nand2 gate2530(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2531(.a(s_283), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2532(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2533(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2534(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1023(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1024(.a(gate283inter0), .b(s_68), .O(gate283inter1));
  and2  gate1025(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1026(.a(s_68), .O(gate283inter3));
  inv1  gate1027(.a(s_69), .O(gate283inter4));
  nand2 gate1028(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1029(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1030(.a(G657), .O(gate283inter7));
  inv1  gate1031(.a(G809), .O(gate283inter8));
  nand2 gate1032(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1033(.a(s_69), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1034(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1035(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1036(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1709(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1710(.a(gate284inter0), .b(s_166), .O(gate284inter1));
  and2  gate1711(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1712(.a(s_166), .O(gate284inter3));
  inv1  gate1713(.a(s_167), .O(gate284inter4));
  nand2 gate1714(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1715(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1716(.a(G785), .O(gate284inter7));
  inv1  gate1717(.a(G809), .O(gate284inter8));
  nand2 gate1718(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1719(.a(s_167), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1720(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1721(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1722(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1247(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1248(.a(gate285inter0), .b(s_100), .O(gate285inter1));
  and2  gate1249(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1250(.a(s_100), .O(gate285inter3));
  inv1  gate1251(.a(s_101), .O(gate285inter4));
  nand2 gate1252(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1253(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1254(.a(G660), .O(gate285inter7));
  inv1  gate1255(.a(G812), .O(gate285inter8));
  nand2 gate1256(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1257(.a(s_101), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1258(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1259(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1260(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1373(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1374(.a(gate288inter0), .b(s_118), .O(gate288inter1));
  and2  gate1375(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1376(.a(s_118), .O(gate288inter3));
  inv1  gate1377(.a(s_119), .O(gate288inter4));
  nand2 gate1378(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1379(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1380(.a(G791), .O(gate288inter7));
  inv1  gate1381(.a(G815), .O(gate288inter8));
  nand2 gate1382(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1383(.a(s_119), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1384(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1385(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1386(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2927(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2928(.a(gate290inter0), .b(s_340), .O(gate290inter1));
  and2  gate2929(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2930(.a(s_340), .O(gate290inter3));
  inv1  gate2931(.a(s_341), .O(gate290inter4));
  nand2 gate2932(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2933(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2934(.a(G820), .O(gate290inter7));
  inv1  gate2935(.a(G821), .O(gate290inter8));
  nand2 gate2936(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2937(.a(s_341), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2938(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2939(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2940(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1541(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1542(.a(gate291inter0), .b(s_142), .O(gate291inter1));
  and2  gate1543(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1544(.a(s_142), .O(gate291inter3));
  inv1  gate1545(.a(s_143), .O(gate291inter4));
  nand2 gate1546(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1547(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1548(.a(G822), .O(gate291inter7));
  inv1  gate1549(.a(G823), .O(gate291inter8));
  nand2 gate1550(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1551(.a(s_143), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1552(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1553(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1554(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate2689(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2690(.a(gate292inter0), .b(s_306), .O(gate292inter1));
  and2  gate2691(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2692(.a(s_306), .O(gate292inter3));
  inv1  gate2693(.a(s_307), .O(gate292inter4));
  nand2 gate2694(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2695(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2696(.a(G824), .O(gate292inter7));
  inv1  gate2697(.a(G825), .O(gate292inter8));
  nand2 gate2698(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2699(.a(s_307), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2700(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2701(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2702(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1107(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1108(.a(gate295inter0), .b(s_80), .O(gate295inter1));
  and2  gate1109(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1110(.a(s_80), .O(gate295inter3));
  inv1  gate1111(.a(s_81), .O(gate295inter4));
  nand2 gate1112(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1113(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1114(.a(G830), .O(gate295inter7));
  inv1  gate1115(.a(G831), .O(gate295inter8));
  nand2 gate1116(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1117(.a(s_81), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1118(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1119(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1120(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1975(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1976(.a(gate296inter0), .b(s_204), .O(gate296inter1));
  and2  gate1977(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1978(.a(s_204), .O(gate296inter3));
  inv1  gate1979(.a(s_205), .O(gate296inter4));
  nand2 gate1980(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1981(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1982(.a(G826), .O(gate296inter7));
  inv1  gate1983(.a(G827), .O(gate296inter8));
  nand2 gate1984(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1985(.a(s_205), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1986(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1987(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1988(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1681(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1682(.a(gate388inter0), .b(s_162), .O(gate388inter1));
  and2  gate1683(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1684(.a(s_162), .O(gate388inter3));
  inv1  gate1685(.a(s_163), .O(gate388inter4));
  nand2 gate1686(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1687(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1688(.a(G2), .O(gate388inter7));
  inv1  gate1689(.a(G1039), .O(gate388inter8));
  nand2 gate1690(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1691(.a(s_163), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1692(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1693(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1694(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate687(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate688(.a(gate394inter0), .b(s_20), .O(gate394inter1));
  and2  gate689(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate690(.a(s_20), .O(gate394inter3));
  inv1  gate691(.a(s_21), .O(gate394inter4));
  nand2 gate692(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate693(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate694(.a(G8), .O(gate394inter7));
  inv1  gate695(.a(G1057), .O(gate394inter8));
  nand2 gate696(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate697(.a(s_21), .b(gate394inter3), .O(gate394inter10));
  nor2  gate698(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate699(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate700(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2619(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2620(.a(gate396inter0), .b(s_296), .O(gate396inter1));
  and2  gate2621(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2622(.a(s_296), .O(gate396inter3));
  inv1  gate2623(.a(s_297), .O(gate396inter4));
  nand2 gate2624(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2625(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2626(.a(G10), .O(gate396inter7));
  inv1  gate2627(.a(G1063), .O(gate396inter8));
  nand2 gate2628(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2629(.a(s_297), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2630(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2631(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2632(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1947(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1948(.a(gate398inter0), .b(s_200), .O(gate398inter1));
  and2  gate1949(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1950(.a(s_200), .O(gate398inter3));
  inv1  gate1951(.a(s_201), .O(gate398inter4));
  nand2 gate1952(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1953(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1954(.a(G12), .O(gate398inter7));
  inv1  gate1955(.a(G1069), .O(gate398inter8));
  nand2 gate1956(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1957(.a(s_201), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1958(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1959(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1960(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1289(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1290(.a(gate399inter0), .b(s_106), .O(gate399inter1));
  and2  gate1291(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1292(.a(s_106), .O(gate399inter3));
  inv1  gate1293(.a(s_107), .O(gate399inter4));
  nand2 gate1294(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1295(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1296(.a(G13), .O(gate399inter7));
  inv1  gate1297(.a(G1072), .O(gate399inter8));
  nand2 gate1298(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1299(.a(s_107), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1300(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1301(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1302(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1415(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1416(.a(gate400inter0), .b(s_124), .O(gate400inter1));
  and2  gate1417(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1418(.a(s_124), .O(gate400inter3));
  inv1  gate1419(.a(s_125), .O(gate400inter4));
  nand2 gate1420(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1421(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1422(.a(G14), .O(gate400inter7));
  inv1  gate1423(.a(G1075), .O(gate400inter8));
  nand2 gate1424(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1425(.a(s_125), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1426(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1427(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1428(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2325(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2326(.a(gate401inter0), .b(s_254), .O(gate401inter1));
  and2  gate2327(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2328(.a(s_254), .O(gate401inter3));
  inv1  gate2329(.a(s_255), .O(gate401inter4));
  nand2 gate2330(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2331(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2332(.a(G15), .O(gate401inter7));
  inv1  gate2333(.a(G1078), .O(gate401inter8));
  nand2 gate2334(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2335(.a(s_255), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2336(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2337(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2338(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate2073(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2074(.a(gate402inter0), .b(s_218), .O(gate402inter1));
  and2  gate2075(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2076(.a(s_218), .O(gate402inter3));
  inv1  gate2077(.a(s_219), .O(gate402inter4));
  nand2 gate2078(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2079(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2080(.a(G16), .O(gate402inter7));
  inv1  gate2081(.a(G1081), .O(gate402inter8));
  nand2 gate2082(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2083(.a(s_219), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2084(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2085(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2086(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1639(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1640(.a(gate404inter0), .b(s_156), .O(gate404inter1));
  and2  gate1641(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1642(.a(s_156), .O(gate404inter3));
  inv1  gate1643(.a(s_157), .O(gate404inter4));
  nand2 gate1644(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1645(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1646(.a(G18), .O(gate404inter7));
  inv1  gate1647(.a(G1087), .O(gate404inter8));
  nand2 gate1648(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1649(.a(s_157), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1650(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1651(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1652(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1345(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1346(.a(gate406inter0), .b(s_114), .O(gate406inter1));
  and2  gate1347(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1348(.a(s_114), .O(gate406inter3));
  inv1  gate1349(.a(s_115), .O(gate406inter4));
  nand2 gate1350(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1351(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1352(.a(G20), .O(gate406inter7));
  inv1  gate1353(.a(G1093), .O(gate406inter8));
  nand2 gate1354(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1355(.a(s_115), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1356(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1357(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1358(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1667(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1668(.a(gate407inter0), .b(s_160), .O(gate407inter1));
  and2  gate1669(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1670(.a(s_160), .O(gate407inter3));
  inv1  gate1671(.a(s_161), .O(gate407inter4));
  nand2 gate1672(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1673(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1674(.a(G21), .O(gate407inter7));
  inv1  gate1675(.a(G1096), .O(gate407inter8));
  nand2 gate1676(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1677(.a(s_161), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1678(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1679(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1680(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1919(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1920(.a(gate409inter0), .b(s_196), .O(gate409inter1));
  and2  gate1921(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1922(.a(s_196), .O(gate409inter3));
  inv1  gate1923(.a(s_197), .O(gate409inter4));
  nand2 gate1924(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1925(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1926(.a(G23), .O(gate409inter7));
  inv1  gate1927(.a(G1102), .O(gate409inter8));
  nand2 gate1928(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1929(.a(s_197), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1930(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1931(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1932(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2913(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2914(.a(gate410inter0), .b(s_338), .O(gate410inter1));
  and2  gate2915(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2916(.a(s_338), .O(gate410inter3));
  inv1  gate2917(.a(s_339), .O(gate410inter4));
  nand2 gate2918(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2919(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2920(.a(G24), .O(gate410inter7));
  inv1  gate2921(.a(G1105), .O(gate410inter8));
  nand2 gate2922(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2923(.a(s_339), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2924(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2925(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2926(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2493(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2494(.a(gate413inter0), .b(s_278), .O(gate413inter1));
  and2  gate2495(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2496(.a(s_278), .O(gate413inter3));
  inv1  gate2497(.a(s_279), .O(gate413inter4));
  nand2 gate2498(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2499(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2500(.a(G27), .O(gate413inter7));
  inv1  gate2501(.a(G1114), .O(gate413inter8));
  nand2 gate2502(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2503(.a(s_279), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2504(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2505(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2506(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1765(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1766(.a(gate414inter0), .b(s_174), .O(gate414inter1));
  and2  gate1767(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1768(.a(s_174), .O(gate414inter3));
  inv1  gate1769(.a(s_175), .O(gate414inter4));
  nand2 gate1770(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1771(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1772(.a(G28), .O(gate414inter7));
  inv1  gate1773(.a(G1117), .O(gate414inter8));
  nand2 gate1774(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1775(.a(s_175), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1776(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1777(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1778(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2311(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2312(.a(gate416inter0), .b(s_252), .O(gate416inter1));
  and2  gate2313(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2314(.a(s_252), .O(gate416inter3));
  inv1  gate2315(.a(s_253), .O(gate416inter4));
  nand2 gate2316(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2317(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2318(.a(G30), .O(gate416inter7));
  inv1  gate2319(.a(G1123), .O(gate416inter8));
  nand2 gate2320(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2321(.a(s_253), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2322(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2323(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2324(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1905(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1906(.a(gate418inter0), .b(s_194), .O(gate418inter1));
  and2  gate1907(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1908(.a(s_194), .O(gate418inter3));
  inv1  gate1909(.a(s_195), .O(gate418inter4));
  nand2 gate1910(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1911(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1912(.a(G32), .O(gate418inter7));
  inv1  gate1913(.a(G1129), .O(gate418inter8));
  nand2 gate1914(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1915(.a(s_195), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1916(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1917(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1918(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1135(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1136(.a(gate419inter0), .b(s_84), .O(gate419inter1));
  and2  gate1137(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1138(.a(s_84), .O(gate419inter3));
  inv1  gate1139(.a(s_85), .O(gate419inter4));
  nand2 gate1140(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1141(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1142(.a(G1), .O(gate419inter7));
  inv1  gate1143(.a(G1132), .O(gate419inter8));
  nand2 gate1144(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1145(.a(s_85), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1146(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1147(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1148(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2171(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2172(.a(gate426inter0), .b(s_232), .O(gate426inter1));
  and2  gate2173(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2174(.a(s_232), .O(gate426inter3));
  inv1  gate2175(.a(s_233), .O(gate426inter4));
  nand2 gate2176(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2177(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2178(.a(G1045), .O(gate426inter7));
  inv1  gate2179(.a(G1141), .O(gate426inter8));
  nand2 gate2180(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2181(.a(s_233), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2182(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2183(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2184(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2899(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2900(.a(gate430inter0), .b(s_336), .O(gate430inter1));
  and2  gate2901(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2902(.a(s_336), .O(gate430inter3));
  inv1  gate2903(.a(s_337), .O(gate430inter4));
  nand2 gate2904(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2905(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2906(.a(G1051), .O(gate430inter7));
  inv1  gate2907(.a(G1147), .O(gate430inter8));
  nand2 gate2908(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2909(.a(s_337), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2910(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2911(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2912(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2451(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2452(.a(gate432inter0), .b(s_272), .O(gate432inter1));
  and2  gate2453(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2454(.a(s_272), .O(gate432inter3));
  inv1  gate2455(.a(s_273), .O(gate432inter4));
  nand2 gate2456(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2457(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2458(.a(G1054), .O(gate432inter7));
  inv1  gate2459(.a(G1150), .O(gate432inter8));
  nand2 gate2460(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2461(.a(s_273), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2462(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2463(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2464(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1989(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1990(.a(gate434inter0), .b(s_206), .O(gate434inter1));
  and2  gate1991(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1992(.a(s_206), .O(gate434inter3));
  inv1  gate1993(.a(s_207), .O(gate434inter4));
  nand2 gate1994(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1995(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1996(.a(G1057), .O(gate434inter7));
  inv1  gate1997(.a(G1153), .O(gate434inter8));
  nand2 gate1998(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1999(.a(s_207), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2000(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2001(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2002(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate2829(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2830(.a(gate437inter0), .b(s_326), .O(gate437inter1));
  and2  gate2831(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2832(.a(s_326), .O(gate437inter3));
  inv1  gate2833(.a(s_327), .O(gate437inter4));
  nand2 gate2834(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2835(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2836(.a(G10), .O(gate437inter7));
  inv1  gate2837(.a(G1159), .O(gate437inter8));
  nand2 gate2838(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2839(.a(s_327), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2840(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2841(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2842(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2731(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2732(.a(gate439inter0), .b(s_312), .O(gate439inter1));
  and2  gate2733(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2734(.a(s_312), .O(gate439inter3));
  inv1  gate2735(.a(s_313), .O(gate439inter4));
  nand2 gate2736(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2737(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2738(.a(G11), .O(gate439inter7));
  inv1  gate2739(.a(G1162), .O(gate439inter8));
  nand2 gate2740(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2741(.a(s_313), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2742(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2743(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2744(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1625(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1626(.a(gate440inter0), .b(s_154), .O(gate440inter1));
  and2  gate1627(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1628(.a(s_154), .O(gate440inter3));
  inv1  gate1629(.a(s_155), .O(gate440inter4));
  nand2 gate1630(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1631(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1632(.a(G1066), .O(gate440inter7));
  inv1  gate1633(.a(G1162), .O(gate440inter8));
  nand2 gate1634(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1635(.a(s_155), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1636(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1637(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1638(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate715(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate716(.a(gate442inter0), .b(s_24), .O(gate442inter1));
  and2  gate717(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate718(.a(s_24), .O(gate442inter3));
  inv1  gate719(.a(s_25), .O(gate442inter4));
  nand2 gate720(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate721(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate722(.a(G1069), .O(gate442inter7));
  inv1  gate723(.a(G1165), .O(gate442inter8));
  nand2 gate724(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate725(.a(s_25), .b(gate442inter3), .O(gate442inter10));
  nor2  gate726(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate727(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate728(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2941(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2942(.a(gate444inter0), .b(s_342), .O(gate444inter1));
  and2  gate2943(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2944(.a(s_342), .O(gate444inter3));
  inv1  gate2945(.a(s_343), .O(gate444inter4));
  nand2 gate2946(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2947(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2948(.a(G1072), .O(gate444inter7));
  inv1  gate2949(.a(G1168), .O(gate444inter8));
  nand2 gate2950(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2951(.a(s_343), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2952(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2953(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2954(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate827(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate828(.a(gate450inter0), .b(s_40), .O(gate450inter1));
  and2  gate829(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate830(.a(s_40), .O(gate450inter3));
  inv1  gate831(.a(s_41), .O(gate450inter4));
  nand2 gate832(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate833(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate834(.a(G1081), .O(gate450inter7));
  inv1  gate835(.a(G1177), .O(gate450inter8));
  nand2 gate836(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate837(.a(s_41), .b(gate450inter3), .O(gate450inter10));
  nor2  gate838(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate839(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate840(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2983(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2984(.a(gate452inter0), .b(s_348), .O(gate452inter1));
  and2  gate2985(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2986(.a(s_348), .O(gate452inter3));
  inv1  gate2987(.a(s_349), .O(gate452inter4));
  nand2 gate2988(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2989(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2990(.a(G1084), .O(gate452inter7));
  inv1  gate2991(.a(G1180), .O(gate452inter8));
  nand2 gate2992(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2993(.a(s_349), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2994(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2995(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2996(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate617(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate618(.a(gate453inter0), .b(s_10), .O(gate453inter1));
  and2  gate619(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate620(.a(s_10), .O(gate453inter3));
  inv1  gate621(.a(s_11), .O(gate453inter4));
  nand2 gate622(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate623(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate624(.a(G18), .O(gate453inter7));
  inv1  gate625(.a(G1183), .O(gate453inter8));
  nand2 gate626(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate627(.a(s_11), .b(gate453inter3), .O(gate453inter10));
  nor2  gate628(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate629(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate630(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1079(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1080(.a(gate454inter0), .b(s_76), .O(gate454inter1));
  and2  gate1081(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1082(.a(s_76), .O(gate454inter3));
  inv1  gate1083(.a(s_77), .O(gate454inter4));
  nand2 gate1084(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1085(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1086(.a(G1087), .O(gate454inter7));
  inv1  gate1087(.a(G1183), .O(gate454inter8));
  nand2 gate1088(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1089(.a(s_77), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1090(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1091(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1092(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1751(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1752(.a(gate458inter0), .b(s_172), .O(gate458inter1));
  and2  gate1753(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1754(.a(s_172), .O(gate458inter3));
  inv1  gate1755(.a(s_173), .O(gate458inter4));
  nand2 gate1756(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1757(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1758(.a(G1093), .O(gate458inter7));
  inv1  gate1759(.a(G1189), .O(gate458inter8));
  nand2 gate1760(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1761(.a(s_173), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1762(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1763(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1764(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2801(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2802(.a(gate462inter0), .b(s_322), .O(gate462inter1));
  and2  gate2803(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2804(.a(s_322), .O(gate462inter3));
  inv1  gate2805(.a(s_323), .O(gate462inter4));
  nand2 gate2806(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2807(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2808(.a(G1099), .O(gate462inter7));
  inv1  gate2809(.a(G1195), .O(gate462inter8));
  nand2 gate2810(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2811(.a(s_323), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2812(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2813(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2814(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2563(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2564(.a(gate466inter0), .b(s_288), .O(gate466inter1));
  and2  gate2565(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2566(.a(s_288), .O(gate466inter3));
  inv1  gate2567(.a(s_289), .O(gate466inter4));
  nand2 gate2568(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2569(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2570(.a(G1105), .O(gate466inter7));
  inv1  gate2571(.a(G1201), .O(gate466inter8));
  nand2 gate2572(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2573(.a(s_289), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2574(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2575(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2576(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate575(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate576(.a(gate467inter0), .b(s_4), .O(gate467inter1));
  and2  gate577(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate578(.a(s_4), .O(gate467inter3));
  inv1  gate579(.a(s_5), .O(gate467inter4));
  nand2 gate580(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate581(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate582(.a(G25), .O(gate467inter7));
  inv1  gate583(.a(G1204), .O(gate467inter8));
  nand2 gate584(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate585(.a(s_5), .b(gate467inter3), .O(gate467inter10));
  nor2  gate586(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate587(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate588(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2241(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2242(.a(gate470inter0), .b(s_242), .O(gate470inter1));
  and2  gate2243(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2244(.a(s_242), .O(gate470inter3));
  inv1  gate2245(.a(s_243), .O(gate470inter4));
  nand2 gate2246(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2247(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2248(.a(G1111), .O(gate470inter7));
  inv1  gate2249(.a(G1207), .O(gate470inter8));
  nand2 gate2250(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2251(.a(s_243), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2252(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2253(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2254(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate729(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate730(.a(gate471inter0), .b(s_26), .O(gate471inter1));
  and2  gate731(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate732(.a(s_26), .O(gate471inter3));
  inv1  gate733(.a(s_27), .O(gate471inter4));
  nand2 gate734(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate735(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate736(.a(G27), .O(gate471inter7));
  inv1  gate737(.a(G1210), .O(gate471inter8));
  nand2 gate738(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate739(.a(s_27), .b(gate471inter3), .O(gate471inter10));
  nor2  gate740(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate741(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate742(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1233(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1234(.a(gate476inter0), .b(s_98), .O(gate476inter1));
  and2  gate1235(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1236(.a(s_98), .O(gate476inter3));
  inv1  gate1237(.a(s_99), .O(gate476inter4));
  nand2 gate1238(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1239(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1240(.a(G1120), .O(gate476inter7));
  inv1  gate1241(.a(G1216), .O(gate476inter8));
  nand2 gate1242(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1243(.a(s_99), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1244(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1245(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1246(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2423(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2424(.a(gate478inter0), .b(s_268), .O(gate478inter1));
  and2  gate2425(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2426(.a(s_268), .O(gate478inter3));
  inv1  gate2427(.a(s_269), .O(gate478inter4));
  nand2 gate2428(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2429(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2430(.a(G1123), .O(gate478inter7));
  inv1  gate2431(.a(G1219), .O(gate478inter8));
  nand2 gate2432(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2433(.a(s_269), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2434(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2435(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2436(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2339(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2340(.a(gate480inter0), .b(s_256), .O(gate480inter1));
  and2  gate2341(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2342(.a(s_256), .O(gate480inter3));
  inv1  gate2343(.a(s_257), .O(gate480inter4));
  nand2 gate2344(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2345(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2346(.a(G1126), .O(gate480inter7));
  inv1  gate2347(.a(G1222), .O(gate480inter8));
  nand2 gate2348(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2349(.a(s_257), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2350(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2351(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2352(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1443(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1444(.a(gate482inter0), .b(s_128), .O(gate482inter1));
  and2  gate1445(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1446(.a(s_128), .O(gate482inter3));
  inv1  gate1447(.a(s_129), .O(gate482inter4));
  nand2 gate1448(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1449(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1450(.a(G1129), .O(gate482inter7));
  inv1  gate1451(.a(G1225), .O(gate482inter8));
  nand2 gate1452(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1453(.a(s_129), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1454(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1455(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1456(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1653(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1654(.a(gate483inter0), .b(s_158), .O(gate483inter1));
  and2  gate1655(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1656(.a(s_158), .O(gate483inter3));
  inv1  gate1657(.a(s_159), .O(gate483inter4));
  nand2 gate1658(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1659(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1660(.a(G1228), .O(gate483inter7));
  inv1  gate1661(.a(G1229), .O(gate483inter8));
  nand2 gate1662(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1663(.a(s_159), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1664(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1665(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1666(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2367(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2368(.a(gate485inter0), .b(s_260), .O(gate485inter1));
  and2  gate2369(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2370(.a(s_260), .O(gate485inter3));
  inv1  gate2371(.a(s_261), .O(gate485inter4));
  nand2 gate2372(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2373(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2374(.a(G1232), .O(gate485inter7));
  inv1  gate2375(.a(G1233), .O(gate485inter8));
  nand2 gate2376(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2377(.a(s_261), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2378(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2379(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2380(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2017(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2018(.a(gate489inter0), .b(s_210), .O(gate489inter1));
  and2  gate2019(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2020(.a(s_210), .O(gate489inter3));
  inv1  gate2021(.a(s_211), .O(gate489inter4));
  nand2 gate2022(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2023(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2024(.a(G1240), .O(gate489inter7));
  inv1  gate2025(.a(G1241), .O(gate489inter8));
  nand2 gate2026(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2027(.a(s_211), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2028(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2029(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2030(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2143(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2144(.a(gate491inter0), .b(s_228), .O(gate491inter1));
  and2  gate2145(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2146(.a(s_228), .O(gate491inter3));
  inv1  gate2147(.a(s_229), .O(gate491inter4));
  nand2 gate2148(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2149(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2150(.a(G1244), .O(gate491inter7));
  inv1  gate2151(.a(G1245), .O(gate491inter8));
  nand2 gate2152(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2153(.a(s_229), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2154(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2155(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2156(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1933(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1934(.a(gate494inter0), .b(s_198), .O(gate494inter1));
  and2  gate1935(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1936(.a(s_198), .O(gate494inter3));
  inv1  gate1937(.a(s_199), .O(gate494inter4));
  nand2 gate1938(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1939(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1940(.a(G1250), .O(gate494inter7));
  inv1  gate1941(.a(G1251), .O(gate494inter8));
  nand2 gate1942(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1943(.a(s_199), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1944(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1945(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1946(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1695(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1696(.a(gate496inter0), .b(s_164), .O(gate496inter1));
  and2  gate1697(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1698(.a(s_164), .O(gate496inter3));
  inv1  gate1699(.a(s_165), .O(gate496inter4));
  nand2 gate1700(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1701(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1702(.a(G1254), .O(gate496inter7));
  inv1  gate1703(.a(G1255), .O(gate496inter8));
  nand2 gate1704(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1705(.a(s_165), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1706(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1707(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1708(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate701(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate702(.a(gate497inter0), .b(s_22), .O(gate497inter1));
  and2  gate703(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate704(.a(s_22), .O(gate497inter3));
  inv1  gate705(.a(s_23), .O(gate497inter4));
  nand2 gate706(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate707(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate708(.a(G1256), .O(gate497inter7));
  inv1  gate709(.a(G1257), .O(gate497inter8));
  nand2 gate710(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate711(.a(s_23), .b(gate497inter3), .O(gate497inter10));
  nor2  gate712(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate713(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate714(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2185(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2186(.a(gate499inter0), .b(s_234), .O(gate499inter1));
  and2  gate2187(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2188(.a(s_234), .O(gate499inter3));
  inv1  gate2189(.a(s_235), .O(gate499inter4));
  nand2 gate2190(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2191(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2192(.a(G1260), .O(gate499inter7));
  inv1  gate2193(.a(G1261), .O(gate499inter8));
  nand2 gate2194(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2195(.a(s_235), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2196(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2197(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2198(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1401(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1402(.a(gate500inter0), .b(s_122), .O(gate500inter1));
  and2  gate1403(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1404(.a(s_122), .O(gate500inter3));
  inv1  gate1405(.a(s_123), .O(gate500inter4));
  nand2 gate1406(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1407(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1408(.a(G1262), .O(gate500inter7));
  inv1  gate1409(.a(G1263), .O(gate500inter8));
  nand2 gate1410(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1411(.a(s_123), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1412(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1413(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1414(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2353(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2354(.a(gate501inter0), .b(s_258), .O(gate501inter1));
  and2  gate2355(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2356(.a(s_258), .O(gate501inter3));
  inv1  gate2357(.a(s_259), .O(gate501inter4));
  nand2 gate2358(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2359(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2360(.a(G1264), .O(gate501inter7));
  inv1  gate2361(.a(G1265), .O(gate501inter8));
  nand2 gate2362(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2363(.a(s_259), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2364(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2365(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2366(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate967(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate968(.a(gate502inter0), .b(s_60), .O(gate502inter1));
  and2  gate969(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate970(.a(s_60), .O(gate502inter3));
  inv1  gate971(.a(s_61), .O(gate502inter4));
  nand2 gate972(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate973(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate974(.a(G1266), .O(gate502inter7));
  inv1  gate975(.a(G1267), .O(gate502inter8));
  nand2 gate976(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate977(.a(s_61), .b(gate502inter3), .O(gate502inter10));
  nor2  gate978(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate979(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate980(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1275(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1276(.a(gate504inter0), .b(s_104), .O(gate504inter1));
  and2  gate1277(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1278(.a(s_104), .O(gate504inter3));
  inv1  gate1279(.a(s_105), .O(gate504inter4));
  nand2 gate1280(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1281(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1282(.a(G1270), .O(gate504inter7));
  inv1  gate1283(.a(G1271), .O(gate504inter8));
  nand2 gate1284(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1285(.a(s_105), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1286(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1287(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1288(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2591(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2592(.a(gate508inter0), .b(s_292), .O(gate508inter1));
  and2  gate2593(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2594(.a(s_292), .O(gate508inter3));
  inv1  gate2595(.a(s_293), .O(gate508inter4));
  nand2 gate2596(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2597(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2598(.a(G1278), .O(gate508inter7));
  inv1  gate2599(.a(G1279), .O(gate508inter8));
  nand2 gate2600(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2601(.a(s_293), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2602(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2603(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2604(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1611(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1612(.a(gate509inter0), .b(s_152), .O(gate509inter1));
  and2  gate1613(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1614(.a(s_152), .O(gate509inter3));
  inv1  gate1615(.a(s_153), .O(gate509inter4));
  nand2 gate1616(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1617(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1618(.a(G1280), .O(gate509inter7));
  inv1  gate1619(.a(G1281), .O(gate509inter8));
  nand2 gate1620(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1621(.a(s_153), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1622(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1623(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1624(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule