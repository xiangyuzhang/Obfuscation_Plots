module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2577(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2578(.a(gate11inter0), .b(s_290), .O(gate11inter1));
  and2  gate2579(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2580(.a(s_290), .O(gate11inter3));
  inv1  gate2581(.a(s_291), .O(gate11inter4));
  nand2 gate2582(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2583(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2584(.a(G5), .O(gate11inter7));
  inv1  gate2585(.a(G6), .O(gate11inter8));
  nand2 gate2586(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2587(.a(s_291), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2588(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2589(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2590(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1569(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1570(.a(gate13inter0), .b(s_146), .O(gate13inter1));
  and2  gate1571(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1572(.a(s_146), .O(gate13inter3));
  inv1  gate1573(.a(s_147), .O(gate13inter4));
  nand2 gate1574(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1575(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1576(.a(G9), .O(gate13inter7));
  inv1  gate1577(.a(G10), .O(gate13inter8));
  nand2 gate1578(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1579(.a(s_147), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1580(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1581(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1582(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1457(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1458(.a(gate16inter0), .b(s_130), .O(gate16inter1));
  and2  gate1459(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1460(.a(s_130), .O(gate16inter3));
  inv1  gate1461(.a(s_131), .O(gate16inter4));
  nand2 gate1462(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1463(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1464(.a(G15), .O(gate16inter7));
  inv1  gate1465(.a(G16), .O(gate16inter8));
  nand2 gate1466(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1467(.a(s_131), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1468(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1469(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1470(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1611(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1612(.a(gate20inter0), .b(s_152), .O(gate20inter1));
  and2  gate1613(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1614(.a(s_152), .O(gate20inter3));
  inv1  gate1615(.a(s_153), .O(gate20inter4));
  nand2 gate1616(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1617(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1618(.a(G23), .O(gate20inter7));
  inv1  gate1619(.a(G24), .O(gate20inter8));
  nand2 gate1620(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1621(.a(s_153), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1622(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1623(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1624(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2591(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2592(.a(gate22inter0), .b(s_292), .O(gate22inter1));
  and2  gate2593(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2594(.a(s_292), .O(gate22inter3));
  inv1  gate2595(.a(s_293), .O(gate22inter4));
  nand2 gate2596(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2597(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2598(.a(G27), .O(gate22inter7));
  inv1  gate2599(.a(G28), .O(gate22inter8));
  nand2 gate2600(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2601(.a(s_293), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2602(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2603(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2604(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2745(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2746(.a(gate29inter0), .b(s_314), .O(gate29inter1));
  and2  gate2747(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2748(.a(s_314), .O(gate29inter3));
  inv1  gate2749(.a(s_315), .O(gate29inter4));
  nand2 gate2750(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2751(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2752(.a(G3), .O(gate29inter7));
  inv1  gate2753(.a(G7), .O(gate29inter8));
  nand2 gate2754(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2755(.a(s_315), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2756(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2757(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2758(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2269(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2270(.a(gate32inter0), .b(s_246), .O(gate32inter1));
  and2  gate2271(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2272(.a(s_246), .O(gate32inter3));
  inv1  gate2273(.a(s_247), .O(gate32inter4));
  nand2 gate2274(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2275(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2276(.a(G12), .O(gate32inter7));
  inv1  gate2277(.a(G16), .O(gate32inter8));
  nand2 gate2278(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2279(.a(s_247), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2280(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2281(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2282(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1317(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1318(.a(gate33inter0), .b(s_110), .O(gate33inter1));
  and2  gate1319(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1320(.a(s_110), .O(gate33inter3));
  inv1  gate1321(.a(s_111), .O(gate33inter4));
  nand2 gate1322(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1323(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1324(.a(G17), .O(gate33inter7));
  inv1  gate1325(.a(G21), .O(gate33inter8));
  nand2 gate1326(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1327(.a(s_111), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1328(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1329(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1330(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1639(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1640(.a(gate34inter0), .b(s_156), .O(gate34inter1));
  and2  gate1641(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1642(.a(s_156), .O(gate34inter3));
  inv1  gate1643(.a(s_157), .O(gate34inter4));
  nand2 gate1644(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1645(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1646(.a(G25), .O(gate34inter7));
  inv1  gate1647(.a(G29), .O(gate34inter8));
  nand2 gate1648(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1649(.a(s_157), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1650(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1651(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1652(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2409(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2410(.a(gate36inter0), .b(s_266), .O(gate36inter1));
  and2  gate2411(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2412(.a(s_266), .O(gate36inter3));
  inv1  gate2413(.a(s_267), .O(gate36inter4));
  nand2 gate2414(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2415(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2416(.a(G26), .O(gate36inter7));
  inv1  gate2417(.a(G30), .O(gate36inter8));
  nand2 gate2418(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2419(.a(s_267), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2420(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2421(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2422(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1471(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1472(.a(gate37inter0), .b(s_132), .O(gate37inter1));
  and2  gate1473(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1474(.a(s_132), .O(gate37inter3));
  inv1  gate1475(.a(s_133), .O(gate37inter4));
  nand2 gate1476(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1477(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1478(.a(G19), .O(gate37inter7));
  inv1  gate1479(.a(G23), .O(gate37inter8));
  nand2 gate1480(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1481(.a(s_133), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1482(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1483(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1484(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1079(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1080(.a(gate40inter0), .b(s_76), .O(gate40inter1));
  and2  gate1081(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1082(.a(s_76), .O(gate40inter3));
  inv1  gate1083(.a(s_77), .O(gate40inter4));
  nand2 gate1084(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1085(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1086(.a(G28), .O(gate40inter7));
  inv1  gate1087(.a(G32), .O(gate40inter8));
  nand2 gate1088(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1089(.a(s_77), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1090(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1091(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1092(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2689(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2690(.a(gate41inter0), .b(s_306), .O(gate41inter1));
  and2  gate2691(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2692(.a(s_306), .O(gate41inter3));
  inv1  gate2693(.a(s_307), .O(gate41inter4));
  nand2 gate2694(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2695(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2696(.a(G1), .O(gate41inter7));
  inv1  gate2697(.a(G266), .O(gate41inter8));
  nand2 gate2698(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2699(.a(s_307), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2700(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2701(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2702(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2395(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2396(.a(gate47inter0), .b(s_264), .O(gate47inter1));
  and2  gate2397(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2398(.a(s_264), .O(gate47inter3));
  inv1  gate2399(.a(s_265), .O(gate47inter4));
  nand2 gate2400(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2401(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2402(.a(G7), .O(gate47inter7));
  inv1  gate2403(.a(G275), .O(gate47inter8));
  nand2 gate2404(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2405(.a(s_265), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2406(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2407(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2408(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1443(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1444(.a(gate48inter0), .b(s_128), .O(gate48inter1));
  and2  gate1445(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1446(.a(s_128), .O(gate48inter3));
  inv1  gate1447(.a(s_129), .O(gate48inter4));
  nand2 gate1448(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1449(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1450(.a(G8), .O(gate48inter7));
  inv1  gate1451(.a(G275), .O(gate48inter8));
  nand2 gate1452(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1453(.a(s_129), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1454(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1455(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1456(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2157(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2158(.a(gate49inter0), .b(s_230), .O(gate49inter1));
  and2  gate2159(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2160(.a(s_230), .O(gate49inter3));
  inv1  gate2161(.a(s_231), .O(gate49inter4));
  nand2 gate2162(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2163(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2164(.a(G9), .O(gate49inter7));
  inv1  gate2165(.a(G278), .O(gate49inter8));
  nand2 gate2166(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2167(.a(s_231), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2168(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2169(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2170(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1919(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1920(.a(gate50inter0), .b(s_196), .O(gate50inter1));
  and2  gate1921(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1922(.a(s_196), .O(gate50inter3));
  inv1  gate1923(.a(s_197), .O(gate50inter4));
  nand2 gate1924(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1925(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1926(.a(G10), .O(gate50inter7));
  inv1  gate1927(.a(G278), .O(gate50inter8));
  nand2 gate1928(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1929(.a(s_197), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1930(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1931(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1932(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1051(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1052(.a(gate52inter0), .b(s_72), .O(gate52inter1));
  and2  gate1053(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1054(.a(s_72), .O(gate52inter3));
  inv1  gate1055(.a(s_73), .O(gate52inter4));
  nand2 gate1056(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1057(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1058(.a(G12), .O(gate52inter7));
  inv1  gate1059(.a(G281), .O(gate52inter8));
  nand2 gate1060(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1061(.a(s_73), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1062(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1063(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1064(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1261(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1262(.a(gate58inter0), .b(s_102), .O(gate58inter1));
  and2  gate1263(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1264(.a(s_102), .O(gate58inter3));
  inv1  gate1265(.a(s_103), .O(gate58inter4));
  nand2 gate1266(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1267(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1268(.a(G18), .O(gate58inter7));
  inv1  gate1269(.a(G290), .O(gate58inter8));
  nand2 gate1270(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1271(.a(s_103), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1272(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1273(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1274(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1205(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1206(.a(gate63inter0), .b(s_94), .O(gate63inter1));
  and2  gate1207(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1208(.a(s_94), .O(gate63inter3));
  inv1  gate1209(.a(s_95), .O(gate63inter4));
  nand2 gate1210(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1211(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1212(.a(G23), .O(gate63inter7));
  inv1  gate1213(.a(G299), .O(gate63inter8));
  nand2 gate1214(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1215(.a(s_95), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1216(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1217(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1218(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2521(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2522(.a(gate67inter0), .b(s_282), .O(gate67inter1));
  and2  gate2523(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2524(.a(s_282), .O(gate67inter3));
  inv1  gate2525(.a(s_283), .O(gate67inter4));
  nand2 gate2526(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2527(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2528(.a(G27), .O(gate67inter7));
  inv1  gate2529(.a(G305), .O(gate67inter8));
  nand2 gate2530(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2531(.a(s_283), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2532(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2533(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2534(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate589(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate590(.a(gate69inter0), .b(s_6), .O(gate69inter1));
  and2  gate591(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate592(.a(s_6), .O(gate69inter3));
  inv1  gate593(.a(s_7), .O(gate69inter4));
  nand2 gate594(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate595(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate596(.a(G29), .O(gate69inter7));
  inv1  gate597(.a(G308), .O(gate69inter8));
  nand2 gate598(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate599(.a(s_7), .b(gate69inter3), .O(gate69inter10));
  nor2  gate600(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate601(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate602(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1681(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1682(.a(gate73inter0), .b(s_162), .O(gate73inter1));
  and2  gate1683(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1684(.a(s_162), .O(gate73inter3));
  inv1  gate1685(.a(s_163), .O(gate73inter4));
  nand2 gate1686(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1687(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1688(.a(G1), .O(gate73inter7));
  inv1  gate1689(.a(G314), .O(gate73inter8));
  nand2 gate1690(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1691(.a(s_163), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1692(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1693(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1694(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1933(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1934(.a(gate74inter0), .b(s_198), .O(gate74inter1));
  and2  gate1935(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1936(.a(s_198), .O(gate74inter3));
  inv1  gate1937(.a(s_199), .O(gate74inter4));
  nand2 gate1938(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1939(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1940(.a(G5), .O(gate74inter7));
  inv1  gate1941(.a(G314), .O(gate74inter8));
  nand2 gate1942(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1943(.a(s_199), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1944(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1945(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1946(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2199(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2200(.a(gate77inter0), .b(s_236), .O(gate77inter1));
  and2  gate2201(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2202(.a(s_236), .O(gate77inter3));
  inv1  gate2203(.a(s_237), .O(gate77inter4));
  nand2 gate2204(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2205(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2206(.a(G2), .O(gate77inter7));
  inv1  gate2207(.a(G320), .O(gate77inter8));
  nand2 gate2208(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2209(.a(s_237), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2210(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2211(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2212(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate911(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate912(.a(gate79inter0), .b(s_52), .O(gate79inter1));
  and2  gate913(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate914(.a(s_52), .O(gate79inter3));
  inv1  gate915(.a(s_53), .O(gate79inter4));
  nand2 gate916(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate917(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate918(.a(G10), .O(gate79inter7));
  inv1  gate919(.a(G323), .O(gate79inter8));
  nand2 gate920(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate921(.a(s_53), .b(gate79inter3), .O(gate79inter10));
  nor2  gate922(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate923(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate924(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate2031(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2032(.a(gate80inter0), .b(s_212), .O(gate80inter1));
  and2  gate2033(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2034(.a(s_212), .O(gate80inter3));
  inv1  gate2035(.a(s_213), .O(gate80inter4));
  nand2 gate2036(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2037(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2038(.a(G14), .O(gate80inter7));
  inv1  gate2039(.a(G323), .O(gate80inter8));
  nand2 gate2040(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2041(.a(s_213), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2042(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2043(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2044(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1177(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1178(.a(gate84inter0), .b(s_90), .O(gate84inter1));
  and2  gate1179(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1180(.a(s_90), .O(gate84inter3));
  inv1  gate1181(.a(s_91), .O(gate84inter4));
  nand2 gate1182(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1183(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1184(.a(G15), .O(gate84inter7));
  inv1  gate1185(.a(G329), .O(gate84inter8));
  nand2 gate1186(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1187(.a(s_91), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1188(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1189(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1190(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate659(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate660(.a(gate85inter0), .b(s_16), .O(gate85inter1));
  and2  gate661(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate662(.a(s_16), .O(gate85inter3));
  inv1  gate663(.a(s_17), .O(gate85inter4));
  nand2 gate664(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate665(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate666(.a(G4), .O(gate85inter7));
  inv1  gate667(.a(G332), .O(gate85inter8));
  nand2 gate668(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate669(.a(s_17), .b(gate85inter3), .O(gate85inter10));
  nor2  gate670(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate671(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate672(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate827(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate828(.a(gate86inter0), .b(s_40), .O(gate86inter1));
  and2  gate829(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate830(.a(s_40), .O(gate86inter3));
  inv1  gate831(.a(s_41), .O(gate86inter4));
  nand2 gate832(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate833(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate834(.a(G8), .O(gate86inter7));
  inv1  gate835(.a(G332), .O(gate86inter8));
  nand2 gate836(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate837(.a(s_41), .b(gate86inter3), .O(gate86inter10));
  nor2  gate838(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate839(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate840(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate841(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate842(.a(gate91inter0), .b(s_42), .O(gate91inter1));
  and2  gate843(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate844(.a(s_42), .O(gate91inter3));
  inv1  gate845(.a(s_43), .O(gate91inter4));
  nand2 gate846(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate847(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate848(.a(G25), .O(gate91inter7));
  inv1  gate849(.a(G341), .O(gate91inter8));
  nand2 gate850(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate851(.a(s_43), .b(gate91inter3), .O(gate91inter10));
  nor2  gate852(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate853(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate854(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1135(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1136(.a(gate95inter0), .b(s_84), .O(gate95inter1));
  and2  gate1137(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1138(.a(s_84), .O(gate95inter3));
  inv1  gate1139(.a(s_85), .O(gate95inter4));
  nand2 gate1140(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1141(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1142(.a(G26), .O(gate95inter7));
  inv1  gate1143(.a(G347), .O(gate95inter8));
  nand2 gate1144(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1145(.a(s_85), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1146(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1147(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1148(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2549(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2550(.a(gate99inter0), .b(s_286), .O(gate99inter1));
  and2  gate2551(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2552(.a(s_286), .O(gate99inter3));
  inv1  gate2553(.a(s_287), .O(gate99inter4));
  nand2 gate2554(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2555(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2556(.a(G27), .O(gate99inter7));
  inv1  gate2557(.a(G353), .O(gate99inter8));
  nand2 gate2558(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2559(.a(s_287), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2560(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2561(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2562(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate939(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate940(.a(gate100inter0), .b(s_56), .O(gate100inter1));
  and2  gate941(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate942(.a(s_56), .O(gate100inter3));
  inv1  gate943(.a(s_57), .O(gate100inter4));
  nand2 gate944(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate945(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate946(.a(G31), .O(gate100inter7));
  inv1  gate947(.a(G353), .O(gate100inter8));
  nand2 gate948(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate949(.a(s_57), .b(gate100inter3), .O(gate100inter10));
  nor2  gate950(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate951(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate952(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1555(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1556(.a(gate103inter0), .b(s_144), .O(gate103inter1));
  and2  gate1557(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1558(.a(s_144), .O(gate103inter3));
  inv1  gate1559(.a(s_145), .O(gate103inter4));
  nand2 gate1560(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1561(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1562(.a(G28), .O(gate103inter7));
  inv1  gate1563(.a(G359), .O(gate103inter8));
  nand2 gate1564(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1565(.a(s_145), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1566(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1567(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1568(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate631(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate632(.a(gate104inter0), .b(s_12), .O(gate104inter1));
  and2  gate633(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate634(.a(s_12), .O(gate104inter3));
  inv1  gate635(.a(s_13), .O(gate104inter4));
  nand2 gate636(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate637(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate638(.a(G32), .O(gate104inter7));
  inv1  gate639(.a(G359), .O(gate104inter8));
  nand2 gate640(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate641(.a(s_13), .b(gate104inter3), .O(gate104inter10));
  nor2  gate642(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate643(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate644(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate883(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate884(.a(gate107inter0), .b(s_48), .O(gate107inter1));
  and2  gate885(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate886(.a(s_48), .O(gate107inter3));
  inv1  gate887(.a(s_49), .O(gate107inter4));
  nand2 gate888(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate889(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate890(.a(G366), .O(gate107inter7));
  inv1  gate891(.a(G367), .O(gate107inter8));
  nand2 gate892(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate893(.a(s_49), .b(gate107inter3), .O(gate107inter10));
  nor2  gate894(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate895(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate896(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate813(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate814(.a(gate109inter0), .b(s_38), .O(gate109inter1));
  and2  gate815(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate816(.a(s_38), .O(gate109inter3));
  inv1  gate817(.a(s_39), .O(gate109inter4));
  nand2 gate818(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate819(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate820(.a(G370), .O(gate109inter7));
  inv1  gate821(.a(G371), .O(gate109inter8));
  nand2 gate822(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate823(.a(s_39), .b(gate109inter3), .O(gate109inter10));
  nor2  gate824(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate825(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate826(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1709(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1710(.a(gate110inter0), .b(s_166), .O(gate110inter1));
  and2  gate1711(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1712(.a(s_166), .O(gate110inter3));
  inv1  gate1713(.a(s_167), .O(gate110inter4));
  nand2 gate1714(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1715(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1716(.a(G372), .O(gate110inter7));
  inv1  gate1717(.a(G373), .O(gate110inter8));
  nand2 gate1718(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1719(.a(s_167), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1720(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1721(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1722(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate785(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate786(.a(gate111inter0), .b(s_34), .O(gate111inter1));
  and2  gate787(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate788(.a(s_34), .O(gate111inter3));
  inv1  gate789(.a(s_35), .O(gate111inter4));
  nand2 gate790(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate791(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate792(.a(G374), .O(gate111inter7));
  inv1  gate793(.a(G375), .O(gate111inter8));
  nand2 gate794(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate795(.a(s_35), .b(gate111inter3), .O(gate111inter10));
  nor2  gate796(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate797(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate798(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1653(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1654(.a(gate115inter0), .b(s_158), .O(gate115inter1));
  and2  gate1655(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1656(.a(s_158), .O(gate115inter3));
  inv1  gate1657(.a(s_159), .O(gate115inter4));
  nand2 gate1658(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1659(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1660(.a(G382), .O(gate115inter7));
  inv1  gate1661(.a(G383), .O(gate115inter8));
  nand2 gate1662(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1663(.a(s_159), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1664(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1665(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1666(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1331(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1332(.a(gate116inter0), .b(s_112), .O(gate116inter1));
  and2  gate1333(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1334(.a(s_112), .O(gate116inter3));
  inv1  gate1335(.a(s_113), .O(gate116inter4));
  nand2 gate1336(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1337(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1338(.a(G384), .O(gate116inter7));
  inv1  gate1339(.a(G385), .O(gate116inter8));
  nand2 gate1340(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1341(.a(s_113), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1342(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1343(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1344(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1625(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1626(.a(gate117inter0), .b(s_154), .O(gate117inter1));
  and2  gate1627(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1628(.a(s_154), .O(gate117inter3));
  inv1  gate1629(.a(s_155), .O(gate117inter4));
  nand2 gate1630(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1631(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1632(.a(G386), .O(gate117inter7));
  inv1  gate1633(.a(G387), .O(gate117inter8));
  nand2 gate1634(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1635(.a(s_155), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1636(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1637(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1638(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate2465(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2466(.a(gate118inter0), .b(s_274), .O(gate118inter1));
  and2  gate2467(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2468(.a(s_274), .O(gate118inter3));
  inv1  gate2469(.a(s_275), .O(gate118inter4));
  nand2 gate2470(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2471(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2472(.a(G388), .O(gate118inter7));
  inv1  gate2473(.a(G389), .O(gate118inter8));
  nand2 gate2474(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2475(.a(s_275), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2476(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2477(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2478(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2045(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2046(.a(gate121inter0), .b(s_214), .O(gate121inter1));
  and2  gate2047(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2048(.a(s_214), .O(gate121inter3));
  inv1  gate2049(.a(s_215), .O(gate121inter4));
  nand2 gate2050(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2051(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2052(.a(G394), .O(gate121inter7));
  inv1  gate2053(.a(G395), .O(gate121inter8));
  nand2 gate2054(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2055(.a(s_215), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2056(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2057(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2058(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2017(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2018(.a(gate122inter0), .b(s_210), .O(gate122inter1));
  and2  gate2019(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2020(.a(s_210), .O(gate122inter3));
  inv1  gate2021(.a(s_211), .O(gate122inter4));
  nand2 gate2022(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2023(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2024(.a(G396), .O(gate122inter7));
  inv1  gate2025(.a(G397), .O(gate122inter8));
  nand2 gate2026(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2027(.a(s_211), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2028(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2029(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2030(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2129(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2130(.a(gate124inter0), .b(s_226), .O(gate124inter1));
  and2  gate2131(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2132(.a(s_226), .O(gate124inter3));
  inv1  gate2133(.a(s_227), .O(gate124inter4));
  nand2 gate2134(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2135(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2136(.a(G400), .O(gate124inter7));
  inv1  gate2137(.a(G401), .O(gate124inter8));
  nand2 gate2138(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2139(.a(s_227), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2140(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2141(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2142(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate575(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate576(.a(gate125inter0), .b(s_4), .O(gate125inter1));
  and2  gate577(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate578(.a(s_4), .O(gate125inter3));
  inv1  gate579(.a(s_5), .O(gate125inter4));
  nand2 gate580(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate581(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate582(.a(G402), .O(gate125inter7));
  inv1  gate583(.a(G403), .O(gate125inter8));
  nand2 gate584(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate585(.a(s_5), .b(gate125inter3), .O(gate125inter10));
  nor2  gate586(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate587(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate588(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate701(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate702(.a(gate127inter0), .b(s_22), .O(gate127inter1));
  and2  gate703(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate704(.a(s_22), .O(gate127inter3));
  inv1  gate705(.a(s_23), .O(gate127inter4));
  nand2 gate706(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate707(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate708(.a(G406), .O(gate127inter7));
  inv1  gate709(.a(G407), .O(gate127inter8));
  nand2 gate710(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate711(.a(s_23), .b(gate127inter3), .O(gate127inter10));
  nor2  gate712(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate713(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate714(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate2731(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2732(.a(gate130inter0), .b(s_312), .O(gate130inter1));
  and2  gate2733(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2734(.a(s_312), .O(gate130inter3));
  inv1  gate2735(.a(s_313), .O(gate130inter4));
  nand2 gate2736(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2737(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2738(.a(G412), .O(gate130inter7));
  inv1  gate2739(.a(G413), .O(gate130inter8));
  nand2 gate2740(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2741(.a(s_313), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2742(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2743(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2744(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2353(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2354(.a(gate131inter0), .b(s_258), .O(gate131inter1));
  and2  gate2355(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2356(.a(s_258), .O(gate131inter3));
  inv1  gate2357(.a(s_259), .O(gate131inter4));
  nand2 gate2358(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2359(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2360(.a(G414), .O(gate131inter7));
  inv1  gate2361(.a(G415), .O(gate131inter8));
  nand2 gate2362(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2363(.a(s_259), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2364(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2365(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2366(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1219(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1220(.a(gate139inter0), .b(s_96), .O(gate139inter1));
  and2  gate1221(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1222(.a(s_96), .O(gate139inter3));
  inv1  gate1223(.a(s_97), .O(gate139inter4));
  nand2 gate1224(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1225(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1226(.a(G438), .O(gate139inter7));
  inv1  gate1227(.a(G441), .O(gate139inter8));
  nand2 gate1228(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1229(.a(s_97), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1230(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1231(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1232(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2759(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2760(.a(gate143inter0), .b(s_316), .O(gate143inter1));
  and2  gate2761(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2762(.a(s_316), .O(gate143inter3));
  inv1  gate2763(.a(s_317), .O(gate143inter4));
  nand2 gate2764(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2765(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2766(.a(G462), .O(gate143inter7));
  inv1  gate2767(.a(G465), .O(gate143inter8));
  nand2 gate2768(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2769(.a(s_317), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2770(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2771(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2772(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2423(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2424(.a(gate147inter0), .b(s_268), .O(gate147inter1));
  and2  gate2425(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2426(.a(s_268), .O(gate147inter3));
  inv1  gate2427(.a(s_269), .O(gate147inter4));
  nand2 gate2428(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2429(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2430(.a(G486), .O(gate147inter7));
  inv1  gate2431(.a(G489), .O(gate147inter8));
  nand2 gate2432(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2433(.a(s_269), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2434(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2435(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2436(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1247(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1248(.a(gate148inter0), .b(s_100), .O(gate148inter1));
  and2  gate1249(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1250(.a(s_100), .O(gate148inter3));
  inv1  gate1251(.a(s_101), .O(gate148inter4));
  nand2 gate1252(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1253(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1254(.a(G492), .O(gate148inter7));
  inv1  gate1255(.a(G495), .O(gate148inter8));
  nand2 gate1256(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1257(.a(s_101), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1258(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1259(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1260(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate673(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate674(.a(gate149inter0), .b(s_18), .O(gate149inter1));
  and2  gate675(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate676(.a(s_18), .O(gate149inter3));
  inv1  gate677(.a(s_19), .O(gate149inter4));
  nand2 gate678(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate679(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate680(.a(G498), .O(gate149inter7));
  inv1  gate681(.a(G501), .O(gate149inter8));
  nand2 gate682(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate683(.a(s_19), .b(gate149inter3), .O(gate149inter10));
  nor2  gate684(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate685(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate686(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2339(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2340(.a(gate155inter0), .b(s_256), .O(gate155inter1));
  and2  gate2341(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2342(.a(s_256), .O(gate155inter3));
  inv1  gate2343(.a(s_257), .O(gate155inter4));
  nand2 gate2344(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2345(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2346(.a(G432), .O(gate155inter7));
  inv1  gate2347(.a(G525), .O(gate155inter8));
  nand2 gate2348(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2349(.a(s_257), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2350(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2351(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2352(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate743(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate744(.a(gate160inter0), .b(s_28), .O(gate160inter1));
  and2  gate745(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate746(.a(s_28), .O(gate160inter3));
  inv1  gate747(.a(s_29), .O(gate160inter4));
  nand2 gate748(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate749(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate750(.a(G447), .O(gate160inter7));
  inv1  gate751(.a(G531), .O(gate160inter8));
  nand2 gate752(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate753(.a(s_29), .b(gate160inter3), .O(gate160inter10));
  nor2  gate754(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate755(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate756(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate953(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate954(.a(gate162inter0), .b(s_58), .O(gate162inter1));
  and2  gate955(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate956(.a(s_58), .O(gate162inter3));
  inv1  gate957(.a(s_59), .O(gate162inter4));
  nand2 gate958(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate959(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate960(.a(G453), .O(gate162inter7));
  inv1  gate961(.a(G534), .O(gate162inter8));
  nand2 gate962(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate963(.a(s_59), .b(gate162inter3), .O(gate162inter10));
  nor2  gate964(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate965(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate966(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2073(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2074(.a(gate164inter0), .b(s_218), .O(gate164inter1));
  and2  gate2075(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2076(.a(s_218), .O(gate164inter3));
  inv1  gate2077(.a(s_219), .O(gate164inter4));
  nand2 gate2078(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2079(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2080(.a(G459), .O(gate164inter7));
  inv1  gate2081(.a(G537), .O(gate164inter8));
  nand2 gate2082(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2083(.a(s_219), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2084(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2085(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2086(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1485(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1486(.a(gate168inter0), .b(s_134), .O(gate168inter1));
  and2  gate1487(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1488(.a(s_134), .O(gate168inter3));
  inv1  gate1489(.a(s_135), .O(gate168inter4));
  nand2 gate1490(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1491(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1492(.a(G471), .O(gate168inter7));
  inv1  gate1493(.a(G543), .O(gate168inter8));
  nand2 gate1494(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1495(.a(s_135), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1496(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1497(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1498(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1947(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1948(.a(gate174inter0), .b(s_200), .O(gate174inter1));
  and2  gate1949(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1950(.a(s_200), .O(gate174inter3));
  inv1  gate1951(.a(s_201), .O(gate174inter4));
  nand2 gate1952(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1953(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1954(.a(G489), .O(gate174inter7));
  inv1  gate1955(.a(G552), .O(gate174inter8));
  nand2 gate1956(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1957(.a(s_201), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1958(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1959(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1960(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2605(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2606(.a(gate175inter0), .b(s_294), .O(gate175inter1));
  and2  gate2607(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2608(.a(s_294), .O(gate175inter3));
  inv1  gate2609(.a(s_295), .O(gate175inter4));
  nand2 gate2610(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2611(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2612(.a(G492), .O(gate175inter7));
  inv1  gate2613(.a(G555), .O(gate175inter8));
  nand2 gate2614(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2615(.a(s_295), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2616(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2617(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2618(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1359(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1360(.a(gate177inter0), .b(s_116), .O(gate177inter1));
  and2  gate1361(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1362(.a(s_116), .O(gate177inter3));
  inv1  gate1363(.a(s_117), .O(gate177inter4));
  nand2 gate1364(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1365(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1366(.a(G498), .O(gate177inter7));
  inv1  gate1367(.a(G558), .O(gate177inter8));
  nand2 gate1368(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1369(.a(s_117), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1370(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1371(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1372(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1723(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1724(.a(gate179inter0), .b(s_168), .O(gate179inter1));
  and2  gate1725(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1726(.a(s_168), .O(gate179inter3));
  inv1  gate1727(.a(s_169), .O(gate179inter4));
  nand2 gate1728(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1729(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1730(.a(G504), .O(gate179inter7));
  inv1  gate1731(.a(G561), .O(gate179inter8));
  nand2 gate1732(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1733(.a(s_169), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1734(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1735(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1736(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1149(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1150(.a(gate182inter0), .b(s_86), .O(gate182inter1));
  and2  gate1151(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1152(.a(s_86), .O(gate182inter3));
  inv1  gate1153(.a(s_87), .O(gate182inter4));
  nand2 gate1154(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1155(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1156(.a(G513), .O(gate182inter7));
  inv1  gate1157(.a(G564), .O(gate182inter8));
  nand2 gate1158(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1159(.a(s_87), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1160(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1161(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1162(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1415(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1416(.a(gate184inter0), .b(s_124), .O(gate184inter1));
  and2  gate1417(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1418(.a(s_124), .O(gate184inter3));
  inv1  gate1419(.a(s_125), .O(gate184inter4));
  nand2 gate1420(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1421(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1422(.a(G519), .O(gate184inter7));
  inv1  gate1423(.a(G567), .O(gate184inter8));
  nand2 gate1424(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1425(.a(s_125), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1426(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1427(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1428(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1891(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1892(.a(gate192inter0), .b(s_192), .O(gate192inter1));
  and2  gate1893(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1894(.a(s_192), .O(gate192inter3));
  inv1  gate1895(.a(s_193), .O(gate192inter4));
  nand2 gate1896(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1897(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1898(.a(G584), .O(gate192inter7));
  inv1  gate1899(.a(G585), .O(gate192inter8));
  nand2 gate1900(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1901(.a(s_193), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1902(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1903(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1904(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1821(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1822(.a(gate193inter0), .b(s_182), .O(gate193inter1));
  and2  gate1823(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1824(.a(s_182), .O(gate193inter3));
  inv1  gate1825(.a(s_183), .O(gate193inter4));
  nand2 gate1826(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1827(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1828(.a(G586), .O(gate193inter7));
  inv1  gate1829(.a(G587), .O(gate193inter8));
  nand2 gate1830(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1831(.a(s_183), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1832(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1833(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1834(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1499(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1500(.a(gate200inter0), .b(s_136), .O(gate200inter1));
  and2  gate1501(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1502(.a(s_136), .O(gate200inter3));
  inv1  gate1503(.a(s_137), .O(gate200inter4));
  nand2 gate1504(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1505(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1506(.a(G600), .O(gate200inter7));
  inv1  gate1507(.a(G601), .O(gate200inter8));
  nand2 gate1508(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1509(.a(s_137), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1510(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1511(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1512(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2185(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2186(.a(gate205inter0), .b(s_234), .O(gate205inter1));
  and2  gate2187(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2188(.a(s_234), .O(gate205inter3));
  inv1  gate2189(.a(s_235), .O(gate205inter4));
  nand2 gate2190(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2191(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2192(.a(G622), .O(gate205inter7));
  inv1  gate2193(.a(G627), .O(gate205inter8));
  nand2 gate2194(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2195(.a(s_235), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2196(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2197(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2198(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1779(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1780(.a(gate206inter0), .b(s_176), .O(gate206inter1));
  and2  gate1781(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1782(.a(s_176), .O(gate206inter3));
  inv1  gate1783(.a(s_177), .O(gate206inter4));
  nand2 gate1784(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1785(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1786(.a(G632), .O(gate206inter7));
  inv1  gate1787(.a(G637), .O(gate206inter8));
  nand2 gate1788(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1789(.a(s_177), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1790(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1791(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1792(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1737(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1738(.a(gate210inter0), .b(s_170), .O(gate210inter1));
  and2  gate1739(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1740(.a(s_170), .O(gate210inter3));
  inv1  gate1741(.a(s_171), .O(gate210inter4));
  nand2 gate1742(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1743(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1744(.a(G607), .O(gate210inter7));
  inv1  gate1745(.a(G666), .O(gate210inter8));
  nand2 gate1746(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1747(.a(s_171), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1748(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1749(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1750(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate981(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate982(.a(gate211inter0), .b(s_62), .O(gate211inter1));
  and2  gate983(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate984(.a(s_62), .O(gate211inter3));
  inv1  gate985(.a(s_63), .O(gate211inter4));
  nand2 gate986(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate987(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate988(.a(G612), .O(gate211inter7));
  inv1  gate989(.a(G669), .O(gate211inter8));
  nand2 gate990(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate991(.a(s_63), .b(gate211inter3), .O(gate211inter10));
  nor2  gate992(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate993(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate994(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2493(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2494(.a(gate214inter0), .b(s_278), .O(gate214inter1));
  and2  gate2495(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2496(.a(s_278), .O(gate214inter3));
  inv1  gate2497(.a(s_279), .O(gate214inter4));
  nand2 gate2498(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2499(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2500(.a(G612), .O(gate214inter7));
  inv1  gate2501(.a(G672), .O(gate214inter8));
  nand2 gate2502(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2503(.a(s_279), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2504(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2505(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2506(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2479(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2480(.a(gate215inter0), .b(s_276), .O(gate215inter1));
  and2  gate2481(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2482(.a(s_276), .O(gate215inter3));
  inv1  gate2483(.a(s_277), .O(gate215inter4));
  nand2 gate2484(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2485(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2486(.a(G607), .O(gate215inter7));
  inv1  gate2487(.a(G675), .O(gate215inter8));
  nand2 gate2488(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2489(.a(s_277), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2490(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2491(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2492(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1233(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1234(.a(gate221inter0), .b(s_98), .O(gate221inter1));
  and2  gate1235(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1236(.a(s_98), .O(gate221inter3));
  inv1  gate1237(.a(s_99), .O(gate221inter4));
  nand2 gate1238(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1239(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1240(.a(G622), .O(gate221inter7));
  inv1  gate1241(.a(G684), .O(gate221inter8));
  nand2 gate1242(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1243(.a(s_99), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1244(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1245(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1246(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate2311(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate2312(.a(gate226inter0), .b(s_252), .O(gate226inter1));
  and2  gate2313(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate2314(.a(s_252), .O(gate226inter3));
  inv1  gate2315(.a(s_253), .O(gate226inter4));
  nand2 gate2316(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate2317(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate2318(.a(G692), .O(gate226inter7));
  inv1  gate2319(.a(G693), .O(gate226inter8));
  nand2 gate2320(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate2321(.a(s_253), .b(gate226inter3), .O(gate226inter10));
  nor2  gate2322(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate2323(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate2324(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2535(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2536(.a(gate228inter0), .b(s_284), .O(gate228inter1));
  and2  gate2537(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2538(.a(s_284), .O(gate228inter3));
  inv1  gate2539(.a(s_285), .O(gate228inter4));
  nand2 gate2540(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2541(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2542(.a(G696), .O(gate228inter7));
  inv1  gate2543(.a(G697), .O(gate228inter8));
  nand2 gate2544(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2545(.a(s_285), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2546(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2547(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2548(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate799(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate800(.a(gate237inter0), .b(s_36), .O(gate237inter1));
  and2  gate801(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate802(.a(s_36), .O(gate237inter3));
  inv1  gate803(.a(s_37), .O(gate237inter4));
  nand2 gate804(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate805(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate806(.a(G254), .O(gate237inter7));
  inv1  gate807(.a(G706), .O(gate237inter8));
  nand2 gate808(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate809(.a(s_37), .b(gate237inter3), .O(gate237inter10));
  nor2  gate810(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate811(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate812(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate2115(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2116(.a(gate238inter0), .b(s_224), .O(gate238inter1));
  and2  gate2117(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2118(.a(s_224), .O(gate238inter3));
  inv1  gate2119(.a(s_225), .O(gate238inter4));
  nand2 gate2120(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2121(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2122(.a(G257), .O(gate238inter7));
  inv1  gate2123(.a(G709), .O(gate238inter8));
  nand2 gate2124(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2125(.a(s_225), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2126(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2127(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2128(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2619(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2620(.a(gate239inter0), .b(s_296), .O(gate239inter1));
  and2  gate2621(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2622(.a(s_296), .O(gate239inter3));
  inv1  gate2623(.a(s_297), .O(gate239inter4));
  nand2 gate2624(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2625(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2626(.a(G260), .O(gate239inter7));
  inv1  gate2627(.a(G712), .O(gate239inter8));
  nand2 gate2628(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2629(.a(s_297), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2630(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2631(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2632(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1303(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1304(.a(gate243inter0), .b(s_108), .O(gate243inter1));
  and2  gate1305(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1306(.a(s_108), .O(gate243inter3));
  inv1  gate1307(.a(s_109), .O(gate243inter4));
  nand2 gate1308(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1309(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1310(.a(G245), .O(gate243inter7));
  inv1  gate1311(.a(G733), .O(gate243inter8));
  nand2 gate1312(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1313(.a(s_109), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1314(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1315(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1316(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1093(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1094(.a(gate244inter0), .b(s_78), .O(gate244inter1));
  and2  gate1095(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1096(.a(s_78), .O(gate244inter3));
  inv1  gate1097(.a(s_79), .O(gate244inter4));
  nand2 gate1098(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1099(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1100(.a(G721), .O(gate244inter7));
  inv1  gate1101(.a(G733), .O(gate244inter8));
  nand2 gate1102(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1103(.a(s_79), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1104(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1105(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1106(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2633(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2634(.a(gate248inter0), .b(s_298), .O(gate248inter1));
  and2  gate2635(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2636(.a(s_298), .O(gate248inter3));
  inv1  gate2637(.a(s_299), .O(gate248inter4));
  nand2 gate2638(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2639(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2640(.a(G727), .O(gate248inter7));
  inv1  gate2641(.a(G739), .O(gate248inter8));
  nand2 gate2642(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2643(.a(s_299), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2644(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2645(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2646(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1989(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1990(.a(gate251inter0), .b(s_206), .O(gate251inter1));
  and2  gate1991(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1992(.a(s_206), .O(gate251inter3));
  inv1  gate1993(.a(s_207), .O(gate251inter4));
  nand2 gate1994(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1995(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1996(.a(G257), .O(gate251inter7));
  inv1  gate1997(.a(G745), .O(gate251inter8));
  nand2 gate1998(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1999(.a(s_207), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2000(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2001(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2002(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1121(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1122(.a(gate254inter0), .b(s_82), .O(gate254inter1));
  and2  gate1123(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1124(.a(s_82), .O(gate254inter3));
  inv1  gate1125(.a(s_83), .O(gate254inter4));
  nand2 gate1126(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1127(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1128(.a(G712), .O(gate254inter7));
  inv1  gate1129(.a(G748), .O(gate254inter8));
  nand2 gate1130(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1131(.a(s_83), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1132(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1133(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1134(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1009(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1010(.a(gate255inter0), .b(s_66), .O(gate255inter1));
  and2  gate1011(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1012(.a(s_66), .O(gate255inter3));
  inv1  gate1013(.a(s_67), .O(gate255inter4));
  nand2 gate1014(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1015(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1016(.a(G263), .O(gate255inter7));
  inv1  gate1017(.a(G751), .O(gate255inter8));
  nand2 gate1018(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1019(.a(s_67), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1020(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1021(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1022(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1345(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1346(.a(gate257inter0), .b(s_114), .O(gate257inter1));
  and2  gate1347(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1348(.a(s_114), .O(gate257inter3));
  inv1  gate1349(.a(s_115), .O(gate257inter4));
  nand2 gate1350(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1351(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1352(.a(G754), .O(gate257inter7));
  inv1  gate1353(.a(G755), .O(gate257inter8));
  nand2 gate1354(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1355(.a(s_115), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1356(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1357(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1358(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate869(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate870(.a(gate258inter0), .b(s_46), .O(gate258inter1));
  and2  gate871(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate872(.a(s_46), .O(gate258inter3));
  inv1  gate873(.a(s_47), .O(gate258inter4));
  nand2 gate874(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate875(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate876(.a(G756), .O(gate258inter7));
  inv1  gate877(.a(G757), .O(gate258inter8));
  nand2 gate878(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate879(.a(s_47), .b(gate258inter3), .O(gate258inter10));
  nor2  gate880(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate881(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate882(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1807(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1808(.a(gate259inter0), .b(s_180), .O(gate259inter1));
  and2  gate1809(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1810(.a(s_180), .O(gate259inter3));
  inv1  gate1811(.a(s_181), .O(gate259inter4));
  nand2 gate1812(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1813(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1814(.a(G758), .O(gate259inter7));
  inv1  gate1815(.a(G759), .O(gate259inter8));
  nand2 gate1816(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1817(.a(s_181), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1818(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1819(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1820(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate967(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate968(.a(gate260inter0), .b(s_60), .O(gate260inter1));
  and2  gate969(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate970(.a(s_60), .O(gate260inter3));
  inv1  gate971(.a(s_61), .O(gate260inter4));
  nand2 gate972(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate973(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate974(.a(G760), .O(gate260inter7));
  inv1  gate975(.a(G761), .O(gate260inter8));
  nand2 gate976(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate977(.a(s_61), .b(gate260inter3), .O(gate260inter10));
  nor2  gate978(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate979(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate980(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1065(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1066(.a(gate265inter0), .b(s_74), .O(gate265inter1));
  and2  gate1067(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1068(.a(s_74), .O(gate265inter3));
  inv1  gate1069(.a(s_75), .O(gate265inter4));
  nand2 gate1070(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1071(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1072(.a(G642), .O(gate265inter7));
  inv1  gate1073(.a(G770), .O(gate265inter8));
  nand2 gate1074(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1075(.a(s_75), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1076(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1077(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1078(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1527(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1528(.a(gate266inter0), .b(s_140), .O(gate266inter1));
  and2  gate1529(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1530(.a(s_140), .O(gate266inter3));
  inv1  gate1531(.a(s_141), .O(gate266inter4));
  nand2 gate1532(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1533(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1534(.a(G645), .O(gate266inter7));
  inv1  gate1535(.a(G773), .O(gate266inter8));
  nand2 gate1536(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1537(.a(s_141), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1538(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1539(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1540(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1513(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1514(.a(gate267inter0), .b(s_138), .O(gate267inter1));
  and2  gate1515(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1516(.a(s_138), .O(gate267inter3));
  inv1  gate1517(.a(s_139), .O(gate267inter4));
  nand2 gate1518(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1519(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1520(.a(G648), .O(gate267inter7));
  inv1  gate1521(.a(G776), .O(gate267inter8));
  nand2 gate1522(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1523(.a(s_139), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1524(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1525(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1526(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1961(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1962(.a(gate268inter0), .b(s_202), .O(gate268inter1));
  and2  gate1963(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1964(.a(s_202), .O(gate268inter3));
  inv1  gate1965(.a(s_203), .O(gate268inter4));
  nand2 gate1966(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1967(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1968(.a(G651), .O(gate268inter7));
  inv1  gate1969(.a(G779), .O(gate268inter8));
  nand2 gate1970(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1971(.a(s_203), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1972(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1973(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1974(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2647(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2648(.a(gate269inter0), .b(s_300), .O(gate269inter1));
  and2  gate2649(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2650(.a(s_300), .O(gate269inter3));
  inv1  gate2651(.a(s_301), .O(gate269inter4));
  nand2 gate2652(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2653(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2654(.a(G654), .O(gate269inter7));
  inv1  gate2655(.a(G782), .O(gate269inter8));
  nand2 gate2656(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2657(.a(s_301), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2658(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2659(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2660(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2325(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2326(.a(gate275inter0), .b(s_254), .O(gate275inter1));
  and2  gate2327(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2328(.a(s_254), .O(gate275inter3));
  inv1  gate2329(.a(s_255), .O(gate275inter4));
  nand2 gate2330(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2331(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2332(.a(G645), .O(gate275inter7));
  inv1  gate2333(.a(G797), .O(gate275inter8));
  nand2 gate2334(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2335(.a(s_255), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2336(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2337(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2338(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1289(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1290(.a(gate277inter0), .b(s_106), .O(gate277inter1));
  and2  gate1291(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1292(.a(s_106), .O(gate277inter3));
  inv1  gate1293(.a(s_107), .O(gate277inter4));
  nand2 gate1294(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1295(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1296(.a(G648), .O(gate277inter7));
  inv1  gate1297(.a(G800), .O(gate277inter8));
  nand2 gate1298(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1299(.a(s_107), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1300(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1301(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1302(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate897(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate898(.a(gate282inter0), .b(s_50), .O(gate282inter1));
  and2  gate899(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate900(.a(s_50), .O(gate282inter3));
  inv1  gate901(.a(s_51), .O(gate282inter4));
  nand2 gate902(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate903(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate904(.a(G782), .O(gate282inter7));
  inv1  gate905(.a(G806), .O(gate282inter8));
  nand2 gate906(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate907(.a(s_51), .b(gate282inter3), .O(gate282inter10));
  nor2  gate908(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate909(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate910(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1695(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1696(.a(gate285inter0), .b(s_164), .O(gate285inter1));
  and2  gate1697(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1698(.a(s_164), .O(gate285inter3));
  inv1  gate1699(.a(s_165), .O(gate285inter4));
  nand2 gate1700(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1701(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1702(.a(G660), .O(gate285inter7));
  inv1  gate1703(.a(G812), .O(gate285inter8));
  nand2 gate1704(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1705(.a(s_165), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1706(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1707(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1708(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2507(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2508(.a(gate286inter0), .b(s_280), .O(gate286inter1));
  and2  gate2509(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2510(.a(s_280), .O(gate286inter3));
  inv1  gate2511(.a(s_281), .O(gate286inter4));
  nand2 gate2512(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2513(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2514(.a(G788), .O(gate286inter7));
  inv1  gate2515(.a(G812), .O(gate286inter8));
  nand2 gate2516(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2517(.a(s_281), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2518(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2519(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2520(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2171(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2172(.a(gate287inter0), .b(s_232), .O(gate287inter1));
  and2  gate2173(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2174(.a(s_232), .O(gate287inter3));
  inv1  gate2175(.a(s_233), .O(gate287inter4));
  nand2 gate2176(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2177(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2178(.a(G663), .O(gate287inter7));
  inv1  gate2179(.a(G815), .O(gate287inter8));
  nand2 gate2180(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2181(.a(s_233), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2182(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2183(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2184(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1541(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1542(.a(gate288inter0), .b(s_142), .O(gate288inter1));
  and2  gate1543(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1544(.a(s_142), .O(gate288inter3));
  inv1  gate1545(.a(s_143), .O(gate288inter4));
  nand2 gate1546(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1547(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1548(.a(G791), .O(gate288inter7));
  inv1  gate1549(.a(G815), .O(gate288inter8));
  nand2 gate1550(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1551(.a(s_143), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1552(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1553(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1554(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1597(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1598(.a(gate290inter0), .b(s_150), .O(gate290inter1));
  and2  gate1599(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1600(.a(s_150), .O(gate290inter3));
  inv1  gate1601(.a(s_151), .O(gate290inter4));
  nand2 gate1602(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1603(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1604(.a(G820), .O(gate290inter7));
  inv1  gate1605(.a(G821), .O(gate290inter8));
  nand2 gate1606(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1607(.a(s_151), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1608(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1609(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1610(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1429(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1430(.a(gate291inter0), .b(s_126), .O(gate291inter1));
  and2  gate1431(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1432(.a(s_126), .O(gate291inter3));
  inv1  gate1433(.a(s_127), .O(gate291inter4));
  nand2 gate1434(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1435(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1436(.a(G822), .O(gate291inter7));
  inv1  gate1437(.a(G823), .O(gate291inter8));
  nand2 gate1438(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1439(.a(s_127), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1440(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1441(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1442(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1905(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1906(.a(gate292inter0), .b(s_194), .O(gate292inter1));
  and2  gate1907(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1908(.a(s_194), .O(gate292inter3));
  inv1  gate1909(.a(s_195), .O(gate292inter4));
  nand2 gate1910(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1911(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1912(.a(G824), .O(gate292inter7));
  inv1  gate1913(.a(G825), .O(gate292inter8));
  nand2 gate1914(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1915(.a(s_195), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1916(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1917(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1918(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate645(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate646(.a(gate293inter0), .b(s_14), .O(gate293inter1));
  and2  gate647(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate648(.a(s_14), .O(gate293inter3));
  inv1  gate649(.a(s_15), .O(gate293inter4));
  nand2 gate650(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate651(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate652(.a(G828), .O(gate293inter7));
  inv1  gate653(.a(G829), .O(gate293inter8));
  nand2 gate654(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate655(.a(s_15), .b(gate293inter3), .O(gate293inter10));
  nor2  gate656(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate657(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate658(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2003(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2004(.a(gate294inter0), .b(s_208), .O(gate294inter1));
  and2  gate2005(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2006(.a(s_208), .O(gate294inter3));
  inv1  gate2007(.a(s_209), .O(gate294inter4));
  nand2 gate2008(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2009(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2010(.a(G832), .O(gate294inter7));
  inv1  gate2011(.a(G833), .O(gate294inter8));
  nand2 gate2012(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2013(.a(s_209), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2014(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2015(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2016(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1751(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1752(.a(gate391inter0), .b(s_172), .O(gate391inter1));
  and2  gate1753(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1754(.a(s_172), .O(gate391inter3));
  inv1  gate1755(.a(s_173), .O(gate391inter4));
  nand2 gate1756(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1757(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1758(.a(G5), .O(gate391inter7));
  inv1  gate1759(.a(G1048), .O(gate391inter8));
  nand2 gate1760(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1761(.a(s_173), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1762(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1763(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1764(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate561(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate562(.a(gate392inter0), .b(s_2), .O(gate392inter1));
  and2  gate563(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate564(.a(s_2), .O(gate392inter3));
  inv1  gate565(.a(s_3), .O(gate392inter4));
  nand2 gate566(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate567(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate568(.a(G6), .O(gate392inter7));
  inv1  gate569(.a(G1051), .O(gate392inter8));
  nand2 gate570(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate571(.a(s_3), .b(gate392inter3), .O(gate392inter10));
  nor2  gate572(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate573(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate574(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate2059(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2060(.a(gate393inter0), .b(s_216), .O(gate393inter1));
  and2  gate2061(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2062(.a(s_216), .O(gate393inter3));
  inv1  gate2063(.a(s_217), .O(gate393inter4));
  nand2 gate2064(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2065(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2066(.a(G7), .O(gate393inter7));
  inv1  gate2067(.a(G1054), .O(gate393inter8));
  nand2 gate2068(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2069(.a(s_217), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2070(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2071(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2072(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1373(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1374(.a(gate398inter0), .b(s_118), .O(gate398inter1));
  and2  gate1375(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1376(.a(s_118), .O(gate398inter3));
  inv1  gate1377(.a(s_119), .O(gate398inter4));
  nand2 gate1378(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1379(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1380(.a(G12), .O(gate398inter7));
  inv1  gate1381(.a(G1069), .O(gate398inter8));
  nand2 gate1382(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1383(.a(s_119), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1384(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1385(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1386(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1765(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1766(.a(gate399inter0), .b(s_174), .O(gate399inter1));
  and2  gate1767(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1768(.a(s_174), .O(gate399inter3));
  inv1  gate1769(.a(s_175), .O(gate399inter4));
  nand2 gate1770(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1771(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1772(.a(G13), .O(gate399inter7));
  inv1  gate1773(.a(G1072), .O(gate399inter8));
  nand2 gate1774(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1775(.a(s_175), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1776(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1777(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1778(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2297(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2298(.a(gate401inter0), .b(s_250), .O(gate401inter1));
  and2  gate2299(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2300(.a(s_250), .O(gate401inter3));
  inv1  gate2301(.a(s_251), .O(gate401inter4));
  nand2 gate2302(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2303(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2304(.a(G15), .O(gate401inter7));
  inv1  gate2305(.a(G1078), .O(gate401inter8));
  nand2 gate2306(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2307(.a(s_251), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2308(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2309(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2310(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate855(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate856(.a(gate403inter0), .b(s_44), .O(gate403inter1));
  and2  gate857(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate858(.a(s_44), .O(gate403inter3));
  inv1  gate859(.a(s_45), .O(gate403inter4));
  nand2 gate860(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate861(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate862(.a(G17), .O(gate403inter7));
  inv1  gate863(.a(G1084), .O(gate403inter8));
  nand2 gate864(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate865(.a(s_45), .b(gate403inter3), .O(gate403inter10));
  nor2  gate866(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate867(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate868(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate757(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate758(.a(gate405inter0), .b(s_30), .O(gate405inter1));
  and2  gate759(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate760(.a(s_30), .O(gate405inter3));
  inv1  gate761(.a(s_31), .O(gate405inter4));
  nand2 gate762(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate763(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate764(.a(G19), .O(gate405inter7));
  inv1  gate765(.a(G1090), .O(gate405inter8));
  nand2 gate766(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate767(.a(s_31), .b(gate405inter3), .O(gate405inter10));
  nor2  gate768(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate769(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate770(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2717(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2718(.a(gate406inter0), .b(s_310), .O(gate406inter1));
  and2  gate2719(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2720(.a(s_310), .O(gate406inter3));
  inv1  gate2721(.a(s_311), .O(gate406inter4));
  nand2 gate2722(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2723(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2724(.a(G20), .O(gate406inter7));
  inv1  gate2725(.a(G1093), .O(gate406inter8));
  nand2 gate2726(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2727(.a(s_311), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2728(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2729(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2730(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2773(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2774(.a(gate408inter0), .b(s_318), .O(gate408inter1));
  and2  gate2775(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2776(.a(s_318), .O(gate408inter3));
  inv1  gate2777(.a(s_319), .O(gate408inter4));
  nand2 gate2778(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2779(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2780(.a(G22), .O(gate408inter7));
  inv1  gate2781(.a(G1099), .O(gate408inter8));
  nand2 gate2782(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2783(.a(s_319), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2784(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2785(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2786(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1387(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1388(.a(gate410inter0), .b(s_120), .O(gate410inter1));
  and2  gate1389(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1390(.a(s_120), .O(gate410inter3));
  inv1  gate1391(.a(s_121), .O(gate410inter4));
  nand2 gate1392(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1393(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1394(.a(G24), .O(gate410inter7));
  inv1  gate1395(.a(G1105), .O(gate410inter8));
  nand2 gate1396(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1397(.a(s_121), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1398(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1399(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1400(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1849(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1850(.a(gate411inter0), .b(s_186), .O(gate411inter1));
  and2  gate1851(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1852(.a(s_186), .O(gate411inter3));
  inv1  gate1853(.a(s_187), .O(gate411inter4));
  nand2 gate1854(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1855(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1856(.a(G25), .O(gate411inter7));
  inv1  gate1857(.a(G1108), .O(gate411inter8));
  nand2 gate1858(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1859(.a(s_187), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1860(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1861(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1862(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate995(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate996(.a(gate412inter0), .b(s_64), .O(gate412inter1));
  and2  gate997(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate998(.a(s_64), .O(gate412inter3));
  inv1  gate999(.a(s_65), .O(gate412inter4));
  nand2 gate1000(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1001(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1002(.a(G26), .O(gate412inter7));
  inv1  gate1003(.a(G1111), .O(gate412inter8));
  nand2 gate1004(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1005(.a(s_65), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1006(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1007(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1008(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2563(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2564(.a(gate414inter0), .b(s_288), .O(gate414inter1));
  and2  gate2565(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2566(.a(s_288), .O(gate414inter3));
  inv1  gate2567(.a(s_289), .O(gate414inter4));
  nand2 gate2568(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2569(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2570(.a(G28), .O(gate414inter7));
  inv1  gate2571(.a(G1117), .O(gate414inter8));
  nand2 gate2572(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2573(.a(s_289), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2574(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2575(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2576(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate729(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate730(.a(gate418inter0), .b(s_26), .O(gate418inter1));
  and2  gate731(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate732(.a(s_26), .O(gate418inter3));
  inv1  gate733(.a(s_27), .O(gate418inter4));
  nand2 gate734(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate735(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate736(.a(G32), .O(gate418inter7));
  inv1  gate737(.a(G1129), .O(gate418inter8));
  nand2 gate738(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate739(.a(s_27), .b(gate418inter3), .O(gate418inter10));
  nor2  gate740(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate741(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate742(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1023(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1024(.a(gate419inter0), .b(s_68), .O(gate419inter1));
  and2  gate1025(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1026(.a(s_68), .O(gate419inter3));
  inv1  gate1027(.a(s_69), .O(gate419inter4));
  nand2 gate1028(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1029(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1030(.a(G1), .O(gate419inter7));
  inv1  gate1031(.a(G1132), .O(gate419inter8));
  nand2 gate1032(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1033(.a(s_69), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1034(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1035(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1036(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate771(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate772(.a(gate420inter0), .b(s_32), .O(gate420inter1));
  and2  gate773(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate774(.a(s_32), .O(gate420inter3));
  inv1  gate775(.a(s_33), .O(gate420inter4));
  nand2 gate776(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate777(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate778(.a(G1036), .O(gate420inter7));
  inv1  gate779(.a(G1132), .O(gate420inter8));
  nand2 gate780(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate781(.a(s_33), .b(gate420inter3), .O(gate420inter10));
  nor2  gate782(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate783(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate784(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate603(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate604(.a(gate422inter0), .b(s_8), .O(gate422inter1));
  and2  gate605(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate606(.a(s_8), .O(gate422inter3));
  inv1  gate607(.a(s_9), .O(gate422inter4));
  nand2 gate608(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate609(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate610(.a(G1039), .O(gate422inter7));
  inv1  gate611(.a(G1135), .O(gate422inter8));
  nand2 gate612(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate613(.a(s_9), .b(gate422inter3), .O(gate422inter10));
  nor2  gate614(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate615(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate616(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2283(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2284(.a(gate426inter0), .b(s_248), .O(gate426inter1));
  and2  gate2285(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2286(.a(s_248), .O(gate426inter3));
  inv1  gate2287(.a(s_249), .O(gate426inter4));
  nand2 gate2288(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2289(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2290(.a(G1045), .O(gate426inter7));
  inv1  gate2291(.a(G1141), .O(gate426inter8));
  nand2 gate2292(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2293(.a(s_249), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2294(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2295(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2296(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2087(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2088(.a(gate427inter0), .b(s_220), .O(gate427inter1));
  and2  gate2089(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2090(.a(s_220), .O(gate427inter3));
  inv1  gate2091(.a(s_221), .O(gate427inter4));
  nand2 gate2092(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2093(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2094(.a(G5), .O(gate427inter7));
  inv1  gate2095(.a(G1144), .O(gate427inter8));
  nand2 gate2096(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2097(.a(s_221), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2098(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2099(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2100(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2213(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2214(.a(gate429inter0), .b(s_238), .O(gate429inter1));
  and2  gate2215(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2216(.a(s_238), .O(gate429inter3));
  inv1  gate2217(.a(s_239), .O(gate429inter4));
  nand2 gate2218(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2219(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2220(.a(G6), .O(gate429inter7));
  inv1  gate2221(.a(G1147), .O(gate429inter8));
  nand2 gate2222(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2223(.a(s_239), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2224(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2225(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2226(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1191(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1192(.a(gate433inter0), .b(s_92), .O(gate433inter1));
  and2  gate1193(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1194(.a(s_92), .O(gate433inter3));
  inv1  gate1195(.a(s_93), .O(gate433inter4));
  nand2 gate1196(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1197(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1198(.a(G8), .O(gate433inter7));
  inv1  gate1199(.a(G1153), .O(gate433inter8));
  nand2 gate1200(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1201(.a(s_93), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1202(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1203(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1204(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2367(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2368(.a(gate443inter0), .b(s_260), .O(gate443inter1));
  and2  gate2369(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2370(.a(s_260), .O(gate443inter3));
  inv1  gate2371(.a(s_261), .O(gate443inter4));
  nand2 gate2372(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2373(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2374(.a(G13), .O(gate443inter7));
  inv1  gate2375(.a(G1168), .O(gate443inter8));
  nand2 gate2376(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2377(.a(s_261), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2378(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2379(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2380(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2675(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2676(.a(gate444inter0), .b(s_304), .O(gate444inter1));
  and2  gate2677(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2678(.a(s_304), .O(gate444inter3));
  inv1  gate2679(.a(s_305), .O(gate444inter4));
  nand2 gate2680(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2681(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2682(.a(G1072), .O(gate444inter7));
  inv1  gate2683(.a(G1168), .O(gate444inter8));
  nand2 gate2684(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2685(.a(s_305), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2686(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2687(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2688(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2787(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2788(.a(gate448inter0), .b(s_320), .O(gate448inter1));
  and2  gate2789(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2790(.a(s_320), .O(gate448inter3));
  inv1  gate2791(.a(s_321), .O(gate448inter4));
  nand2 gate2792(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2793(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2794(.a(G1078), .O(gate448inter7));
  inv1  gate2795(.a(G1174), .O(gate448inter8));
  nand2 gate2796(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2797(.a(s_321), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2798(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2799(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2800(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2255(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2256(.a(gate450inter0), .b(s_244), .O(gate450inter1));
  and2  gate2257(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2258(.a(s_244), .O(gate450inter3));
  inv1  gate2259(.a(s_245), .O(gate450inter4));
  nand2 gate2260(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2261(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2262(.a(G1081), .O(gate450inter7));
  inv1  gate2263(.a(G1177), .O(gate450inter8));
  nand2 gate2264(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2265(.a(s_245), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2266(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2267(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2268(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2451(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2452(.a(gate452inter0), .b(s_272), .O(gate452inter1));
  and2  gate2453(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2454(.a(s_272), .O(gate452inter3));
  inv1  gate2455(.a(s_273), .O(gate452inter4));
  nand2 gate2456(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2457(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2458(.a(G1084), .O(gate452inter7));
  inv1  gate2459(.a(G1180), .O(gate452inter8));
  nand2 gate2460(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2461(.a(s_273), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2462(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2463(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2464(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1863(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1864(.a(gate455inter0), .b(s_188), .O(gate455inter1));
  and2  gate1865(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1866(.a(s_188), .O(gate455inter3));
  inv1  gate1867(.a(s_189), .O(gate455inter4));
  nand2 gate1868(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1869(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1870(.a(G19), .O(gate455inter7));
  inv1  gate1871(.a(G1186), .O(gate455inter8));
  nand2 gate1872(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1873(.a(s_189), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1874(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1875(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1876(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1275(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1276(.a(gate458inter0), .b(s_104), .O(gate458inter1));
  and2  gate1277(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1278(.a(s_104), .O(gate458inter3));
  inv1  gate1279(.a(s_105), .O(gate458inter4));
  nand2 gate1280(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1281(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1282(.a(G1093), .O(gate458inter7));
  inv1  gate1283(.a(G1189), .O(gate458inter8));
  nand2 gate1284(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1285(.a(s_105), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1286(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1287(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1288(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2241(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2242(.a(gate462inter0), .b(s_242), .O(gate462inter1));
  and2  gate2243(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2244(.a(s_242), .O(gate462inter3));
  inv1  gate2245(.a(s_243), .O(gate462inter4));
  nand2 gate2246(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2247(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2248(.a(G1099), .O(gate462inter7));
  inv1  gate2249(.a(G1195), .O(gate462inter8));
  nand2 gate2250(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2251(.a(s_243), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2252(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2253(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2254(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1583(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1584(.a(gate464inter0), .b(s_148), .O(gate464inter1));
  and2  gate1585(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1586(.a(s_148), .O(gate464inter3));
  inv1  gate1587(.a(s_149), .O(gate464inter4));
  nand2 gate1588(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1589(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1590(.a(G1102), .O(gate464inter7));
  inv1  gate1591(.a(G1198), .O(gate464inter8));
  nand2 gate1592(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1593(.a(s_149), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1594(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1595(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1596(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2227(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2228(.a(gate465inter0), .b(s_240), .O(gate465inter1));
  and2  gate2229(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2230(.a(s_240), .O(gate465inter3));
  inv1  gate2231(.a(s_241), .O(gate465inter4));
  nand2 gate2232(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2233(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2234(.a(G24), .O(gate465inter7));
  inv1  gate2235(.a(G1201), .O(gate465inter8));
  nand2 gate2236(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2237(.a(s_241), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2238(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2239(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2240(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1877(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1878(.a(gate468inter0), .b(s_190), .O(gate468inter1));
  and2  gate1879(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1880(.a(s_190), .O(gate468inter3));
  inv1  gate1881(.a(s_191), .O(gate468inter4));
  nand2 gate1882(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1883(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1884(.a(G1108), .O(gate468inter7));
  inv1  gate1885(.a(G1204), .O(gate468inter8));
  nand2 gate1886(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1887(.a(s_191), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1888(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1889(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1890(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1835(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1836(.a(gate470inter0), .b(s_184), .O(gate470inter1));
  and2  gate1837(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1838(.a(s_184), .O(gate470inter3));
  inv1  gate1839(.a(s_185), .O(gate470inter4));
  nand2 gate1840(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1841(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1842(.a(G1111), .O(gate470inter7));
  inv1  gate1843(.a(G1207), .O(gate470inter8));
  nand2 gate1844(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1845(.a(s_185), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1846(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1847(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1848(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1793(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1794(.a(gate472inter0), .b(s_178), .O(gate472inter1));
  and2  gate1795(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1796(.a(s_178), .O(gate472inter3));
  inv1  gate1797(.a(s_179), .O(gate472inter4));
  nand2 gate1798(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1799(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1800(.a(G1114), .O(gate472inter7));
  inv1  gate1801(.a(G1210), .O(gate472inter8));
  nand2 gate1802(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1803(.a(s_179), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1804(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1805(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1806(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2703(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2704(.a(gate474inter0), .b(s_308), .O(gate474inter1));
  and2  gate2705(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2706(.a(s_308), .O(gate474inter3));
  inv1  gate2707(.a(s_309), .O(gate474inter4));
  nand2 gate2708(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2709(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2710(.a(G1117), .O(gate474inter7));
  inv1  gate2711(.a(G1213), .O(gate474inter8));
  nand2 gate2712(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2713(.a(s_309), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2714(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2715(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2716(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1163(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1164(.a(gate478inter0), .b(s_88), .O(gate478inter1));
  and2  gate1165(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1166(.a(s_88), .O(gate478inter3));
  inv1  gate1167(.a(s_89), .O(gate478inter4));
  nand2 gate1168(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1169(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1170(.a(G1123), .O(gate478inter7));
  inv1  gate1171(.a(G1219), .O(gate478inter8));
  nand2 gate1172(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1173(.a(s_89), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1174(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1175(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1176(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2381(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2382(.a(gate482inter0), .b(s_262), .O(gate482inter1));
  and2  gate2383(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2384(.a(s_262), .O(gate482inter3));
  inv1  gate2385(.a(s_263), .O(gate482inter4));
  nand2 gate2386(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2387(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2388(.a(G1129), .O(gate482inter7));
  inv1  gate2389(.a(G1225), .O(gate482inter8));
  nand2 gate2390(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2391(.a(s_263), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2392(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2393(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2394(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1667(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1668(.a(gate485inter0), .b(s_160), .O(gate485inter1));
  and2  gate1669(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1670(.a(s_160), .O(gate485inter3));
  inv1  gate1671(.a(s_161), .O(gate485inter4));
  nand2 gate1672(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1673(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1674(.a(G1232), .O(gate485inter7));
  inv1  gate1675(.a(G1233), .O(gate485inter8));
  nand2 gate1676(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1677(.a(s_161), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1678(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1679(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1680(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate2101(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2102(.a(gate486inter0), .b(s_222), .O(gate486inter1));
  and2  gate2103(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2104(.a(s_222), .O(gate486inter3));
  inv1  gate2105(.a(s_223), .O(gate486inter4));
  nand2 gate2106(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2107(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2108(.a(G1234), .O(gate486inter7));
  inv1  gate2109(.a(G1235), .O(gate486inter8));
  nand2 gate2110(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2111(.a(s_223), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2112(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2113(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2114(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate715(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate716(.a(gate487inter0), .b(s_24), .O(gate487inter1));
  and2  gate717(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate718(.a(s_24), .O(gate487inter3));
  inv1  gate719(.a(s_25), .O(gate487inter4));
  nand2 gate720(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate721(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate722(.a(G1236), .O(gate487inter7));
  inv1  gate723(.a(G1237), .O(gate487inter8));
  nand2 gate724(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate725(.a(s_25), .b(gate487inter3), .O(gate487inter10));
  nor2  gate726(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate727(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate728(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate547(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate548(.a(gate488inter0), .b(s_0), .O(gate488inter1));
  and2  gate549(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate550(.a(s_0), .O(gate488inter3));
  inv1  gate551(.a(s_1), .O(gate488inter4));
  nand2 gate552(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate553(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate554(.a(G1238), .O(gate488inter7));
  inv1  gate555(.a(G1239), .O(gate488inter8));
  nand2 gate556(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate557(.a(s_1), .b(gate488inter3), .O(gate488inter10));
  nor2  gate558(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate559(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate560(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate687(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate688(.a(gate492inter0), .b(s_20), .O(gate492inter1));
  and2  gate689(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate690(.a(s_20), .O(gate492inter3));
  inv1  gate691(.a(s_21), .O(gate492inter4));
  nand2 gate692(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate693(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate694(.a(G1246), .O(gate492inter7));
  inv1  gate695(.a(G1247), .O(gate492inter8));
  nand2 gate696(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate697(.a(s_21), .b(gate492inter3), .O(gate492inter10));
  nor2  gate698(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate699(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate700(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1401(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1402(.a(gate494inter0), .b(s_122), .O(gate494inter1));
  and2  gate1403(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1404(.a(s_122), .O(gate494inter3));
  inv1  gate1405(.a(s_123), .O(gate494inter4));
  nand2 gate1406(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1407(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1408(.a(G1250), .O(gate494inter7));
  inv1  gate1409(.a(G1251), .O(gate494inter8));
  nand2 gate1410(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1411(.a(s_123), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1412(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1413(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1414(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate925(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate926(.a(gate495inter0), .b(s_54), .O(gate495inter1));
  and2  gate927(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate928(.a(s_54), .O(gate495inter3));
  inv1  gate929(.a(s_55), .O(gate495inter4));
  nand2 gate930(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate931(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate932(.a(G1252), .O(gate495inter7));
  inv1  gate933(.a(G1253), .O(gate495inter8));
  nand2 gate934(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate935(.a(s_55), .b(gate495inter3), .O(gate495inter10));
  nor2  gate936(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate937(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate938(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate617(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate618(.a(gate497inter0), .b(s_10), .O(gate497inter1));
  and2  gate619(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate620(.a(s_10), .O(gate497inter3));
  inv1  gate621(.a(s_11), .O(gate497inter4));
  nand2 gate622(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate623(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate624(.a(G1256), .O(gate497inter7));
  inv1  gate625(.a(G1257), .O(gate497inter8));
  nand2 gate626(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate627(.a(s_11), .b(gate497inter3), .O(gate497inter10));
  nor2  gate628(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate629(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate630(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1107(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1108(.a(gate499inter0), .b(s_80), .O(gate499inter1));
  and2  gate1109(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1110(.a(s_80), .O(gate499inter3));
  inv1  gate1111(.a(s_81), .O(gate499inter4));
  nand2 gate1112(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1113(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1114(.a(G1260), .O(gate499inter7));
  inv1  gate1115(.a(G1261), .O(gate499inter8));
  nand2 gate1116(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1117(.a(s_81), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1118(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1119(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1120(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate2661(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2662(.a(gate504inter0), .b(s_302), .O(gate504inter1));
  and2  gate2663(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2664(.a(s_302), .O(gate504inter3));
  inv1  gate2665(.a(s_303), .O(gate504inter4));
  nand2 gate2666(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2667(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2668(.a(G1270), .O(gate504inter7));
  inv1  gate2669(.a(G1271), .O(gate504inter8));
  nand2 gate2670(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2671(.a(s_303), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2672(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2673(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2674(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1975(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1976(.a(gate507inter0), .b(s_204), .O(gate507inter1));
  and2  gate1977(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1978(.a(s_204), .O(gate507inter3));
  inv1  gate1979(.a(s_205), .O(gate507inter4));
  nand2 gate1980(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1981(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1982(.a(G1276), .O(gate507inter7));
  inv1  gate1983(.a(G1277), .O(gate507inter8));
  nand2 gate1984(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1985(.a(s_205), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1986(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1987(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1988(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1037(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1038(.a(gate508inter0), .b(s_70), .O(gate508inter1));
  and2  gate1039(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1040(.a(s_70), .O(gate508inter3));
  inv1  gate1041(.a(s_71), .O(gate508inter4));
  nand2 gate1042(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1043(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1044(.a(G1278), .O(gate508inter7));
  inv1  gate1045(.a(G1279), .O(gate508inter8));
  nand2 gate1046(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1047(.a(s_71), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1048(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1049(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1050(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2437(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2438(.a(gate510inter0), .b(s_270), .O(gate510inter1));
  and2  gate2439(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2440(.a(s_270), .O(gate510inter3));
  inv1  gate2441(.a(s_271), .O(gate510inter4));
  nand2 gate2442(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2443(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2444(.a(G1282), .O(gate510inter7));
  inv1  gate2445(.a(G1283), .O(gate510inter8));
  nand2 gate2446(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2447(.a(s_271), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2448(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2449(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2450(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate2143(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2144(.a(gate511inter0), .b(s_228), .O(gate511inter1));
  and2  gate2145(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2146(.a(s_228), .O(gate511inter3));
  inv1  gate2147(.a(s_229), .O(gate511inter4));
  nand2 gate2148(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2149(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2150(.a(G1284), .O(gate511inter7));
  inv1  gate2151(.a(G1285), .O(gate511inter8));
  nand2 gate2152(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2153(.a(s_229), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2154(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2155(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2156(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule