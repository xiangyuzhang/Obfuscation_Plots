module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1149(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1150(.a(gate24inter0), .b(s_86), .O(gate24inter1));
  and2  gate1151(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1152(.a(s_86), .O(gate24inter3));
  inv1  gate1153(.a(s_87), .O(gate24inter4));
  nand2 gate1154(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1155(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1156(.a(G31), .O(gate24inter7));
  inv1  gate1157(.a(G32), .O(gate24inter8));
  nand2 gate1158(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1159(.a(s_87), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1160(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1161(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1162(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate771(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate772(.a(gate43inter0), .b(s_32), .O(gate43inter1));
  and2  gate773(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate774(.a(s_32), .O(gate43inter3));
  inv1  gate775(.a(s_33), .O(gate43inter4));
  nand2 gate776(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate777(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate778(.a(G3), .O(gate43inter7));
  inv1  gate779(.a(G269), .O(gate43inter8));
  nand2 gate780(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate781(.a(s_33), .b(gate43inter3), .O(gate43inter10));
  nor2  gate782(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate783(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate784(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate743(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate744(.a(gate62inter0), .b(s_28), .O(gate62inter1));
  and2  gate745(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate746(.a(s_28), .O(gate62inter3));
  inv1  gate747(.a(s_29), .O(gate62inter4));
  nand2 gate748(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate749(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate750(.a(G22), .O(gate62inter7));
  inv1  gate751(.a(G296), .O(gate62inter8));
  nand2 gate752(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate753(.a(s_29), .b(gate62inter3), .O(gate62inter10));
  nor2  gate754(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate755(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate756(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate925(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate926(.a(gate65inter0), .b(s_54), .O(gate65inter1));
  and2  gate927(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate928(.a(s_54), .O(gate65inter3));
  inv1  gate929(.a(s_55), .O(gate65inter4));
  nand2 gate930(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate931(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate932(.a(G25), .O(gate65inter7));
  inv1  gate933(.a(G302), .O(gate65inter8));
  nand2 gate934(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate935(.a(s_55), .b(gate65inter3), .O(gate65inter10));
  nor2  gate936(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate937(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate938(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1079(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1080(.a(gate68inter0), .b(s_76), .O(gate68inter1));
  and2  gate1081(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1082(.a(s_76), .O(gate68inter3));
  inv1  gate1083(.a(s_77), .O(gate68inter4));
  nand2 gate1084(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1085(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1086(.a(G28), .O(gate68inter7));
  inv1  gate1087(.a(G305), .O(gate68inter8));
  nand2 gate1088(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1089(.a(s_77), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1090(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1091(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1092(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate953(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate954(.a(gate74inter0), .b(s_58), .O(gate74inter1));
  and2  gate955(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate956(.a(s_58), .O(gate74inter3));
  inv1  gate957(.a(s_59), .O(gate74inter4));
  nand2 gate958(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate959(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate960(.a(G5), .O(gate74inter7));
  inv1  gate961(.a(G314), .O(gate74inter8));
  nand2 gate962(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate963(.a(s_59), .b(gate74inter3), .O(gate74inter10));
  nor2  gate964(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate965(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate966(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate701(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate702(.a(gate75inter0), .b(s_22), .O(gate75inter1));
  and2  gate703(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate704(.a(s_22), .O(gate75inter3));
  inv1  gate705(.a(s_23), .O(gate75inter4));
  nand2 gate706(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate707(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate708(.a(G9), .O(gate75inter7));
  inv1  gate709(.a(G317), .O(gate75inter8));
  nand2 gate710(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate711(.a(s_23), .b(gate75inter3), .O(gate75inter10));
  nor2  gate712(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate713(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate714(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate673(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate674(.a(gate77inter0), .b(s_18), .O(gate77inter1));
  and2  gate675(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate676(.a(s_18), .O(gate77inter3));
  inv1  gate677(.a(s_19), .O(gate77inter4));
  nand2 gate678(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate679(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate680(.a(G2), .O(gate77inter7));
  inv1  gate681(.a(G320), .O(gate77inter8));
  nand2 gate682(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate683(.a(s_19), .b(gate77inter3), .O(gate77inter10));
  nor2  gate684(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate685(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate686(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate785(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate786(.a(gate79inter0), .b(s_34), .O(gate79inter1));
  and2  gate787(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate788(.a(s_34), .O(gate79inter3));
  inv1  gate789(.a(s_35), .O(gate79inter4));
  nand2 gate790(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate791(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate792(.a(G10), .O(gate79inter7));
  inv1  gate793(.a(G323), .O(gate79inter8));
  nand2 gate794(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate795(.a(s_35), .b(gate79inter3), .O(gate79inter10));
  nor2  gate796(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate797(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate798(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate841(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate842(.a(gate81inter0), .b(s_42), .O(gate81inter1));
  and2  gate843(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate844(.a(s_42), .O(gate81inter3));
  inv1  gate845(.a(s_43), .O(gate81inter4));
  nand2 gate846(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate847(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate848(.a(G3), .O(gate81inter7));
  inv1  gate849(.a(G326), .O(gate81inter8));
  nand2 gate850(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate851(.a(s_43), .b(gate81inter3), .O(gate81inter10));
  nor2  gate852(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate853(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate854(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1065(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1066(.a(gate123inter0), .b(s_74), .O(gate123inter1));
  and2  gate1067(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1068(.a(s_74), .O(gate123inter3));
  inv1  gate1069(.a(s_75), .O(gate123inter4));
  nand2 gate1070(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1071(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1072(.a(G398), .O(gate123inter7));
  inv1  gate1073(.a(G399), .O(gate123inter8));
  nand2 gate1074(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1075(.a(s_75), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1076(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1077(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1078(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate575(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate576(.a(gate154inter0), .b(s_4), .O(gate154inter1));
  and2  gate577(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate578(.a(s_4), .O(gate154inter3));
  inv1  gate579(.a(s_5), .O(gate154inter4));
  nand2 gate580(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate581(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate582(.a(G429), .O(gate154inter7));
  inv1  gate583(.a(G522), .O(gate154inter8));
  nand2 gate584(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate585(.a(s_5), .b(gate154inter3), .O(gate154inter10));
  nor2  gate586(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate587(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate588(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate799(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate800(.a(gate155inter0), .b(s_36), .O(gate155inter1));
  and2  gate801(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate802(.a(s_36), .O(gate155inter3));
  inv1  gate803(.a(s_37), .O(gate155inter4));
  nand2 gate804(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate805(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate806(.a(G432), .O(gate155inter7));
  inv1  gate807(.a(G525), .O(gate155inter8));
  nand2 gate808(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate809(.a(s_37), .b(gate155inter3), .O(gate155inter10));
  nor2  gate810(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate811(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate812(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1037(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1038(.a(gate160inter0), .b(s_70), .O(gate160inter1));
  and2  gate1039(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1040(.a(s_70), .O(gate160inter3));
  inv1  gate1041(.a(s_71), .O(gate160inter4));
  nand2 gate1042(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1043(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1044(.a(G447), .O(gate160inter7));
  inv1  gate1045(.a(G531), .O(gate160inter8));
  nand2 gate1046(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1047(.a(s_71), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1048(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1049(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1050(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate603(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate604(.a(gate180inter0), .b(s_8), .O(gate180inter1));
  and2  gate605(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate606(.a(s_8), .O(gate180inter3));
  inv1  gate607(.a(s_9), .O(gate180inter4));
  nand2 gate608(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate609(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate610(.a(G507), .O(gate180inter7));
  inv1  gate611(.a(G561), .O(gate180inter8));
  nand2 gate612(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate613(.a(s_9), .b(gate180inter3), .O(gate180inter10));
  nor2  gate614(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate615(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate616(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1023(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1024(.a(gate182inter0), .b(s_68), .O(gate182inter1));
  and2  gate1025(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1026(.a(s_68), .O(gate182inter3));
  inv1  gate1027(.a(s_69), .O(gate182inter4));
  nand2 gate1028(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1029(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1030(.a(G513), .O(gate182inter7));
  inv1  gate1031(.a(G564), .O(gate182inter8));
  nand2 gate1032(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1033(.a(s_69), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1034(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1035(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1036(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate995(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate996(.a(gate185inter0), .b(s_64), .O(gate185inter1));
  and2  gate997(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate998(.a(s_64), .O(gate185inter3));
  inv1  gate999(.a(s_65), .O(gate185inter4));
  nand2 gate1000(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1001(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1002(.a(G570), .O(gate185inter7));
  inv1  gate1003(.a(G571), .O(gate185inter8));
  nand2 gate1004(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1005(.a(s_65), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1006(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1007(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1008(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1051(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1052(.a(gate191inter0), .b(s_72), .O(gate191inter1));
  and2  gate1053(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1054(.a(s_72), .O(gate191inter3));
  inv1  gate1055(.a(s_73), .O(gate191inter4));
  nand2 gate1056(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1057(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1058(.a(G582), .O(gate191inter7));
  inv1  gate1059(.a(G583), .O(gate191inter8));
  nand2 gate1060(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1061(.a(s_73), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1062(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1063(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1064(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate897(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate898(.a(gate203inter0), .b(s_50), .O(gate203inter1));
  and2  gate899(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate900(.a(s_50), .O(gate203inter3));
  inv1  gate901(.a(s_51), .O(gate203inter4));
  nand2 gate902(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate903(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate904(.a(G602), .O(gate203inter7));
  inv1  gate905(.a(G612), .O(gate203inter8));
  nand2 gate906(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate907(.a(s_51), .b(gate203inter3), .O(gate203inter10));
  nor2  gate908(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate909(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate910(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate813(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate814(.a(gate205inter0), .b(s_38), .O(gate205inter1));
  and2  gate815(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate816(.a(s_38), .O(gate205inter3));
  inv1  gate817(.a(s_39), .O(gate205inter4));
  nand2 gate818(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate819(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate820(.a(G622), .O(gate205inter7));
  inv1  gate821(.a(G627), .O(gate205inter8));
  nand2 gate822(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate823(.a(s_39), .b(gate205inter3), .O(gate205inter10));
  nor2  gate824(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate825(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate826(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1107(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1108(.a(gate210inter0), .b(s_80), .O(gate210inter1));
  and2  gate1109(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1110(.a(s_80), .O(gate210inter3));
  inv1  gate1111(.a(s_81), .O(gate210inter4));
  nand2 gate1112(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1113(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1114(.a(G607), .O(gate210inter7));
  inv1  gate1115(.a(G666), .O(gate210inter8));
  nand2 gate1116(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1117(.a(s_81), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1118(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1119(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1120(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate869(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate870(.a(gate229inter0), .b(s_46), .O(gate229inter1));
  and2  gate871(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate872(.a(s_46), .O(gate229inter3));
  inv1  gate873(.a(s_47), .O(gate229inter4));
  nand2 gate874(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate875(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate876(.a(G698), .O(gate229inter7));
  inv1  gate877(.a(G699), .O(gate229inter8));
  nand2 gate878(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate879(.a(s_47), .b(gate229inter3), .O(gate229inter10));
  nor2  gate880(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate881(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate882(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate715(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate716(.a(gate233inter0), .b(s_24), .O(gate233inter1));
  and2  gate717(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate718(.a(s_24), .O(gate233inter3));
  inv1  gate719(.a(s_25), .O(gate233inter4));
  nand2 gate720(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate721(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate722(.a(G242), .O(gate233inter7));
  inv1  gate723(.a(G718), .O(gate233inter8));
  nand2 gate724(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate725(.a(s_25), .b(gate233inter3), .O(gate233inter10));
  nor2  gate726(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate727(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate728(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1121(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1122(.a(gate248inter0), .b(s_82), .O(gate248inter1));
  and2  gate1123(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1124(.a(s_82), .O(gate248inter3));
  inv1  gate1125(.a(s_83), .O(gate248inter4));
  nand2 gate1126(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1127(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1128(.a(G727), .O(gate248inter7));
  inv1  gate1129(.a(G739), .O(gate248inter8));
  nand2 gate1130(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1131(.a(s_83), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1132(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1133(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1134(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate645(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate646(.a(gate250inter0), .b(s_14), .O(gate250inter1));
  and2  gate647(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate648(.a(s_14), .O(gate250inter3));
  inv1  gate649(.a(s_15), .O(gate250inter4));
  nand2 gate650(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate651(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate652(.a(G706), .O(gate250inter7));
  inv1  gate653(.a(G742), .O(gate250inter8));
  nand2 gate654(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate655(.a(s_15), .b(gate250inter3), .O(gate250inter10));
  nor2  gate656(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate657(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate658(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1009(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1010(.a(gate254inter0), .b(s_66), .O(gate254inter1));
  and2  gate1011(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1012(.a(s_66), .O(gate254inter3));
  inv1  gate1013(.a(s_67), .O(gate254inter4));
  nand2 gate1014(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1015(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1016(.a(G712), .O(gate254inter7));
  inv1  gate1017(.a(G748), .O(gate254inter8));
  nand2 gate1018(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1019(.a(s_67), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1020(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1021(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1022(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1163(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1164(.a(gate265inter0), .b(s_88), .O(gate265inter1));
  and2  gate1165(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1166(.a(s_88), .O(gate265inter3));
  inv1  gate1167(.a(s_89), .O(gate265inter4));
  nand2 gate1168(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1169(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1170(.a(G642), .O(gate265inter7));
  inv1  gate1171(.a(G770), .O(gate265inter8));
  nand2 gate1172(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1173(.a(s_89), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1174(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1175(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1176(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1093(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1094(.a(gate269inter0), .b(s_78), .O(gate269inter1));
  and2  gate1095(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1096(.a(s_78), .O(gate269inter3));
  inv1  gate1097(.a(s_79), .O(gate269inter4));
  nand2 gate1098(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1099(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1100(.a(G654), .O(gate269inter7));
  inv1  gate1101(.a(G782), .O(gate269inter8));
  nand2 gate1102(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1103(.a(s_79), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1104(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1105(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1106(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate547(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate548(.a(gate272inter0), .b(s_0), .O(gate272inter1));
  and2  gate549(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate550(.a(s_0), .O(gate272inter3));
  inv1  gate551(.a(s_1), .O(gate272inter4));
  nand2 gate552(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate553(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate554(.a(G663), .O(gate272inter7));
  inv1  gate555(.a(G791), .O(gate272inter8));
  nand2 gate556(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate557(.a(s_1), .b(gate272inter3), .O(gate272inter10));
  nor2  gate558(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate559(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate560(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate911(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate912(.a(gate281inter0), .b(s_52), .O(gate281inter1));
  and2  gate913(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate914(.a(s_52), .O(gate281inter3));
  inv1  gate915(.a(s_53), .O(gate281inter4));
  nand2 gate916(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate917(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate918(.a(G654), .O(gate281inter7));
  inv1  gate919(.a(G806), .O(gate281inter8));
  nand2 gate920(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate921(.a(s_53), .b(gate281inter3), .O(gate281inter10));
  nor2  gate922(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate923(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate924(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1177(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1178(.a(gate292inter0), .b(s_90), .O(gate292inter1));
  and2  gate1179(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1180(.a(s_90), .O(gate292inter3));
  inv1  gate1181(.a(s_91), .O(gate292inter4));
  nand2 gate1182(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1183(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1184(.a(G824), .O(gate292inter7));
  inv1  gate1185(.a(G825), .O(gate292inter8));
  nand2 gate1186(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1187(.a(s_91), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1188(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1189(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1190(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate589(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate590(.a(gate394inter0), .b(s_6), .O(gate394inter1));
  and2  gate591(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate592(.a(s_6), .O(gate394inter3));
  inv1  gate593(.a(s_7), .O(gate394inter4));
  nand2 gate594(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate595(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate596(.a(G8), .O(gate394inter7));
  inv1  gate597(.a(G1057), .O(gate394inter8));
  nand2 gate598(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate599(.a(s_7), .b(gate394inter3), .O(gate394inter10));
  nor2  gate600(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate601(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate602(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate939(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate940(.a(gate397inter0), .b(s_56), .O(gate397inter1));
  and2  gate941(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate942(.a(s_56), .O(gate397inter3));
  inv1  gate943(.a(s_57), .O(gate397inter4));
  nand2 gate944(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate945(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate946(.a(G11), .O(gate397inter7));
  inv1  gate947(.a(G1066), .O(gate397inter8));
  nand2 gate948(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate949(.a(s_57), .b(gate397inter3), .O(gate397inter10));
  nor2  gate950(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate951(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate952(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate687(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate688(.a(gate399inter0), .b(s_20), .O(gate399inter1));
  and2  gate689(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate690(.a(s_20), .O(gate399inter3));
  inv1  gate691(.a(s_21), .O(gate399inter4));
  nand2 gate692(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate693(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate694(.a(G13), .O(gate399inter7));
  inv1  gate695(.a(G1072), .O(gate399inter8));
  nand2 gate696(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate697(.a(s_21), .b(gate399inter3), .O(gate399inter10));
  nor2  gate698(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate699(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate700(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate659(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate660(.a(gate408inter0), .b(s_16), .O(gate408inter1));
  and2  gate661(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate662(.a(s_16), .O(gate408inter3));
  inv1  gate663(.a(s_17), .O(gate408inter4));
  nand2 gate664(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate665(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate666(.a(G22), .O(gate408inter7));
  inv1  gate667(.a(G1099), .O(gate408inter8));
  nand2 gate668(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate669(.a(s_17), .b(gate408inter3), .O(gate408inter10));
  nor2  gate670(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate671(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate672(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate967(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate968(.a(gate419inter0), .b(s_60), .O(gate419inter1));
  and2  gate969(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate970(.a(s_60), .O(gate419inter3));
  inv1  gate971(.a(s_61), .O(gate419inter4));
  nand2 gate972(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate973(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate974(.a(G1), .O(gate419inter7));
  inv1  gate975(.a(G1132), .O(gate419inter8));
  nand2 gate976(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate977(.a(s_61), .b(gate419inter3), .O(gate419inter10));
  nor2  gate978(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate979(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate980(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate729(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate730(.a(gate455inter0), .b(s_26), .O(gate455inter1));
  and2  gate731(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate732(.a(s_26), .O(gate455inter3));
  inv1  gate733(.a(s_27), .O(gate455inter4));
  nand2 gate734(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate735(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate736(.a(G19), .O(gate455inter7));
  inv1  gate737(.a(G1186), .O(gate455inter8));
  nand2 gate738(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate739(.a(s_27), .b(gate455inter3), .O(gate455inter10));
  nor2  gate740(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate741(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate742(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate855(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate856(.a(gate461inter0), .b(s_44), .O(gate461inter1));
  and2  gate857(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate858(.a(s_44), .O(gate461inter3));
  inv1  gate859(.a(s_45), .O(gate461inter4));
  nand2 gate860(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate861(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate862(.a(G22), .O(gate461inter7));
  inv1  gate863(.a(G1195), .O(gate461inter8));
  nand2 gate864(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate865(.a(s_45), .b(gate461inter3), .O(gate461inter10));
  nor2  gate866(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate867(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate868(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate757(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate758(.a(gate462inter0), .b(s_30), .O(gate462inter1));
  and2  gate759(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate760(.a(s_30), .O(gate462inter3));
  inv1  gate761(.a(s_31), .O(gate462inter4));
  nand2 gate762(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate763(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate764(.a(G1099), .O(gate462inter7));
  inv1  gate765(.a(G1195), .O(gate462inter8));
  nand2 gate766(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate767(.a(s_31), .b(gate462inter3), .O(gate462inter10));
  nor2  gate768(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate769(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate770(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate883(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate884(.a(gate464inter0), .b(s_48), .O(gate464inter1));
  and2  gate885(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate886(.a(s_48), .O(gate464inter3));
  inv1  gate887(.a(s_49), .O(gate464inter4));
  nand2 gate888(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate889(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate890(.a(G1102), .O(gate464inter7));
  inv1  gate891(.a(G1198), .O(gate464inter8));
  nand2 gate892(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate893(.a(s_49), .b(gate464inter3), .O(gate464inter10));
  nor2  gate894(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate895(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate896(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate631(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate632(.a(gate478inter0), .b(s_12), .O(gate478inter1));
  and2  gate633(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate634(.a(s_12), .O(gate478inter3));
  inv1  gate635(.a(s_13), .O(gate478inter4));
  nand2 gate636(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate637(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate638(.a(G1123), .O(gate478inter7));
  inv1  gate639(.a(G1219), .O(gate478inter8));
  nand2 gate640(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate641(.a(s_13), .b(gate478inter3), .O(gate478inter10));
  nor2  gate642(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate643(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate644(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate617(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate618(.a(gate491inter0), .b(s_10), .O(gate491inter1));
  and2  gate619(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate620(.a(s_10), .O(gate491inter3));
  inv1  gate621(.a(s_11), .O(gate491inter4));
  nand2 gate622(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate623(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate624(.a(G1244), .O(gate491inter7));
  inv1  gate625(.a(G1245), .O(gate491inter8));
  nand2 gate626(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate627(.a(s_11), .b(gate491inter3), .O(gate491inter10));
  nor2  gate628(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate629(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate630(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate827(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate828(.a(gate494inter0), .b(s_40), .O(gate494inter1));
  and2  gate829(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate830(.a(s_40), .O(gate494inter3));
  inv1  gate831(.a(s_41), .O(gate494inter4));
  nand2 gate832(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate833(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate834(.a(G1250), .O(gate494inter7));
  inv1  gate835(.a(G1251), .O(gate494inter8));
  nand2 gate836(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate837(.a(s_41), .b(gate494inter3), .O(gate494inter10));
  nor2  gate838(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate839(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate840(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1135(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1136(.a(gate495inter0), .b(s_84), .O(gate495inter1));
  and2  gate1137(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1138(.a(s_84), .O(gate495inter3));
  inv1  gate1139(.a(s_85), .O(gate495inter4));
  nand2 gate1140(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1141(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1142(.a(G1252), .O(gate495inter7));
  inv1  gate1143(.a(G1253), .O(gate495inter8));
  nand2 gate1144(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1145(.a(s_85), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1146(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1147(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1148(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate561(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate562(.a(gate497inter0), .b(s_2), .O(gate497inter1));
  and2  gate563(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate564(.a(s_2), .O(gate497inter3));
  inv1  gate565(.a(s_3), .O(gate497inter4));
  nand2 gate566(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate567(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate568(.a(G1256), .O(gate497inter7));
  inv1  gate569(.a(G1257), .O(gate497inter8));
  nand2 gate570(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate571(.a(s_3), .b(gate497inter3), .O(gate497inter10));
  nor2  gate572(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate573(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate574(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate981(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate982(.a(gate511inter0), .b(s_62), .O(gate511inter1));
  and2  gate983(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate984(.a(s_62), .O(gate511inter3));
  inv1  gate985(.a(s_63), .O(gate511inter4));
  nand2 gate986(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate987(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate988(.a(G1284), .O(gate511inter7));
  inv1  gate989(.a(G1285), .O(gate511inter8));
  nand2 gate990(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate991(.a(s_63), .b(gate511inter3), .O(gate511inter10));
  nor2  gate992(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate993(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate994(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule