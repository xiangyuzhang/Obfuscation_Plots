module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1681(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1682(.a(gate10inter0), .b(s_162), .O(gate10inter1));
  and2  gate1683(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1684(.a(s_162), .O(gate10inter3));
  inv1  gate1685(.a(s_163), .O(gate10inter4));
  nand2 gate1686(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1687(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1688(.a(G3), .O(gate10inter7));
  inv1  gate1689(.a(G4), .O(gate10inter8));
  nand2 gate1690(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1691(.a(s_163), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1692(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1693(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1694(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2073(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2074(.a(gate12inter0), .b(s_218), .O(gate12inter1));
  and2  gate2075(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2076(.a(s_218), .O(gate12inter3));
  inv1  gate2077(.a(s_219), .O(gate12inter4));
  nand2 gate2078(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2079(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2080(.a(G7), .O(gate12inter7));
  inv1  gate2081(.a(G8), .O(gate12inter8));
  nand2 gate2082(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2083(.a(s_219), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2084(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2085(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2086(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1037(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1038(.a(gate15inter0), .b(s_70), .O(gate15inter1));
  and2  gate1039(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1040(.a(s_70), .O(gate15inter3));
  inv1  gate1041(.a(s_71), .O(gate15inter4));
  nand2 gate1042(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1043(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1044(.a(G13), .O(gate15inter7));
  inv1  gate1045(.a(G14), .O(gate15inter8));
  nand2 gate1046(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1047(.a(s_71), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1048(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1049(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1050(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate869(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate870(.a(gate16inter0), .b(s_46), .O(gate16inter1));
  and2  gate871(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate872(.a(s_46), .O(gate16inter3));
  inv1  gate873(.a(s_47), .O(gate16inter4));
  nand2 gate874(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate875(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate876(.a(G15), .O(gate16inter7));
  inv1  gate877(.a(G16), .O(gate16inter8));
  nand2 gate878(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate879(.a(s_47), .b(gate16inter3), .O(gate16inter10));
  nor2  gate880(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate881(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate882(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2003(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2004(.a(gate17inter0), .b(s_208), .O(gate17inter1));
  and2  gate2005(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2006(.a(s_208), .O(gate17inter3));
  inv1  gate2007(.a(s_209), .O(gate17inter4));
  nand2 gate2008(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2009(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2010(.a(G17), .O(gate17inter7));
  inv1  gate2011(.a(G18), .O(gate17inter8));
  nand2 gate2012(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2013(.a(s_209), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2014(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2015(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2016(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1163(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1164(.a(gate20inter0), .b(s_88), .O(gate20inter1));
  and2  gate1165(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1166(.a(s_88), .O(gate20inter3));
  inv1  gate1167(.a(s_89), .O(gate20inter4));
  nand2 gate1168(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1169(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1170(.a(G23), .O(gate20inter7));
  inv1  gate1171(.a(G24), .O(gate20inter8));
  nand2 gate1172(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1173(.a(s_89), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1174(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1175(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1176(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1751(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1752(.a(gate21inter0), .b(s_172), .O(gate21inter1));
  and2  gate1753(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1754(.a(s_172), .O(gate21inter3));
  inv1  gate1755(.a(s_173), .O(gate21inter4));
  nand2 gate1756(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1757(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1758(.a(G25), .O(gate21inter7));
  inv1  gate1759(.a(G26), .O(gate21inter8));
  nand2 gate1760(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1761(.a(s_173), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1762(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1763(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1764(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1905(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1906(.a(gate22inter0), .b(s_194), .O(gate22inter1));
  and2  gate1907(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1908(.a(s_194), .O(gate22inter3));
  inv1  gate1909(.a(s_195), .O(gate22inter4));
  nand2 gate1910(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1911(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1912(.a(G27), .O(gate22inter7));
  inv1  gate1913(.a(G28), .O(gate22inter8));
  nand2 gate1914(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1915(.a(s_195), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1916(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1917(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1918(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1989(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1990(.a(gate25inter0), .b(s_206), .O(gate25inter1));
  and2  gate1991(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1992(.a(s_206), .O(gate25inter3));
  inv1  gate1993(.a(s_207), .O(gate25inter4));
  nand2 gate1994(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1995(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1996(.a(G1), .O(gate25inter7));
  inv1  gate1997(.a(G5), .O(gate25inter8));
  nand2 gate1998(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1999(.a(s_207), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2000(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2001(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2002(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate715(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate716(.a(gate27inter0), .b(s_24), .O(gate27inter1));
  and2  gate717(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate718(.a(s_24), .O(gate27inter3));
  inv1  gate719(.a(s_25), .O(gate27inter4));
  nand2 gate720(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate721(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate722(.a(G2), .O(gate27inter7));
  inv1  gate723(.a(G6), .O(gate27inter8));
  nand2 gate724(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate725(.a(s_25), .b(gate27inter3), .O(gate27inter10));
  nor2  gate726(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate727(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate728(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate575(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate576(.a(gate28inter0), .b(s_4), .O(gate28inter1));
  and2  gate577(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate578(.a(s_4), .O(gate28inter3));
  inv1  gate579(.a(s_5), .O(gate28inter4));
  nand2 gate580(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate581(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate582(.a(G10), .O(gate28inter7));
  inv1  gate583(.a(G14), .O(gate28inter8));
  nand2 gate584(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate585(.a(s_5), .b(gate28inter3), .O(gate28inter10));
  nor2  gate586(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate587(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate588(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1219(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1220(.a(gate32inter0), .b(s_96), .O(gate32inter1));
  and2  gate1221(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1222(.a(s_96), .O(gate32inter3));
  inv1  gate1223(.a(s_97), .O(gate32inter4));
  nand2 gate1224(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1225(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1226(.a(G12), .O(gate32inter7));
  inv1  gate1227(.a(G16), .O(gate32inter8));
  nand2 gate1228(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1229(.a(s_97), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1230(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1231(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1232(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1737(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1738(.a(gate33inter0), .b(s_170), .O(gate33inter1));
  and2  gate1739(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1740(.a(s_170), .O(gate33inter3));
  inv1  gate1741(.a(s_171), .O(gate33inter4));
  nand2 gate1742(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1743(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1744(.a(G17), .O(gate33inter7));
  inv1  gate1745(.a(G21), .O(gate33inter8));
  nand2 gate1746(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1747(.a(s_171), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1748(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1749(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1750(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2171(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2172(.a(gate35inter0), .b(s_232), .O(gate35inter1));
  and2  gate2173(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2174(.a(s_232), .O(gate35inter3));
  inv1  gate2175(.a(s_233), .O(gate35inter4));
  nand2 gate2176(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2177(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2178(.a(G18), .O(gate35inter7));
  inv1  gate2179(.a(G22), .O(gate35inter8));
  nand2 gate2180(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2181(.a(s_233), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2182(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2183(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2184(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate757(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate758(.a(gate36inter0), .b(s_30), .O(gate36inter1));
  and2  gate759(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate760(.a(s_30), .O(gate36inter3));
  inv1  gate761(.a(s_31), .O(gate36inter4));
  nand2 gate762(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate763(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate764(.a(G26), .O(gate36inter7));
  inv1  gate765(.a(G30), .O(gate36inter8));
  nand2 gate766(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate767(.a(s_31), .b(gate36inter3), .O(gate36inter10));
  nor2  gate768(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate769(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate770(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1723(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1724(.a(gate39inter0), .b(s_168), .O(gate39inter1));
  and2  gate1725(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1726(.a(s_168), .O(gate39inter3));
  inv1  gate1727(.a(s_169), .O(gate39inter4));
  nand2 gate1728(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1729(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1730(.a(G20), .O(gate39inter7));
  inv1  gate1731(.a(G24), .O(gate39inter8));
  nand2 gate1732(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1733(.a(s_169), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1734(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1735(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1736(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2101(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2102(.a(gate44inter0), .b(s_222), .O(gate44inter1));
  and2  gate2103(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2104(.a(s_222), .O(gate44inter3));
  inv1  gate2105(.a(s_223), .O(gate44inter4));
  nand2 gate2106(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2107(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2108(.a(G4), .O(gate44inter7));
  inv1  gate2109(.a(G269), .O(gate44inter8));
  nand2 gate2110(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2111(.a(s_223), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2112(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2113(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2114(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate855(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate856(.a(gate45inter0), .b(s_44), .O(gate45inter1));
  and2  gate857(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate858(.a(s_44), .O(gate45inter3));
  inv1  gate859(.a(s_45), .O(gate45inter4));
  nand2 gate860(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate861(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate862(.a(G5), .O(gate45inter7));
  inv1  gate863(.a(G272), .O(gate45inter8));
  nand2 gate864(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate865(.a(s_45), .b(gate45inter3), .O(gate45inter10));
  nor2  gate866(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate867(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate868(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1191(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1192(.a(gate52inter0), .b(s_92), .O(gate52inter1));
  and2  gate1193(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1194(.a(s_92), .O(gate52inter3));
  inv1  gate1195(.a(s_93), .O(gate52inter4));
  nand2 gate1196(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1197(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1198(.a(G12), .O(gate52inter7));
  inv1  gate1199(.a(G281), .O(gate52inter8));
  nand2 gate1200(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1201(.a(s_93), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1202(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1203(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1204(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2045(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2046(.a(gate55inter0), .b(s_214), .O(gate55inter1));
  and2  gate2047(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2048(.a(s_214), .O(gate55inter3));
  inv1  gate2049(.a(s_215), .O(gate55inter4));
  nand2 gate2050(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2051(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2052(.a(G15), .O(gate55inter7));
  inv1  gate2053(.a(G287), .O(gate55inter8));
  nand2 gate2054(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2055(.a(s_215), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2056(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2057(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2058(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1569(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1570(.a(gate56inter0), .b(s_146), .O(gate56inter1));
  and2  gate1571(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1572(.a(s_146), .O(gate56inter3));
  inv1  gate1573(.a(s_147), .O(gate56inter4));
  nand2 gate1574(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1575(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1576(.a(G16), .O(gate56inter7));
  inv1  gate1577(.a(G287), .O(gate56inter8));
  nand2 gate1578(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1579(.a(s_147), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1580(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1581(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1582(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate589(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate590(.a(gate61inter0), .b(s_6), .O(gate61inter1));
  and2  gate591(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate592(.a(s_6), .O(gate61inter3));
  inv1  gate593(.a(s_7), .O(gate61inter4));
  nand2 gate594(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate595(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate596(.a(G21), .O(gate61inter7));
  inv1  gate597(.a(G296), .O(gate61inter8));
  nand2 gate598(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate599(.a(s_7), .b(gate61inter3), .O(gate61inter10));
  nor2  gate600(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate601(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate602(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2423(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2424(.a(gate62inter0), .b(s_268), .O(gate62inter1));
  and2  gate2425(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2426(.a(s_268), .O(gate62inter3));
  inv1  gate2427(.a(s_269), .O(gate62inter4));
  nand2 gate2428(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2429(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2430(.a(G22), .O(gate62inter7));
  inv1  gate2431(.a(G296), .O(gate62inter8));
  nand2 gate2432(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2433(.a(s_269), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2434(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2435(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2436(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate561(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate562(.a(gate68inter0), .b(s_2), .O(gate68inter1));
  and2  gate563(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate564(.a(s_2), .O(gate68inter3));
  inv1  gate565(.a(s_3), .O(gate68inter4));
  nand2 gate566(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate567(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate568(.a(G28), .O(gate68inter7));
  inv1  gate569(.a(G305), .O(gate68inter8));
  nand2 gate570(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate571(.a(s_3), .b(gate68inter3), .O(gate68inter10));
  nor2  gate572(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate573(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate574(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate1205(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1206(.a(gate69inter0), .b(s_94), .O(gate69inter1));
  and2  gate1207(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1208(.a(s_94), .O(gate69inter3));
  inv1  gate1209(.a(s_95), .O(gate69inter4));
  nand2 gate1210(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1211(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1212(.a(G29), .O(gate69inter7));
  inv1  gate1213(.a(G308), .O(gate69inter8));
  nand2 gate1214(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1215(.a(s_95), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1216(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1217(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1218(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1541(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1542(.a(gate72inter0), .b(s_142), .O(gate72inter1));
  and2  gate1543(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1544(.a(s_142), .O(gate72inter3));
  inv1  gate1545(.a(s_143), .O(gate72inter4));
  nand2 gate1546(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1547(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1548(.a(G32), .O(gate72inter7));
  inv1  gate1549(.a(G311), .O(gate72inter8));
  nand2 gate1550(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1551(.a(s_143), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1552(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1553(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1554(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1919(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1920(.a(gate73inter0), .b(s_196), .O(gate73inter1));
  and2  gate1921(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1922(.a(s_196), .O(gate73inter3));
  inv1  gate1923(.a(s_197), .O(gate73inter4));
  nand2 gate1924(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1925(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1926(.a(G1), .O(gate73inter7));
  inv1  gate1927(.a(G314), .O(gate73inter8));
  nand2 gate1928(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1929(.a(s_197), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1930(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1931(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1932(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2087(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2088(.a(gate78inter0), .b(s_220), .O(gate78inter1));
  and2  gate2089(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2090(.a(s_220), .O(gate78inter3));
  inv1  gate2091(.a(s_221), .O(gate78inter4));
  nand2 gate2092(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2093(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2094(.a(G6), .O(gate78inter7));
  inv1  gate2095(.a(G320), .O(gate78inter8));
  nand2 gate2096(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2097(.a(s_221), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2098(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2099(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2100(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2227(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2228(.a(gate82inter0), .b(s_240), .O(gate82inter1));
  and2  gate2229(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2230(.a(s_240), .O(gate82inter3));
  inv1  gate2231(.a(s_241), .O(gate82inter4));
  nand2 gate2232(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2233(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2234(.a(G7), .O(gate82inter7));
  inv1  gate2235(.a(G326), .O(gate82inter8));
  nand2 gate2236(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2237(.a(s_241), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2238(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2239(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2240(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate925(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate926(.a(gate91inter0), .b(s_54), .O(gate91inter1));
  and2  gate927(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate928(.a(s_54), .O(gate91inter3));
  inv1  gate929(.a(s_55), .O(gate91inter4));
  nand2 gate930(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate931(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate932(.a(G25), .O(gate91inter7));
  inv1  gate933(.a(G341), .O(gate91inter8));
  nand2 gate934(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate935(.a(s_55), .b(gate91inter3), .O(gate91inter10));
  nor2  gate936(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate937(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate938(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate673(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate674(.a(gate96inter0), .b(s_18), .O(gate96inter1));
  and2  gate675(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate676(.a(s_18), .O(gate96inter3));
  inv1  gate677(.a(s_19), .O(gate96inter4));
  nand2 gate678(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate679(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate680(.a(G30), .O(gate96inter7));
  inv1  gate681(.a(G347), .O(gate96inter8));
  nand2 gate682(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate683(.a(s_19), .b(gate96inter3), .O(gate96inter10));
  nor2  gate684(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate685(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate686(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2493(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2494(.a(gate97inter0), .b(s_278), .O(gate97inter1));
  and2  gate2495(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2496(.a(s_278), .O(gate97inter3));
  inv1  gate2497(.a(s_279), .O(gate97inter4));
  nand2 gate2498(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2499(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2500(.a(G19), .O(gate97inter7));
  inv1  gate2501(.a(G350), .O(gate97inter8));
  nand2 gate2502(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2503(.a(s_279), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2504(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2505(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2506(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1443(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1444(.a(gate99inter0), .b(s_128), .O(gate99inter1));
  and2  gate1445(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1446(.a(s_128), .O(gate99inter3));
  inv1  gate1447(.a(s_129), .O(gate99inter4));
  nand2 gate1448(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1449(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1450(.a(G27), .O(gate99inter7));
  inv1  gate1451(.a(G353), .O(gate99inter8));
  nand2 gate1452(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1453(.a(s_129), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1454(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1455(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1456(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate981(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate982(.a(gate109inter0), .b(s_62), .O(gate109inter1));
  and2  gate983(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate984(.a(s_62), .O(gate109inter3));
  inv1  gate985(.a(s_63), .O(gate109inter4));
  nand2 gate986(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate987(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate988(.a(G370), .O(gate109inter7));
  inv1  gate989(.a(G371), .O(gate109inter8));
  nand2 gate990(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate991(.a(s_63), .b(gate109inter3), .O(gate109inter10));
  nor2  gate992(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate993(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate994(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1303(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1304(.a(gate112inter0), .b(s_108), .O(gate112inter1));
  and2  gate1305(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1306(.a(s_108), .O(gate112inter3));
  inv1  gate1307(.a(s_109), .O(gate112inter4));
  nand2 gate1308(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1309(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1310(.a(G376), .O(gate112inter7));
  inv1  gate1311(.a(G377), .O(gate112inter8));
  nand2 gate1312(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1313(.a(s_109), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1314(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1315(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1316(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1975(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1976(.a(gate113inter0), .b(s_204), .O(gate113inter1));
  and2  gate1977(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1978(.a(s_204), .O(gate113inter3));
  inv1  gate1979(.a(s_205), .O(gate113inter4));
  nand2 gate1980(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1981(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1982(.a(G378), .O(gate113inter7));
  inv1  gate1983(.a(G379), .O(gate113inter8));
  nand2 gate1984(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1985(.a(s_205), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1986(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1987(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1988(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1065(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1066(.a(gate115inter0), .b(s_74), .O(gate115inter1));
  and2  gate1067(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1068(.a(s_74), .O(gate115inter3));
  inv1  gate1069(.a(s_75), .O(gate115inter4));
  nand2 gate1070(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1071(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1072(.a(G382), .O(gate115inter7));
  inv1  gate1073(.a(G383), .O(gate115inter8));
  nand2 gate1074(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1075(.a(s_75), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1076(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1077(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1078(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1709(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1710(.a(gate116inter0), .b(s_166), .O(gate116inter1));
  and2  gate1711(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1712(.a(s_166), .O(gate116inter3));
  inv1  gate1713(.a(s_167), .O(gate116inter4));
  nand2 gate1714(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1715(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1716(.a(G384), .O(gate116inter7));
  inv1  gate1717(.a(G385), .O(gate116inter8));
  nand2 gate1718(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1719(.a(s_167), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1720(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1721(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1722(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate2143(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2144(.a(gate117inter0), .b(s_228), .O(gate117inter1));
  and2  gate2145(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2146(.a(s_228), .O(gate117inter3));
  inv1  gate2147(.a(s_229), .O(gate117inter4));
  nand2 gate2148(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2149(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2150(.a(G386), .O(gate117inter7));
  inv1  gate2151(.a(G387), .O(gate117inter8));
  nand2 gate2152(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2153(.a(s_229), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2154(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2155(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2156(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate827(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate828(.a(gate122inter0), .b(s_40), .O(gate122inter1));
  and2  gate829(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate830(.a(s_40), .O(gate122inter3));
  inv1  gate831(.a(s_41), .O(gate122inter4));
  nand2 gate832(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate833(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate834(.a(G396), .O(gate122inter7));
  inv1  gate835(.a(G397), .O(gate122inter8));
  nand2 gate836(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate837(.a(s_41), .b(gate122inter3), .O(gate122inter10));
  nor2  gate838(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate839(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate840(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1373(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1374(.a(gate124inter0), .b(s_118), .O(gate124inter1));
  and2  gate1375(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1376(.a(s_118), .O(gate124inter3));
  inv1  gate1377(.a(s_119), .O(gate124inter4));
  nand2 gate1378(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1379(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1380(.a(G400), .O(gate124inter7));
  inv1  gate1381(.a(G401), .O(gate124inter8));
  nand2 gate1382(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1383(.a(s_119), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1384(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1385(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1386(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1149(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1150(.a(gate132inter0), .b(s_86), .O(gate132inter1));
  and2  gate1151(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1152(.a(s_86), .O(gate132inter3));
  inv1  gate1153(.a(s_87), .O(gate132inter4));
  nand2 gate1154(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1155(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1156(.a(G416), .O(gate132inter7));
  inv1  gate1157(.a(G417), .O(gate132inter8));
  nand2 gate1158(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1159(.a(s_87), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1160(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1161(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1162(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1765(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1766(.a(gate134inter0), .b(s_174), .O(gate134inter1));
  and2  gate1767(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1768(.a(s_174), .O(gate134inter3));
  inv1  gate1769(.a(s_175), .O(gate134inter4));
  nand2 gate1770(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1771(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1772(.a(G420), .O(gate134inter7));
  inv1  gate1773(.a(G421), .O(gate134inter8));
  nand2 gate1774(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1775(.a(s_175), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1776(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1777(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1778(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2017(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2018(.a(gate137inter0), .b(s_210), .O(gate137inter1));
  and2  gate2019(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2020(.a(s_210), .O(gate137inter3));
  inv1  gate2021(.a(s_211), .O(gate137inter4));
  nand2 gate2022(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2023(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2024(.a(G426), .O(gate137inter7));
  inv1  gate2025(.a(G429), .O(gate137inter8));
  nand2 gate2026(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2027(.a(s_211), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2028(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2029(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2030(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate967(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate968(.a(gate140inter0), .b(s_60), .O(gate140inter1));
  and2  gate969(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate970(.a(s_60), .O(gate140inter3));
  inv1  gate971(.a(s_61), .O(gate140inter4));
  nand2 gate972(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate973(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate974(.a(G444), .O(gate140inter7));
  inv1  gate975(.a(G447), .O(gate140inter8));
  nand2 gate976(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate977(.a(s_61), .b(gate140inter3), .O(gate140inter10));
  nor2  gate978(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate979(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate980(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1821(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1822(.a(gate142inter0), .b(s_182), .O(gate142inter1));
  and2  gate1823(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1824(.a(s_182), .O(gate142inter3));
  inv1  gate1825(.a(s_183), .O(gate142inter4));
  nand2 gate1826(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1827(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1828(.a(G456), .O(gate142inter7));
  inv1  gate1829(.a(G459), .O(gate142inter8));
  nand2 gate1830(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1831(.a(s_183), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1832(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1833(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1834(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1387(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1388(.a(gate146inter0), .b(s_120), .O(gate146inter1));
  and2  gate1389(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1390(.a(s_120), .O(gate146inter3));
  inv1  gate1391(.a(s_121), .O(gate146inter4));
  nand2 gate1392(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1393(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1394(.a(G480), .O(gate146inter7));
  inv1  gate1395(.a(G483), .O(gate146inter8));
  nand2 gate1396(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1397(.a(s_121), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1398(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1399(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1400(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate687(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate688(.a(gate147inter0), .b(s_20), .O(gate147inter1));
  and2  gate689(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate690(.a(s_20), .O(gate147inter3));
  inv1  gate691(.a(s_21), .O(gate147inter4));
  nand2 gate692(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate693(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate694(.a(G486), .O(gate147inter7));
  inv1  gate695(.a(G489), .O(gate147inter8));
  nand2 gate696(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate697(.a(s_21), .b(gate147inter3), .O(gate147inter10));
  nor2  gate698(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate699(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate700(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1429(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1430(.a(gate148inter0), .b(s_126), .O(gate148inter1));
  and2  gate1431(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1432(.a(s_126), .O(gate148inter3));
  inv1  gate1433(.a(s_127), .O(gate148inter4));
  nand2 gate1434(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1435(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1436(.a(G492), .O(gate148inter7));
  inv1  gate1437(.a(G495), .O(gate148inter8));
  nand2 gate1438(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1439(.a(s_127), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1440(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1441(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1442(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate645(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate646(.a(gate151inter0), .b(s_14), .O(gate151inter1));
  and2  gate647(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate648(.a(s_14), .O(gate151inter3));
  inv1  gate649(.a(s_15), .O(gate151inter4));
  nand2 gate650(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate651(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate652(.a(G510), .O(gate151inter7));
  inv1  gate653(.a(G513), .O(gate151inter8));
  nand2 gate654(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate655(.a(s_15), .b(gate151inter3), .O(gate151inter10));
  nor2  gate656(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate657(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate658(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2199(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2200(.a(gate152inter0), .b(s_236), .O(gate152inter1));
  and2  gate2201(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2202(.a(s_236), .O(gate152inter3));
  inv1  gate2203(.a(s_237), .O(gate152inter4));
  nand2 gate2204(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2205(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2206(.a(G516), .O(gate152inter7));
  inv1  gate2207(.a(G519), .O(gate152inter8));
  nand2 gate2208(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2209(.a(s_237), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2210(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2211(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2212(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate2185(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2186(.a(gate163inter0), .b(s_234), .O(gate163inter1));
  and2  gate2187(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2188(.a(s_234), .O(gate163inter3));
  inv1  gate2189(.a(s_235), .O(gate163inter4));
  nand2 gate2190(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2191(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2192(.a(G456), .O(gate163inter7));
  inv1  gate2193(.a(G537), .O(gate163inter8));
  nand2 gate2194(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2195(.a(s_235), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2196(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2197(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2198(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1877(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1878(.a(gate164inter0), .b(s_190), .O(gate164inter1));
  and2  gate1879(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1880(.a(s_190), .O(gate164inter3));
  inv1  gate1881(.a(s_191), .O(gate164inter4));
  nand2 gate1882(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1883(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1884(.a(G459), .O(gate164inter7));
  inv1  gate1885(.a(G537), .O(gate164inter8));
  nand2 gate1886(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1887(.a(s_191), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1888(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1889(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1890(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate2325(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2326(.a(gate165inter0), .b(s_254), .O(gate165inter1));
  and2  gate2327(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2328(.a(s_254), .O(gate165inter3));
  inv1  gate2329(.a(s_255), .O(gate165inter4));
  nand2 gate2330(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2331(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2332(.a(G462), .O(gate165inter7));
  inv1  gate2333(.a(G540), .O(gate165inter8));
  nand2 gate2334(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2335(.a(s_255), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2336(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2337(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2338(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2465(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2466(.a(gate173inter0), .b(s_274), .O(gate173inter1));
  and2  gate2467(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2468(.a(s_274), .O(gate173inter3));
  inv1  gate2469(.a(s_275), .O(gate173inter4));
  nand2 gate2470(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2471(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2472(.a(G486), .O(gate173inter7));
  inv1  gate2473(.a(G552), .O(gate173inter8));
  nand2 gate2474(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2475(.a(s_275), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2476(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2477(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2478(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2255(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2256(.a(gate174inter0), .b(s_244), .O(gate174inter1));
  and2  gate2257(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2258(.a(s_244), .O(gate174inter3));
  inv1  gate2259(.a(s_245), .O(gate174inter4));
  nand2 gate2260(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2261(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2262(.a(G489), .O(gate174inter7));
  inv1  gate2263(.a(G552), .O(gate174inter8));
  nand2 gate2264(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2265(.a(s_245), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2266(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2267(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2268(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate2395(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2396(.a(gate177inter0), .b(s_264), .O(gate177inter1));
  and2  gate2397(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2398(.a(s_264), .O(gate177inter3));
  inv1  gate2399(.a(s_265), .O(gate177inter4));
  nand2 gate2400(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2401(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2402(.a(G498), .O(gate177inter7));
  inv1  gate2403(.a(G558), .O(gate177inter8));
  nand2 gate2404(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2405(.a(s_265), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2406(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2407(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2408(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2241(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2242(.a(gate181inter0), .b(s_242), .O(gate181inter1));
  and2  gate2243(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2244(.a(s_242), .O(gate181inter3));
  inv1  gate2245(.a(s_243), .O(gate181inter4));
  nand2 gate2246(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2247(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2248(.a(G510), .O(gate181inter7));
  inv1  gate2249(.a(G564), .O(gate181inter8));
  nand2 gate2250(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2251(.a(s_243), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2252(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2253(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2254(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1079(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1080(.a(gate182inter0), .b(s_76), .O(gate182inter1));
  and2  gate1081(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1082(.a(s_76), .O(gate182inter3));
  inv1  gate1083(.a(s_77), .O(gate182inter4));
  nand2 gate1084(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1085(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1086(.a(G513), .O(gate182inter7));
  inv1  gate1087(.a(G564), .O(gate182inter8));
  nand2 gate1088(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1089(.a(s_77), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1090(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1091(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1092(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2507(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2508(.a(gate184inter0), .b(s_280), .O(gate184inter1));
  and2  gate2509(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2510(.a(s_280), .O(gate184inter3));
  inv1  gate2511(.a(s_281), .O(gate184inter4));
  nand2 gate2512(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2513(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2514(.a(G519), .O(gate184inter7));
  inv1  gate2515(.a(G567), .O(gate184inter8));
  nand2 gate2516(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2517(.a(s_281), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2518(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2519(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2520(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate631(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate632(.a(gate186inter0), .b(s_12), .O(gate186inter1));
  and2  gate633(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate634(.a(s_12), .O(gate186inter3));
  inv1  gate635(.a(s_13), .O(gate186inter4));
  nand2 gate636(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate637(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate638(.a(G572), .O(gate186inter7));
  inv1  gate639(.a(G573), .O(gate186inter8));
  nand2 gate640(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate641(.a(s_13), .b(gate186inter3), .O(gate186inter10));
  nor2  gate642(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate643(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate644(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1835(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1836(.a(gate192inter0), .b(s_184), .O(gate192inter1));
  and2  gate1837(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1838(.a(s_184), .O(gate192inter3));
  inv1  gate1839(.a(s_185), .O(gate192inter4));
  nand2 gate1840(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1841(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1842(.a(G584), .O(gate192inter7));
  inv1  gate1843(.a(G585), .O(gate192inter8));
  nand2 gate1844(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1845(.a(s_185), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1846(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1847(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1848(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1653(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1654(.a(gate194inter0), .b(s_158), .O(gate194inter1));
  and2  gate1655(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1656(.a(s_158), .O(gate194inter3));
  inv1  gate1657(.a(s_159), .O(gate194inter4));
  nand2 gate1658(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1659(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1660(.a(G588), .O(gate194inter7));
  inv1  gate1661(.a(G589), .O(gate194inter8));
  nand2 gate1662(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1663(.a(s_159), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1664(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1665(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1666(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1331(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1332(.a(gate198inter0), .b(s_112), .O(gate198inter1));
  and2  gate1333(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1334(.a(s_112), .O(gate198inter3));
  inv1  gate1335(.a(s_113), .O(gate198inter4));
  nand2 gate1336(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1337(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1338(.a(G596), .O(gate198inter7));
  inv1  gate1339(.a(G597), .O(gate198inter8));
  nand2 gate1340(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1341(.a(s_113), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1342(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1343(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1344(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1583(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1584(.a(gate201inter0), .b(s_148), .O(gate201inter1));
  and2  gate1585(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1586(.a(s_148), .O(gate201inter3));
  inv1  gate1587(.a(s_149), .O(gate201inter4));
  nand2 gate1588(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1589(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1590(.a(G602), .O(gate201inter7));
  inv1  gate1591(.a(G607), .O(gate201inter8));
  nand2 gate1592(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1593(.a(s_149), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1594(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1595(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1596(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2059(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2060(.a(gate207inter0), .b(s_216), .O(gate207inter1));
  and2  gate2061(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2062(.a(s_216), .O(gate207inter3));
  inv1  gate2063(.a(s_217), .O(gate207inter4));
  nand2 gate2064(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2065(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2066(.a(G622), .O(gate207inter7));
  inv1  gate2067(.a(G632), .O(gate207inter8));
  nand2 gate2068(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2069(.a(s_217), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2070(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2071(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2072(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate953(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate954(.a(gate208inter0), .b(s_58), .O(gate208inter1));
  and2  gate955(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate956(.a(s_58), .O(gate208inter3));
  inv1  gate957(.a(s_59), .O(gate208inter4));
  nand2 gate958(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate959(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate960(.a(G627), .O(gate208inter7));
  inv1  gate961(.a(G637), .O(gate208inter8));
  nand2 gate962(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate963(.a(s_59), .b(gate208inter3), .O(gate208inter10));
  nor2  gate964(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate965(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate966(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1947(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1948(.a(gate212inter0), .b(s_200), .O(gate212inter1));
  and2  gate1949(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1950(.a(s_200), .O(gate212inter3));
  inv1  gate1951(.a(s_201), .O(gate212inter4));
  nand2 gate1952(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1953(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1954(.a(G617), .O(gate212inter7));
  inv1  gate1955(.a(G669), .O(gate212inter8));
  nand2 gate1956(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1957(.a(s_201), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1958(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1959(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1960(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1457(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1458(.a(gate222inter0), .b(s_130), .O(gate222inter1));
  and2  gate1459(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1460(.a(s_130), .O(gate222inter3));
  inv1  gate1461(.a(s_131), .O(gate222inter4));
  nand2 gate1462(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1463(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1464(.a(G632), .O(gate222inter7));
  inv1  gate1465(.a(G684), .O(gate222inter8));
  nand2 gate1466(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1467(.a(s_131), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1468(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1469(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1470(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1891(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1892(.a(gate223inter0), .b(s_192), .O(gate223inter1));
  and2  gate1893(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1894(.a(s_192), .O(gate223inter3));
  inv1  gate1895(.a(s_193), .O(gate223inter4));
  nand2 gate1896(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1897(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1898(.a(G627), .O(gate223inter7));
  inv1  gate1899(.a(G687), .O(gate223inter8));
  nand2 gate1900(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1901(.a(s_193), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1902(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1903(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1904(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1177(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1178(.a(gate224inter0), .b(s_90), .O(gate224inter1));
  and2  gate1179(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1180(.a(s_90), .O(gate224inter3));
  inv1  gate1181(.a(s_91), .O(gate224inter4));
  nand2 gate1182(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1183(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1184(.a(G637), .O(gate224inter7));
  inv1  gate1185(.a(G687), .O(gate224inter8));
  nand2 gate1186(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1187(.a(s_91), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1188(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1189(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1190(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate743(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate744(.a(gate225inter0), .b(s_28), .O(gate225inter1));
  and2  gate745(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate746(.a(s_28), .O(gate225inter3));
  inv1  gate747(.a(s_29), .O(gate225inter4));
  nand2 gate748(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate749(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate750(.a(G690), .O(gate225inter7));
  inv1  gate751(.a(G691), .O(gate225inter8));
  nand2 gate752(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate753(.a(s_29), .b(gate225inter3), .O(gate225inter10));
  nor2  gate754(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate755(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate756(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate813(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate814(.a(gate226inter0), .b(s_38), .O(gate226inter1));
  and2  gate815(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate816(.a(s_38), .O(gate226inter3));
  inv1  gate817(.a(s_39), .O(gate226inter4));
  nand2 gate818(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate819(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate820(.a(G692), .O(gate226inter7));
  inv1  gate821(.a(G693), .O(gate226inter8));
  nand2 gate822(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate823(.a(s_39), .b(gate226inter3), .O(gate226inter10));
  nor2  gate824(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate825(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate826(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1625(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1626(.a(gate229inter0), .b(s_154), .O(gate229inter1));
  and2  gate1627(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1628(.a(s_154), .O(gate229inter3));
  inv1  gate1629(.a(s_155), .O(gate229inter4));
  nand2 gate1630(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1631(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1632(.a(G698), .O(gate229inter7));
  inv1  gate1633(.a(G699), .O(gate229inter8));
  nand2 gate1634(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1635(.a(s_155), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1636(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1637(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1638(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1639(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1640(.a(gate234inter0), .b(s_156), .O(gate234inter1));
  and2  gate1641(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1642(.a(s_156), .O(gate234inter3));
  inv1  gate1643(.a(s_157), .O(gate234inter4));
  nand2 gate1644(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1645(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1646(.a(G245), .O(gate234inter7));
  inv1  gate1647(.a(G721), .O(gate234inter8));
  nand2 gate1648(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1649(.a(s_157), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1650(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1651(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1652(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1933(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1934(.a(gate240inter0), .b(s_198), .O(gate240inter1));
  and2  gate1935(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1936(.a(s_198), .O(gate240inter3));
  inv1  gate1937(.a(s_199), .O(gate240inter4));
  nand2 gate1938(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1939(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1940(.a(G263), .O(gate240inter7));
  inv1  gate1941(.a(G715), .O(gate240inter8));
  nand2 gate1942(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1943(.a(s_199), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1944(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1945(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1946(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1555(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1556(.a(gate242inter0), .b(s_144), .O(gate242inter1));
  and2  gate1557(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1558(.a(s_144), .O(gate242inter3));
  inv1  gate1559(.a(s_145), .O(gate242inter4));
  nand2 gate1560(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1561(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1562(.a(G718), .O(gate242inter7));
  inv1  gate1563(.a(G730), .O(gate242inter8));
  nand2 gate1564(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1565(.a(s_145), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1566(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1567(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1568(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1317(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1318(.a(gate243inter0), .b(s_110), .O(gate243inter1));
  and2  gate1319(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1320(.a(s_110), .O(gate243inter3));
  inv1  gate1321(.a(s_111), .O(gate243inter4));
  nand2 gate1322(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1323(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1324(.a(G245), .O(gate243inter7));
  inv1  gate1325(.a(G733), .O(gate243inter8));
  nand2 gate1326(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1327(.a(s_111), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1328(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1329(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1330(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1793(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1794(.a(gate248inter0), .b(s_178), .O(gate248inter1));
  and2  gate1795(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1796(.a(s_178), .O(gate248inter3));
  inv1  gate1797(.a(s_179), .O(gate248inter4));
  nand2 gate1798(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1799(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1800(.a(G727), .O(gate248inter7));
  inv1  gate1801(.a(G739), .O(gate248inter8));
  nand2 gate1802(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1803(.a(s_179), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1804(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1805(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1806(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1135(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1136(.a(gate251inter0), .b(s_84), .O(gate251inter1));
  and2  gate1137(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1138(.a(s_84), .O(gate251inter3));
  inv1  gate1139(.a(s_85), .O(gate251inter4));
  nand2 gate1140(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1141(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1142(.a(G257), .O(gate251inter7));
  inv1  gate1143(.a(G745), .O(gate251inter8));
  nand2 gate1144(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1145(.a(s_85), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1146(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1147(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1148(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate603(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate604(.a(gate253inter0), .b(s_8), .O(gate253inter1));
  and2  gate605(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate606(.a(s_8), .O(gate253inter3));
  inv1  gate607(.a(s_9), .O(gate253inter4));
  nand2 gate608(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate609(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate610(.a(G260), .O(gate253inter7));
  inv1  gate611(.a(G748), .O(gate253inter8));
  nand2 gate612(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate613(.a(s_9), .b(gate253inter3), .O(gate253inter10));
  nor2  gate614(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate615(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate616(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1513(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1514(.a(gate254inter0), .b(s_138), .O(gate254inter1));
  and2  gate1515(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1516(.a(s_138), .O(gate254inter3));
  inv1  gate1517(.a(s_139), .O(gate254inter4));
  nand2 gate1518(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1519(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1520(.a(G712), .O(gate254inter7));
  inv1  gate1521(.a(G748), .O(gate254inter8));
  nand2 gate1522(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1523(.a(s_139), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1524(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1525(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1526(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1261(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1262(.a(gate260inter0), .b(s_102), .O(gate260inter1));
  and2  gate1263(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1264(.a(s_102), .O(gate260inter3));
  inv1  gate1265(.a(s_103), .O(gate260inter4));
  nand2 gate1266(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1267(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1268(.a(G760), .O(gate260inter7));
  inv1  gate1269(.a(G761), .O(gate260inter8));
  nand2 gate1270(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1271(.a(s_103), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1272(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1273(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1274(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1667(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1668(.a(gate263inter0), .b(s_160), .O(gate263inter1));
  and2  gate1669(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1670(.a(s_160), .O(gate263inter3));
  inv1  gate1671(.a(s_161), .O(gate263inter4));
  nand2 gate1672(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1673(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1674(.a(G766), .O(gate263inter7));
  inv1  gate1675(.a(G767), .O(gate263inter8));
  nand2 gate1676(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1677(.a(s_161), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1678(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1679(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1680(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2031(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2032(.a(gate269inter0), .b(s_212), .O(gate269inter1));
  and2  gate2033(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2034(.a(s_212), .O(gate269inter3));
  inv1  gate2035(.a(s_213), .O(gate269inter4));
  nand2 gate2036(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2037(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2038(.a(G654), .O(gate269inter7));
  inv1  gate2039(.a(G782), .O(gate269inter8));
  nand2 gate2040(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2041(.a(s_213), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2042(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2043(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2044(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2157(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2158(.a(gate271inter0), .b(s_230), .O(gate271inter1));
  and2  gate2159(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2160(.a(s_230), .O(gate271inter3));
  inv1  gate2161(.a(s_231), .O(gate271inter4));
  nand2 gate2162(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2163(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2164(.a(G660), .O(gate271inter7));
  inv1  gate2165(.a(G788), .O(gate271inter8));
  nand2 gate2166(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2167(.a(s_231), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2168(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2169(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2170(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2297(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2298(.a(gate274inter0), .b(s_250), .O(gate274inter1));
  and2  gate2299(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2300(.a(s_250), .O(gate274inter3));
  inv1  gate2301(.a(s_251), .O(gate274inter4));
  nand2 gate2302(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2303(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2304(.a(G770), .O(gate274inter7));
  inv1  gate2305(.a(G794), .O(gate274inter8));
  nand2 gate2306(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2307(.a(s_251), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2308(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2309(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2310(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2437(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2438(.a(gate275inter0), .b(s_270), .O(gate275inter1));
  and2  gate2439(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2440(.a(s_270), .O(gate275inter3));
  inv1  gate2441(.a(s_271), .O(gate275inter4));
  nand2 gate2442(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2443(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2444(.a(G645), .O(gate275inter7));
  inv1  gate2445(.a(G797), .O(gate275inter8));
  nand2 gate2446(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2447(.a(s_271), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2448(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2449(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2450(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1695(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1696(.a(gate278inter0), .b(s_164), .O(gate278inter1));
  and2  gate1697(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1698(.a(s_164), .O(gate278inter3));
  inv1  gate1699(.a(s_165), .O(gate278inter4));
  nand2 gate1700(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1701(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1702(.a(G776), .O(gate278inter7));
  inv1  gate1703(.a(G800), .O(gate278inter8));
  nand2 gate1704(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1705(.a(s_165), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1706(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1707(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1708(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1359(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1360(.a(gate286inter0), .b(s_116), .O(gate286inter1));
  and2  gate1361(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1362(.a(s_116), .O(gate286inter3));
  inv1  gate1363(.a(s_117), .O(gate286inter4));
  nand2 gate1364(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1365(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1366(.a(G788), .O(gate286inter7));
  inv1  gate1367(.a(G812), .O(gate286inter8));
  nand2 gate1368(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1369(.a(s_117), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1370(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1371(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1372(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2353(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2354(.a(gate287inter0), .b(s_258), .O(gate287inter1));
  and2  gate2355(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2356(.a(s_258), .O(gate287inter3));
  inv1  gate2357(.a(s_259), .O(gate287inter4));
  nand2 gate2358(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2359(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2360(.a(G663), .O(gate287inter7));
  inv1  gate2361(.a(G815), .O(gate287inter8));
  nand2 gate2362(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2363(.a(s_259), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2364(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2365(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2366(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1247(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1248(.a(gate288inter0), .b(s_100), .O(gate288inter1));
  and2  gate1249(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1250(.a(s_100), .O(gate288inter3));
  inv1  gate1251(.a(s_101), .O(gate288inter4));
  nand2 gate1252(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1253(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1254(.a(G791), .O(gate288inter7));
  inv1  gate1255(.a(G815), .O(gate288inter8));
  nand2 gate1256(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1257(.a(s_101), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1258(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1259(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1260(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1121(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1122(.a(gate289inter0), .b(s_82), .O(gate289inter1));
  and2  gate1123(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1124(.a(s_82), .O(gate289inter3));
  inv1  gate1125(.a(s_83), .O(gate289inter4));
  nand2 gate1126(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1127(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1128(.a(G818), .O(gate289inter7));
  inv1  gate1129(.a(G819), .O(gate289inter8));
  nand2 gate1130(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1131(.a(s_83), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1132(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1133(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1134(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate659(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate660(.a(gate293inter0), .b(s_16), .O(gate293inter1));
  and2  gate661(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate662(.a(s_16), .O(gate293inter3));
  inv1  gate663(.a(s_17), .O(gate293inter4));
  nand2 gate664(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate665(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate666(.a(G828), .O(gate293inter7));
  inv1  gate667(.a(G829), .O(gate293inter8));
  nand2 gate668(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate669(.a(s_17), .b(gate293inter3), .O(gate293inter10));
  nor2  gate670(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate671(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate672(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate799(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate800(.a(gate387inter0), .b(s_36), .O(gate387inter1));
  and2  gate801(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate802(.a(s_36), .O(gate387inter3));
  inv1  gate803(.a(s_37), .O(gate387inter4));
  nand2 gate804(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate805(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate806(.a(G1), .O(gate387inter7));
  inv1  gate807(.a(G1036), .O(gate387inter8));
  nand2 gate808(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate809(.a(s_37), .b(gate387inter3), .O(gate387inter10));
  nor2  gate810(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate811(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate812(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2283(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2284(.a(gate389inter0), .b(s_248), .O(gate389inter1));
  and2  gate2285(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2286(.a(s_248), .O(gate389inter3));
  inv1  gate2287(.a(s_249), .O(gate389inter4));
  nand2 gate2288(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2289(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2290(.a(G3), .O(gate389inter7));
  inv1  gate2291(.a(G1042), .O(gate389inter8));
  nand2 gate2292(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2293(.a(s_249), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2294(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2295(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2296(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate785(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate786(.a(gate390inter0), .b(s_34), .O(gate390inter1));
  and2  gate787(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate788(.a(s_34), .O(gate390inter3));
  inv1  gate789(.a(s_35), .O(gate390inter4));
  nand2 gate790(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate791(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate792(.a(G4), .O(gate390inter7));
  inv1  gate793(.a(G1045), .O(gate390inter8));
  nand2 gate794(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate795(.a(s_35), .b(gate390inter3), .O(gate390inter10));
  nor2  gate796(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate797(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate798(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate771(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate772(.a(gate392inter0), .b(s_32), .O(gate392inter1));
  and2  gate773(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate774(.a(s_32), .O(gate392inter3));
  inv1  gate775(.a(s_33), .O(gate392inter4));
  nand2 gate776(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate777(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate778(.a(G6), .O(gate392inter7));
  inv1  gate779(.a(G1051), .O(gate392inter8));
  nand2 gate780(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate781(.a(s_33), .b(gate392inter3), .O(gate392inter10));
  nor2  gate782(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate783(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate784(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate883(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate884(.a(gate393inter0), .b(s_48), .O(gate393inter1));
  and2  gate885(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate886(.a(s_48), .O(gate393inter3));
  inv1  gate887(.a(s_49), .O(gate393inter4));
  nand2 gate888(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate889(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate890(.a(G7), .O(gate393inter7));
  inv1  gate891(.a(G1054), .O(gate393inter8));
  nand2 gate892(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate893(.a(s_49), .b(gate393inter3), .O(gate393inter10));
  nor2  gate894(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate895(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate896(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2213(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2214(.a(gate394inter0), .b(s_238), .O(gate394inter1));
  and2  gate2215(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2216(.a(s_238), .O(gate394inter3));
  inv1  gate2217(.a(s_239), .O(gate394inter4));
  nand2 gate2218(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2219(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2220(.a(G8), .O(gate394inter7));
  inv1  gate2221(.a(G1057), .O(gate394inter8));
  nand2 gate2222(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2223(.a(s_239), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2224(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2225(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2226(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1345(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1346(.a(gate399inter0), .b(s_114), .O(gate399inter1));
  and2  gate1347(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1348(.a(s_114), .O(gate399inter3));
  inv1  gate1349(.a(s_115), .O(gate399inter4));
  nand2 gate1350(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1351(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1352(.a(G13), .O(gate399inter7));
  inv1  gate1353(.a(G1072), .O(gate399inter8));
  nand2 gate1354(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1355(.a(s_115), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1356(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1357(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1358(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2129(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2130(.a(gate401inter0), .b(s_226), .O(gate401inter1));
  and2  gate2131(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2132(.a(s_226), .O(gate401inter3));
  inv1  gate2133(.a(s_227), .O(gate401inter4));
  nand2 gate2134(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2135(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2136(.a(G15), .O(gate401inter7));
  inv1  gate2137(.a(G1078), .O(gate401inter8));
  nand2 gate2138(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2139(.a(s_227), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2140(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2141(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2142(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1275(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1276(.a(gate402inter0), .b(s_104), .O(gate402inter1));
  and2  gate1277(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1278(.a(s_104), .O(gate402inter3));
  inv1  gate1279(.a(s_105), .O(gate402inter4));
  nand2 gate1280(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1281(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1282(.a(G16), .O(gate402inter7));
  inv1  gate1283(.a(G1081), .O(gate402inter8));
  nand2 gate1284(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1285(.a(s_105), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1286(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1287(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1288(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1863(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1864(.a(gate406inter0), .b(s_188), .O(gate406inter1));
  and2  gate1865(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1866(.a(s_188), .O(gate406inter3));
  inv1  gate1867(.a(s_189), .O(gate406inter4));
  nand2 gate1868(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1869(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1870(.a(G20), .O(gate406inter7));
  inv1  gate1871(.a(G1093), .O(gate406inter8));
  nand2 gate1872(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1873(.a(s_189), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1874(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1875(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1876(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1961(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1962(.a(gate407inter0), .b(s_202), .O(gate407inter1));
  and2  gate1963(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1964(.a(s_202), .O(gate407inter3));
  inv1  gate1965(.a(s_203), .O(gate407inter4));
  nand2 gate1966(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1967(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1968(.a(G21), .O(gate407inter7));
  inv1  gate1969(.a(G1096), .O(gate407inter8));
  nand2 gate1970(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1971(.a(s_203), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1972(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1973(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1974(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1093(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1094(.a(gate408inter0), .b(s_78), .O(gate408inter1));
  and2  gate1095(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1096(.a(s_78), .O(gate408inter3));
  inv1  gate1097(.a(s_79), .O(gate408inter4));
  nand2 gate1098(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1099(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1100(.a(G22), .O(gate408inter7));
  inv1  gate1101(.a(G1099), .O(gate408inter8));
  nand2 gate1102(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1103(.a(s_79), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1104(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1105(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1106(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate547(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate548(.a(gate409inter0), .b(s_0), .O(gate409inter1));
  and2  gate549(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate550(.a(s_0), .O(gate409inter3));
  inv1  gate551(.a(s_1), .O(gate409inter4));
  nand2 gate552(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate553(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate554(.a(G23), .O(gate409inter7));
  inv1  gate555(.a(G1102), .O(gate409inter8));
  nand2 gate556(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate557(.a(s_1), .b(gate409inter3), .O(gate409inter10));
  nor2  gate558(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate559(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate560(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate617(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate618(.a(gate410inter0), .b(s_10), .O(gate410inter1));
  and2  gate619(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate620(.a(s_10), .O(gate410inter3));
  inv1  gate621(.a(s_11), .O(gate410inter4));
  nand2 gate622(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate623(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate624(.a(G24), .O(gate410inter7));
  inv1  gate625(.a(G1105), .O(gate410inter8));
  nand2 gate626(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate627(.a(s_11), .b(gate410inter3), .O(gate410inter10));
  nor2  gate628(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate629(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate630(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1051(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1052(.a(gate411inter0), .b(s_72), .O(gate411inter1));
  and2  gate1053(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1054(.a(s_72), .O(gate411inter3));
  inv1  gate1055(.a(s_73), .O(gate411inter4));
  nand2 gate1056(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1057(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1058(.a(G25), .O(gate411inter7));
  inv1  gate1059(.a(G1108), .O(gate411inter8));
  nand2 gate1060(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1061(.a(s_73), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1062(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1063(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1064(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1485(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1486(.a(gate413inter0), .b(s_134), .O(gate413inter1));
  and2  gate1487(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1488(.a(s_134), .O(gate413inter3));
  inv1  gate1489(.a(s_135), .O(gate413inter4));
  nand2 gate1490(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1491(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1492(.a(G27), .O(gate413inter7));
  inv1  gate1493(.a(G1114), .O(gate413inter8));
  nand2 gate1494(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1495(.a(s_135), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1496(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1497(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1498(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1471(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1472(.a(gate420inter0), .b(s_132), .O(gate420inter1));
  and2  gate1473(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1474(.a(s_132), .O(gate420inter3));
  inv1  gate1475(.a(s_133), .O(gate420inter4));
  nand2 gate1476(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1477(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1478(.a(G1036), .O(gate420inter7));
  inv1  gate1479(.a(G1132), .O(gate420inter8));
  nand2 gate1480(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1481(.a(s_133), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1482(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1483(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1484(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2367(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2368(.a(gate423inter0), .b(s_260), .O(gate423inter1));
  and2  gate2369(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2370(.a(s_260), .O(gate423inter3));
  inv1  gate2371(.a(s_261), .O(gate423inter4));
  nand2 gate2372(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2373(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2374(.a(G3), .O(gate423inter7));
  inv1  gate2375(.a(G1138), .O(gate423inter8));
  nand2 gate2376(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2377(.a(s_261), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2378(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2379(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2380(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2479(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2480(.a(gate427inter0), .b(s_276), .O(gate427inter1));
  and2  gate2481(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2482(.a(s_276), .O(gate427inter3));
  inv1  gate2483(.a(s_277), .O(gate427inter4));
  nand2 gate2484(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2485(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2486(.a(G5), .O(gate427inter7));
  inv1  gate2487(.a(G1144), .O(gate427inter8));
  nand2 gate2488(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2489(.a(s_277), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2490(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2491(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2492(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1597(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1598(.a(gate429inter0), .b(s_150), .O(gate429inter1));
  and2  gate1599(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1600(.a(s_150), .O(gate429inter3));
  inv1  gate1601(.a(s_151), .O(gate429inter4));
  nand2 gate1602(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1603(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1604(.a(G6), .O(gate429inter7));
  inv1  gate1605(.a(G1147), .O(gate429inter8));
  nand2 gate1606(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1607(.a(s_151), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1608(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1609(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1610(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1107(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1108(.a(gate430inter0), .b(s_80), .O(gate430inter1));
  and2  gate1109(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1110(.a(s_80), .O(gate430inter3));
  inv1  gate1111(.a(s_81), .O(gate430inter4));
  nand2 gate1112(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1113(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1114(.a(G1051), .O(gate430inter7));
  inv1  gate1115(.a(G1147), .O(gate430inter8));
  nand2 gate1116(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1117(.a(s_81), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1118(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1119(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1120(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1009(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1010(.a(gate436inter0), .b(s_66), .O(gate436inter1));
  and2  gate1011(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1012(.a(s_66), .O(gate436inter3));
  inv1  gate1013(.a(s_67), .O(gate436inter4));
  nand2 gate1014(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1015(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1016(.a(G1060), .O(gate436inter7));
  inv1  gate1017(.a(G1156), .O(gate436inter8));
  nand2 gate1018(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1019(.a(s_67), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1020(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1021(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1022(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate897(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate898(.a(gate438inter0), .b(s_50), .O(gate438inter1));
  and2  gate899(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate900(.a(s_50), .O(gate438inter3));
  inv1  gate901(.a(s_51), .O(gate438inter4));
  nand2 gate902(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate903(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate904(.a(G1063), .O(gate438inter7));
  inv1  gate905(.a(G1159), .O(gate438inter8));
  nand2 gate906(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate907(.a(s_51), .b(gate438inter3), .O(gate438inter10));
  nor2  gate908(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate909(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate910(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1807(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1808(.a(gate440inter0), .b(s_180), .O(gate440inter1));
  and2  gate1809(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1810(.a(s_180), .O(gate440inter3));
  inv1  gate1811(.a(s_181), .O(gate440inter4));
  nand2 gate1812(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1813(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1814(.a(G1066), .O(gate440inter7));
  inv1  gate1815(.a(G1162), .O(gate440inter8));
  nand2 gate1816(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1817(.a(s_181), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1818(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1819(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1820(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1023(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1024(.a(gate442inter0), .b(s_68), .O(gate442inter1));
  and2  gate1025(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1026(.a(s_68), .O(gate442inter3));
  inv1  gate1027(.a(s_69), .O(gate442inter4));
  nand2 gate1028(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1029(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1030(.a(G1069), .O(gate442inter7));
  inv1  gate1031(.a(G1165), .O(gate442inter8));
  nand2 gate1032(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1033(.a(s_69), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1034(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1035(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1036(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate939(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate940(.a(gate444inter0), .b(s_56), .O(gate444inter1));
  and2  gate941(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate942(.a(s_56), .O(gate444inter3));
  inv1  gate943(.a(s_57), .O(gate444inter4));
  nand2 gate944(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate945(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate946(.a(G1072), .O(gate444inter7));
  inv1  gate947(.a(G1168), .O(gate444inter8));
  nand2 gate948(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate949(.a(s_57), .b(gate444inter3), .O(gate444inter10));
  nor2  gate950(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate951(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate952(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate995(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate996(.a(gate450inter0), .b(s_64), .O(gate450inter1));
  and2  gate997(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate998(.a(s_64), .O(gate450inter3));
  inv1  gate999(.a(s_65), .O(gate450inter4));
  nand2 gate1000(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1001(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1002(.a(G1081), .O(gate450inter7));
  inv1  gate1003(.a(G1177), .O(gate450inter8));
  nand2 gate1004(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1005(.a(s_65), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1006(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1007(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1008(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2451(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2452(.a(gate456inter0), .b(s_272), .O(gate456inter1));
  and2  gate2453(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2454(.a(s_272), .O(gate456inter3));
  inv1  gate2455(.a(s_273), .O(gate456inter4));
  nand2 gate2456(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2457(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2458(.a(G1090), .O(gate456inter7));
  inv1  gate2459(.a(G1186), .O(gate456inter8));
  nand2 gate2460(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2461(.a(s_273), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2462(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2463(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2464(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2269(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2270(.a(gate460inter0), .b(s_246), .O(gate460inter1));
  and2  gate2271(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2272(.a(s_246), .O(gate460inter3));
  inv1  gate2273(.a(s_247), .O(gate460inter4));
  nand2 gate2274(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2275(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2276(.a(G1096), .O(gate460inter7));
  inv1  gate2277(.a(G1192), .O(gate460inter8));
  nand2 gate2278(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2279(.a(s_247), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2280(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2281(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2282(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2381(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2382(.a(gate463inter0), .b(s_262), .O(gate463inter1));
  and2  gate2383(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2384(.a(s_262), .O(gate463inter3));
  inv1  gate2385(.a(s_263), .O(gate463inter4));
  nand2 gate2386(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2387(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2388(.a(G23), .O(gate463inter7));
  inv1  gate2389(.a(G1198), .O(gate463inter8));
  nand2 gate2390(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2391(.a(s_263), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2392(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2393(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2394(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate701(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate702(.a(gate467inter0), .b(s_22), .O(gate467inter1));
  and2  gate703(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate704(.a(s_22), .O(gate467inter3));
  inv1  gate705(.a(s_23), .O(gate467inter4));
  nand2 gate706(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate707(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate708(.a(G25), .O(gate467inter7));
  inv1  gate709(.a(G1204), .O(gate467inter8));
  nand2 gate710(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate711(.a(s_23), .b(gate467inter3), .O(gate467inter10));
  nor2  gate712(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate713(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate714(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate729(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate730(.a(gate472inter0), .b(s_26), .O(gate472inter1));
  and2  gate731(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate732(.a(s_26), .O(gate472inter3));
  inv1  gate733(.a(s_27), .O(gate472inter4));
  nand2 gate734(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate735(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate736(.a(G1114), .O(gate472inter7));
  inv1  gate737(.a(G1210), .O(gate472inter8));
  nand2 gate738(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate739(.a(s_27), .b(gate472inter3), .O(gate472inter10));
  nor2  gate740(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate741(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate742(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1499(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1500(.a(gate475inter0), .b(s_136), .O(gate475inter1));
  and2  gate1501(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1502(.a(s_136), .O(gate475inter3));
  inv1  gate1503(.a(s_137), .O(gate475inter4));
  nand2 gate1504(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1505(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1506(.a(G29), .O(gate475inter7));
  inv1  gate1507(.a(G1216), .O(gate475inter8));
  nand2 gate1508(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1509(.a(s_137), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1510(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1511(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1512(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1849(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1850(.a(gate476inter0), .b(s_186), .O(gate476inter1));
  and2  gate1851(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1852(.a(s_186), .O(gate476inter3));
  inv1  gate1853(.a(s_187), .O(gate476inter4));
  nand2 gate1854(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1855(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1856(.a(G1120), .O(gate476inter7));
  inv1  gate1857(.a(G1216), .O(gate476inter8));
  nand2 gate1858(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1859(.a(s_187), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1860(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1861(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1862(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1233(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1234(.a(gate480inter0), .b(s_98), .O(gate480inter1));
  and2  gate1235(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1236(.a(s_98), .O(gate480inter3));
  inv1  gate1237(.a(s_99), .O(gate480inter4));
  nand2 gate1238(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1239(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1240(.a(G1126), .O(gate480inter7));
  inv1  gate1241(.a(G1222), .O(gate480inter8));
  nand2 gate1242(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1243(.a(s_99), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1244(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1245(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1246(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1289(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1290(.a(gate482inter0), .b(s_106), .O(gate482inter1));
  and2  gate1291(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1292(.a(s_106), .O(gate482inter3));
  inv1  gate1293(.a(s_107), .O(gate482inter4));
  nand2 gate1294(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1295(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1296(.a(G1129), .O(gate482inter7));
  inv1  gate1297(.a(G1225), .O(gate482inter8));
  nand2 gate1298(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1299(.a(s_107), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1300(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1301(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1302(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2311(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2312(.a(gate485inter0), .b(s_252), .O(gate485inter1));
  and2  gate2313(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2314(.a(s_252), .O(gate485inter3));
  inv1  gate2315(.a(s_253), .O(gate485inter4));
  nand2 gate2316(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2317(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2318(.a(G1232), .O(gate485inter7));
  inv1  gate2319(.a(G1233), .O(gate485inter8));
  nand2 gate2320(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2321(.a(s_253), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2322(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2323(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2324(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate2409(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2410(.a(gate494inter0), .b(s_266), .O(gate494inter1));
  and2  gate2411(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2412(.a(s_266), .O(gate494inter3));
  inv1  gate2413(.a(s_267), .O(gate494inter4));
  nand2 gate2414(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2415(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2416(.a(G1250), .O(gate494inter7));
  inv1  gate2417(.a(G1251), .O(gate494inter8));
  nand2 gate2418(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2419(.a(s_267), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2420(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2421(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2422(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2339(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2340(.a(gate496inter0), .b(s_256), .O(gate496inter1));
  and2  gate2341(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2342(.a(s_256), .O(gate496inter3));
  inv1  gate2343(.a(s_257), .O(gate496inter4));
  nand2 gate2344(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2345(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2346(.a(G1254), .O(gate496inter7));
  inv1  gate2347(.a(G1255), .O(gate496inter8));
  nand2 gate2348(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2349(.a(s_257), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2350(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2351(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2352(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate841(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate842(.a(gate497inter0), .b(s_42), .O(gate497inter1));
  and2  gate843(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate844(.a(s_42), .O(gate497inter3));
  inv1  gate845(.a(s_43), .O(gate497inter4));
  nand2 gate846(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate847(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate848(.a(G1256), .O(gate497inter7));
  inv1  gate849(.a(G1257), .O(gate497inter8));
  nand2 gate850(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate851(.a(s_43), .b(gate497inter3), .O(gate497inter10));
  nor2  gate852(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate853(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate854(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1611(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1612(.a(gate501inter0), .b(s_152), .O(gate501inter1));
  and2  gate1613(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1614(.a(s_152), .O(gate501inter3));
  inv1  gate1615(.a(s_153), .O(gate501inter4));
  nand2 gate1616(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1617(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1618(.a(G1264), .O(gate501inter7));
  inv1  gate1619(.a(G1265), .O(gate501inter8));
  nand2 gate1620(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1621(.a(s_153), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1622(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1623(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1624(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1401(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1402(.a(gate502inter0), .b(s_122), .O(gate502inter1));
  and2  gate1403(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1404(.a(s_122), .O(gate502inter3));
  inv1  gate1405(.a(s_123), .O(gate502inter4));
  nand2 gate1406(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1407(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1408(.a(G1266), .O(gate502inter7));
  inv1  gate1409(.a(G1267), .O(gate502inter8));
  nand2 gate1410(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1411(.a(s_123), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1412(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1413(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1414(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1779(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1780(.a(gate504inter0), .b(s_176), .O(gate504inter1));
  and2  gate1781(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1782(.a(s_176), .O(gate504inter3));
  inv1  gate1783(.a(s_177), .O(gate504inter4));
  nand2 gate1784(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1785(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1786(.a(G1270), .O(gate504inter7));
  inv1  gate1787(.a(G1271), .O(gate504inter8));
  nand2 gate1788(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1789(.a(s_177), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1790(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1791(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1792(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2115(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2116(.a(gate506inter0), .b(s_224), .O(gate506inter1));
  and2  gate2117(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2118(.a(s_224), .O(gate506inter3));
  inv1  gate2119(.a(s_225), .O(gate506inter4));
  nand2 gate2120(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2121(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2122(.a(G1274), .O(gate506inter7));
  inv1  gate2123(.a(G1275), .O(gate506inter8));
  nand2 gate2124(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2125(.a(s_225), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2126(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2127(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2128(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate911(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate912(.a(gate508inter0), .b(s_52), .O(gate508inter1));
  and2  gate913(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate914(.a(s_52), .O(gate508inter3));
  inv1  gate915(.a(s_53), .O(gate508inter4));
  nand2 gate916(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate917(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate918(.a(G1278), .O(gate508inter7));
  inv1  gate919(.a(G1279), .O(gate508inter8));
  nand2 gate920(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate921(.a(s_53), .b(gate508inter3), .O(gate508inter10));
  nor2  gate922(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate923(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate924(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1527(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1528(.a(gate510inter0), .b(s_140), .O(gate510inter1));
  and2  gate1529(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1530(.a(s_140), .O(gate510inter3));
  inv1  gate1531(.a(s_141), .O(gate510inter4));
  nand2 gate1532(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1533(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1534(.a(G1282), .O(gate510inter7));
  inv1  gate1535(.a(G1283), .O(gate510inter8));
  nand2 gate1536(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1537(.a(s_141), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1538(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1539(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1540(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1415(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1416(.a(gate514inter0), .b(s_124), .O(gate514inter1));
  and2  gate1417(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1418(.a(s_124), .O(gate514inter3));
  inv1  gate1419(.a(s_125), .O(gate514inter4));
  nand2 gate1420(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1421(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1422(.a(G1290), .O(gate514inter7));
  inv1  gate1423(.a(G1291), .O(gate514inter8));
  nand2 gate1424(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1425(.a(s_125), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1426(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1427(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1428(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule