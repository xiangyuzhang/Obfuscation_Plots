module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381, s_382, s_383, s_384, s_385, s_386, s_387, s_388, s_389, s_390, s_391, s_392, s_393, s_394, s_395, s_396, s_397, s_398, s_399, s_400, s_401;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1597(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1598(.a(gate9inter0), .b(s_150), .O(gate9inter1));
  and2  gate1599(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1600(.a(s_150), .O(gate9inter3));
  inv1  gate1601(.a(s_151), .O(gate9inter4));
  nand2 gate1602(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1603(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1604(.a(G1), .O(gate9inter7));
  inv1  gate1605(.a(G2), .O(gate9inter8));
  nand2 gate1606(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1607(.a(s_151), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1608(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1609(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1610(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate715(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate716(.a(gate12inter0), .b(s_24), .O(gate12inter1));
  and2  gate717(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate718(.a(s_24), .O(gate12inter3));
  inv1  gate719(.a(s_25), .O(gate12inter4));
  nand2 gate720(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate721(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate722(.a(G7), .O(gate12inter7));
  inv1  gate723(.a(G8), .O(gate12inter8));
  nand2 gate724(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate725(.a(s_25), .b(gate12inter3), .O(gate12inter10));
  nor2  gate726(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate727(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate728(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2423(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2424(.a(gate17inter0), .b(s_268), .O(gate17inter1));
  and2  gate2425(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2426(.a(s_268), .O(gate17inter3));
  inv1  gate2427(.a(s_269), .O(gate17inter4));
  nand2 gate2428(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2429(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2430(.a(G17), .O(gate17inter7));
  inv1  gate2431(.a(G18), .O(gate17inter8));
  nand2 gate2432(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2433(.a(s_269), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2434(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2435(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2436(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate841(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate842(.a(gate21inter0), .b(s_42), .O(gate21inter1));
  and2  gate843(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate844(.a(s_42), .O(gate21inter3));
  inv1  gate845(.a(s_43), .O(gate21inter4));
  nand2 gate846(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate847(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate848(.a(G25), .O(gate21inter7));
  inv1  gate849(.a(G26), .O(gate21inter8));
  nand2 gate850(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate851(.a(s_43), .b(gate21inter3), .O(gate21inter10));
  nor2  gate852(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate853(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate854(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2983(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2984(.a(gate26inter0), .b(s_348), .O(gate26inter1));
  and2  gate2985(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2986(.a(s_348), .O(gate26inter3));
  inv1  gate2987(.a(s_349), .O(gate26inter4));
  nand2 gate2988(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2989(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2990(.a(G9), .O(gate26inter7));
  inv1  gate2991(.a(G13), .O(gate26inter8));
  nand2 gate2992(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2993(.a(s_349), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2994(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2995(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2996(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1751(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1752(.a(gate28inter0), .b(s_172), .O(gate28inter1));
  and2  gate1753(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1754(.a(s_172), .O(gate28inter3));
  inv1  gate1755(.a(s_173), .O(gate28inter4));
  nand2 gate1756(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1757(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1758(.a(G10), .O(gate28inter7));
  inv1  gate1759(.a(G14), .O(gate28inter8));
  nand2 gate1760(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1761(.a(s_173), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1762(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1763(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1764(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1527(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1528(.a(gate29inter0), .b(s_140), .O(gate29inter1));
  and2  gate1529(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1530(.a(s_140), .O(gate29inter3));
  inv1  gate1531(.a(s_141), .O(gate29inter4));
  nand2 gate1532(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1533(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1534(.a(G3), .O(gate29inter7));
  inv1  gate1535(.a(G7), .O(gate29inter8));
  nand2 gate1536(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1537(.a(s_141), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1538(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1539(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1540(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1821(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1822(.a(gate31inter0), .b(s_182), .O(gate31inter1));
  and2  gate1823(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1824(.a(s_182), .O(gate31inter3));
  inv1  gate1825(.a(s_183), .O(gate31inter4));
  nand2 gate1826(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1827(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1828(.a(G4), .O(gate31inter7));
  inv1  gate1829(.a(G8), .O(gate31inter8));
  nand2 gate1830(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1831(.a(s_183), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1832(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1833(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1834(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2395(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2396(.a(gate35inter0), .b(s_264), .O(gate35inter1));
  and2  gate2397(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2398(.a(s_264), .O(gate35inter3));
  inv1  gate2399(.a(s_265), .O(gate35inter4));
  nand2 gate2400(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2401(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2402(.a(G18), .O(gate35inter7));
  inv1  gate2403(.a(G22), .O(gate35inter8));
  nand2 gate2404(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2405(.a(s_265), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2406(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2407(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2408(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1765(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1766(.a(gate37inter0), .b(s_174), .O(gate37inter1));
  and2  gate1767(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1768(.a(s_174), .O(gate37inter3));
  inv1  gate1769(.a(s_175), .O(gate37inter4));
  nand2 gate1770(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1771(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1772(.a(G19), .O(gate37inter7));
  inv1  gate1773(.a(G23), .O(gate37inter8));
  nand2 gate1774(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1775(.a(s_175), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1776(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1777(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1778(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1331(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1332(.a(gate41inter0), .b(s_112), .O(gate41inter1));
  and2  gate1333(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1334(.a(s_112), .O(gate41inter3));
  inv1  gate1335(.a(s_113), .O(gate41inter4));
  nand2 gate1336(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1337(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1338(.a(G1), .O(gate41inter7));
  inv1  gate1339(.a(G266), .O(gate41inter8));
  nand2 gate1340(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1341(.a(s_113), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1342(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1343(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1344(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2255(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2256(.a(gate42inter0), .b(s_244), .O(gate42inter1));
  and2  gate2257(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2258(.a(s_244), .O(gate42inter3));
  inv1  gate2259(.a(s_245), .O(gate42inter4));
  nand2 gate2260(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2261(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2262(.a(G2), .O(gate42inter7));
  inv1  gate2263(.a(G266), .O(gate42inter8));
  nand2 gate2264(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2265(.a(s_245), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2266(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2267(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2268(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate2731(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2732(.a(gate43inter0), .b(s_312), .O(gate43inter1));
  and2  gate2733(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2734(.a(s_312), .O(gate43inter3));
  inv1  gate2735(.a(s_313), .O(gate43inter4));
  nand2 gate2736(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2737(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2738(.a(G3), .O(gate43inter7));
  inv1  gate2739(.a(G269), .O(gate43inter8));
  nand2 gate2740(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2741(.a(s_313), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2742(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2743(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2744(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1373(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1374(.a(gate44inter0), .b(s_118), .O(gate44inter1));
  and2  gate1375(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1376(.a(s_118), .O(gate44inter3));
  inv1  gate1377(.a(s_119), .O(gate44inter4));
  nand2 gate1378(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1379(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1380(.a(G4), .O(gate44inter7));
  inv1  gate1381(.a(G269), .O(gate44inter8));
  nand2 gate1382(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1383(.a(s_119), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1384(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1385(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1386(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2717(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2718(.a(gate45inter0), .b(s_310), .O(gate45inter1));
  and2  gate2719(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2720(.a(s_310), .O(gate45inter3));
  inv1  gate2721(.a(s_311), .O(gate45inter4));
  nand2 gate2722(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2723(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2724(.a(G5), .O(gate45inter7));
  inv1  gate2725(.a(G272), .O(gate45inter8));
  nand2 gate2726(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2727(.a(s_311), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2728(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2729(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2730(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1611(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1612(.a(gate46inter0), .b(s_152), .O(gate46inter1));
  and2  gate1613(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1614(.a(s_152), .O(gate46inter3));
  inv1  gate1615(.a(s_153), .O(gate46inter4));
  nand2 gate1616(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1617(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1618(.a(G6), .O(gate46inter7));
  inv1  gate1619(.a(G272), .O(gate46inter8));
  nand2 gate1620(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1621(.a(s_153), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1622(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1623(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1624(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1709(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1710(.a(gate49inter0), .b(s_166), .O(gate49inter1));
  and2  gate1711(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1712(.a(s_166), .O(gate49inter3));
  inv1  gate1713(.a(s_167), .O(gate49inter4));
  nand2 gate1714(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1715(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1716(.a(G9), .O(gate49inter7));
  inv1  gate1717(.a(G278), .O(gate49inter8));
  nand2 gate1718(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1719(.a(s_167), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1720(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1721(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1722(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1541(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1542(.a(gate55inter0), .b(s_142), .O(gate55inter1));
  and2  gate1543(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1544(.a(s_142), .O(gate55inter3));
  inv1  gate1545(.a(s_143), .O(gate55inter4));
  nand2 gate1546(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1547(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1548(.a(G15), .O(gate55inter7));
  inv1  gate1549(.a(G287), .O(gate55inter8));
  nand2 gate1550(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1551(.a(s_143), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1552(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1553(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1554(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1863(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1864(.a(gate57inter0), .b(s_188), .O(gate57inter1));
  and2  gate1865(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1866(.a(s_188), .O(gate57inter3));
  inv1  gate1867(.a(s_189), .O(gate57inter4));
  nand2 gate1868(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1869(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1870(.a(G17), .O(gate57inter7));
  inv1  gate1871(.a(G290), .O(gate57inter8));
  nand2 gate1872(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1873(.a(s_189), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1874(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1875(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1876(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate3151(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate3152(.a(gate58inter0), .b(s_372), .O(gate58inter1));
  and2  gate3153(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate3154(.a(s_372), .O(gate58inter3));
  inv1  gate3155(.a(s_373), .O(gate58inter4));
  nand2 gate3156(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate3157(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate3158(.a(G18), .O(gate58inter7));
  inv1  gate3159(.a(G290), .O(gate58inter8));
  nand2 gate3160(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate3161(.a(s_373), .b(gate58inter3), .O(gate58inter10));
  nor2  gate3162(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate3163(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate3164(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1289(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1290(.a(gate60inter0), .b(s_106), .O(gate60inter1));
  and2  gate1291(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1292(.a(s_106), .O(gate60inter3));
  inv1  gate1293(.a(s_107), .O(gate60inter4));
  nand2 gate1294(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1295(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1296(.a(G20), .O(gate60inter7));
  inv1  gate1297(.a(G293), .O(gate60inter8));
  nand2 gate1298(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1299(.a(s_107), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1300(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1301(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1302(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate617(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate618(.a(gate61inter0), .b(s_10), .O(gate61inter1));
  and2  gate619(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate620(.a(s_10), .O(gate61inter3));
  inv1  gate621(.a(s_11), .O(gate61inter4));
  nand2 gate622(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate623(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate624(.a(G21), .O(gate61inter7));
  inv1  gate625(.a(G296), .O(gate61inter8));
  nand2 gate626(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate627(.a(s_11), .b(gate61inter3), .O(gate61inter10));
  nor2  gate628(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate629(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate630(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2115(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2116(.a(gate62inter0), .b(s_224), .O(gate62inter1));
  and2  gate2117(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2118(.a(s_224), .O(gate62inter3));
  inv1  gate2119(.a(s_225), .O(gate62inter4));
  nand2 gate2120(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2121(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2122(.a(G22), .O(gate62inter7));
  inv1  gate2123(.a(G296), .O(gate62inter8));
  nand2 gate2124(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2125(.a(s_225), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2126(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2127(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2128(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2773(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2774(.a(gate63inter0), .b(s_318), .O(gate63inter1));
  and2  gate2775(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2776(.a(s_318), .O(gate63inter3));
  inv1  gate2777(.a(s_319), .O(gate63inter4));
  nand2 gate2778(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2779(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2780(.a(G23), .O(gate63inter7));
  inv1  gate2781(.a(G299), .O(gate63inter8));
  nand2 gate2782(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2783(.a(s_319), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2784(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2785(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2786(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2297(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2298(.a(gate64inter0), .b(s_250), .O(gate64inter1));
  and2  gate2299(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2300(.a(s_250), .O(gate64inter3));
  inv1  gate2301(.a(s_251), .O(gate64inter4));
  nand2 gate2302(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2303(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2304(.a(G24), .O(gate64inter7));
  inv1  gate2305(.a(G299), .O(gate64inter8));
  nand2 gate2306(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2307(.a(s_251), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2308(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2309(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2310(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2969(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2970(.a(gate67inter0), .b(s_346), .O(gate67inter1));
  and2  gate2971(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2972(.a(s_346), .O(gate67inter3));
  inv1  gate2973(.a(s_347), .O(gate67inter4));
  nand2 gate2974(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2975(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2976(.a(G27), .O(gate67inter7));
  inv1  gate2977(.a(G305), .O(gate67inter8));
  nand2 gate2978(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2979(.a(s_347), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2980(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2981(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2982(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1905(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1906(.a(gate68inter0), .b(s_194), .O(gate68inter1));
  and2  gate1907(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1908(.a(s_194), .O(gate68inter3));
  inv1  gate1909(.a(s_195), .O(gate68inter4));
  nand2 gate1910(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1911(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1912(.a(G28), .O(gate68inter7));
  inv1  gate1913(.a(G305), .O(gate68inter8));
  nand2 gate1914(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1915(.a(s_195), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1916(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1917(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1918(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate1499(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1500(.a(gate69inter0), .b(s_136), .O(gate69inter1));
  and2  gate1501(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1502(.a(s_136), .O(gate69inter3));
  inv1  gate1503(.a(s_137), .O(gate69inter4));
  nand2 gate1504(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1505(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1506(.a(G29), .O(gate69inter7));
  inv1  gate1507(.a(G308), .O(gate69inter8));
  nand2 gate1508(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1509(.a(s_137), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1510(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1511(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1512(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate547(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate548(.a(gate73inter0), .b(s_0), .O(gate73inter1));
  and2  gate549(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate550(.a(s_0), .O(gate73inter3));
  inv1  gate551(.a(s_1), .O(gate73inter4));
  nand2 gate552(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate553(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate554(.a(G1), .O(gate73inter7));
  inv1  gate555(.a(G314), .O(gate73inter8));
  nand2 gate556(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate557(.a(s_1), .b(gate73inter3), .O(gate73inter10));
  nor2  gate558(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate559(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate560(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate3305(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate3306(.a(gate75inter0), .b(s_394), .O(gate75inter1));
  and2  gate3307(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate3308(.a(s_394), .O(gate75inter3));
  inv1  gate3309(.a(s_395), .O(gate75inter4));
  nand2 gate3310(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate3311(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate3312(.a(G9), .O(gate75inter7));
  inv1  gate3313(.a(G317), .O(gate75inter8));
  nand2 gate3314(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate3315(.a(s_395), .b(gate75inter3), .O(gate75inter10));
  nor2  gate3316(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate3317(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate3318(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1093(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1094(.a(gate76inter0), .b(s_78), .O(gate76inter1));
  and2  gate1095(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1096(.a(s_78), .O(gate76inter3));
  inv1  gate1097(.a(s_79), .O(gate76inter4));
  nand2 gate1098(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1099(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1100(.a(G13), .O(gate76inter7));
  inv1  gate1101(.a(G317), .O(gate76inter8));
  nand2 gate1102(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1103(.a(s_79), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1104(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1105(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1106(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2759(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2760(.a(gate78inter0), .b(s_316), .O(gate78inter1));
  and2  gate2761(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2762(.a(s_316), .O(gate78inter3));
  inv1  gate2763(.a(s_317), .O(gate78inter4));
  nand2 gate2764(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2765(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2766(.a(G6), .O(gate78inter7));
  inv1  gate2767(.a(G320), .O(gate78inter8));
  nand2 gate2768(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2769(.a(s_317), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2770(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2771(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2772(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2577(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2578(.a(gate81inter0), .b(s_290), .O(gate81inter1));
  and2  gate2579(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2580(.a(s_290), .O(gate81inter3));
  inv1  gate2581(.a(s_291), .O(gate81inter4));
  nand2 gate2582(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2583(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2584(.a(G3), .O(gate81inter7));
  inv1  gate2585(.a(G326), .O(gate81inter8));
  nand2 gate2586(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2587(.a(s_291), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2588(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2589(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2590(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate631(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate632(.a(gate83inter0), .b(s_12), .O(gate83inter1));
  and2  gate633(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate634(.a(s_12), .O(gate83inter3));
  inv1  gate635(.a(s_13), .O(gate83inter4));
  nand2 gate636(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate637(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate638(.a(G11), .O(gate83inter7));
  inv1  gate639(.a(G329), .O(gate83inter8));
  nand2 gate640(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate641(.a(s_13), .b(gate83inter3), .O(gate83inter10));
  nor2  gate642(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate643(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate644(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2493(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2494(.a(gate86inter0), .b(s_278), .O(gate86inter1));
  and2  gate2495(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2496(.a(s_278), .O(gate86inter3));
  inv1  gate2497(.a(s_279), .O(gate86inter4));
  nand2 gate2498(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2499(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2500(.a(G8), .O(gate86inter7));
  inv1  gate2501(.a(G332), .O(gate86inter8));
  nand2 gate2502(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2503(.a(s_279), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2504(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2505(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2506(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1681(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1682(.a(gate88inter0), .b(s_162), .O(gate88inter1));
  and2  gate1683(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1684(.a(s_162), .O(gate88inter3));
  inv1  gate1685(.a(s_163), .O(gate88inter4));
  nand2 gate1686(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1687(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1688(.a(G16), .O(gate88inter7));
  inv1  gate1689(.a(G335), .O(gate88inter8));
  nand2 gate1690(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1691(.a(s_163), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1692(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1693(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1694(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2017(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2018(.a(gate91inter0), .b(s_210), .O(gate91inter1));
  and2  gate2019(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2020(.a(s_210), .O(gate91inter3));
  inv1  gate2021(.a(s_211), .O(gate91inter4));
  nand2 gate2022(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2023(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2024(.a(G25), .O(gate91inter7));
  inv1  gate2025(.a(G341), .O(gate91inter8));
  nand2 gate2026(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2027(.a(s_211), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2028(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2029(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2030(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate883(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate884(.a(gate93inter0), .b(s_48), .O(gate93inter1));
  and2  gate885(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate886(.a(s_48), .O(gate93inter3));
  inv1  gate887(.a(s_49), .O(gate93inter4));
  nand2 gate888(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate889(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate890(.a(G18), .O(gate93inter7));
  inv1  gate891(.a(G344), .O(gate93inter8));
  nand2 gate892(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate893(.a(s_49), .b(gate93inter3), .O(gate93inter10));
  nor2  gate894(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate895(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate896(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate3081(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate3082(.a(gate94inter0), .b(s_362), .O(gate94inter1));
  and2  gate3083(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate3084(.a(s_362), .O(gate94inter3));
  inv1  gate3085(.a(s_363), .O(gate94inter4));
  nand2 gate3086(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate3087(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate3088(.a(G22), .O(gate94inter7));
  inv1  gate3089(.a(G344), .O(gate94inter8));
  nand2 gate3090(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate3091(.a(s_363), .b(gate94inter3), .O(gate94inter10));
  nor2  gate3092(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate3093(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate3094(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate799(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate800(.a(gate97inter0), .b(s_36), .O(gate97inter1));
  and2  gate801(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate802(.a(s_36), .O(gate97inter3));
  inv1  gate803(.a(s_37), .O(gate97inter4));
  nand2 gate804(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate805(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate806(.a(G19), .O(gate97inter7));
  inv1  gate807(.a(G350), .O(gate97inter8));
  nand2 gate808(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate809(.a(s_37), .b(gate97inter3), .O(gate97inter10));
  nor2  gate810(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate811(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate812(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2605(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2606(.a(gate99inter0), .b(s_294), .O(gate99inter1));
  and2  gate2607(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2608(.a(s_294), .O(gate99inter3));
  inv1  gate2609(.a(s_295), .O(gate99inter4));
  nand2 gate2610(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2611(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2612(.a(G27), .O(gate99inter7));
  inv1  gate2613(.a(G353), .O(gate99inter8));
  nand2 gate2614(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2615(.a(s_295), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2616(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2617(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2618(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate3039(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate3040(.a(gate100inter0), .b(s_356), .O(gate100inter1));
  and2  gate3041(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate3042(.a(s_356), .O(gate100inter3));
  inv1  gate3043(.a(s_357), .O(gate100inter4));
  nand2 gate3044(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate3045(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate3046(.a(G31), .O(gate100inter7));
  inv1  gate3047(.a(G353), .O(gate100inter8));
  nand2 gate3048(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate3049(.a(s_357), .b(gate100inter3), .O(gate100inter10));
  nor2  gate3050(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate3051(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate3052(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate771(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate772(.a(gate101inter0), .b(s_32), .O(gate101inter1));
  and2  gate773(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate774(.a(s_32), .O(gate101inter3));
  inv1  gate775(.a(s_33), .O(gate101inter4));
  nand2 gate776(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate777(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate778(.a(G20), .O(gate101inter7));
  inv1  gate779(.a(G356), .O(gate101inter8));
  nand2 gate780(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate781(.a(s_33), .b(gate101inter3), .O(gate101inter10));
  nor2  gate782(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate783(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate784(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate701(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate702(.a(gate103inter0), .b(s_22), .O(gate103inter1));
  and2  gate703(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate704(.a(s_22), .O(gate103inter3));
  inv1  gate705(.a(s_23), .O(gate103inter4));
  nand2 gate706(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate707(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate708(.a(G28), .O(gate103inter7));
  inv1  gate709(.a(G359), .O(gate103inter8));
  nand2 gate710(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate711(.a(s_23), .b(gate103inter3), .O(gate103inter10));
  nor2  gate712(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate713(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate714(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2325(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2326(.a(gate104inter0), .b(s_254), .O(gate104inter1));
  and2  gate2327(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2328(.a(s_254), .O(gate104inter3));
  inv1  gate2329(.a(s_255), .O(gate104inter4));
  nand2 gate2330(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2331(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2332(.a(G32), .O(gate104inter7));
  inv1  gate2333(.a(G359), .O(gate104inter8));
  nand2 gate2334(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2335(.a(s_255), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2336(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2337(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2338(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1107(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1108(.a(gate107inter0), .b(s_80), .O(gate107inter1));
  and2  gate1109(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1110(.a(s_80), .O(gate107inter3));
  inv1  gate1111(.a(s_81), .O(gate107inter4));
  nand2 gate1112(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1113(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1114(.a(G366), .O(gate107inter7));
  inv1  gate1115(.a(G367), .O(gate107inter8));
  nand2 gate1116(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1117(.a(s_81), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1118(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1119(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1120(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2367(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2368(.a(gate110inter0), .b(s_260), .O(gate110inter1));
  and2  gate2369(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2370(.a(s_260), .O(gate110inter3));
  inv1  gate2371(.a(s_261), .O(gate110inter4));
  nand2 gate2372(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2373(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2374(.a(G372), .O(gate110inter7));
  inv1  gate2375(.a(G373), .O(gate110inter8));
  nand2 gate2376(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2377(.a(s_261), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2378(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2379(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2380(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2507(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2508(.a(gate112inter0), .b(s_280), .O(gate112inter1));
  and2  gate2509(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2510(.a(s_280), .O(gate112inter3));
  inv1  gate2511(.a(s_281), .O(gate112inter4));
  nand2 gate2512(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2513(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2514(.a(G376), .O(gate112inter7));
  inv1  gate2515(.a(G377), .O(gate112inter8));
  nand2 gate2516(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2517(.a(s_281), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2518(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2519(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2520(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate575(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate576(.a(gate114inter0), .b(s_4), .O(gate114inter1));
  and2  gate577(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate578(.a(s_4), .O(gate114inter3));
  inv1  gate579(.a(s_5), .O(gate114inter4));
  nand2 gate580(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate581(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate582(.a(G380), .O(gate114inter7));
  inv1  gate583(.a(G381), .O(gate114inter8));
  nand2 gate584(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate585(.a(s_5), .b(gate114inter3), .O(gate114inter10));
  nor2  gate586(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate587(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate588(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate2927(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2928(.a(gate115inter0), .b(s_340), .O(gate115inter1));
  and2  gate2929(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2930(.a(s_340), .O(gate115inter3));
  inv1  gate2931(.a(s_341), .O(gate115inter4));
  nand2 gate2932(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2933(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2934(.a(G382), .O(gate115inter7));
  inv1  gate2935(.a(G383), .O(gate115inter8));
  nand2 gate2936(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2937(.a(s_341), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2938(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2939(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2940(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate2437(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2438(.a(gate116inter0), .b(s_270), .O(gate116inter1));
  and2  gate2439(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2440(.a(s_270), .O(gate116inter3));
  inv1  gate2441(.a(s_271), .O(gate116inter4));
  nand2 gate2442(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2443(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2444(.a(G384), .O(gate116inter7));
  inv1  gate2445(.a(G385), .O(gate116inter8));
  nand2 gate2446(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2447(.a(s_271), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2448(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2449(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2450(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate3137(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate3138(.a(gate118inter0), .b(s_370), .O(gate118inter1));
  and2  gate3139(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate3140(.a(s_370), .O(gate118inter3));
  inv1  gate3141(.a(s_371), .O(gate118inter4));
  nand2 gate3142(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate3143(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate3144(.a(G388), .O(gate118inter7));
  inv1  gate3145(.a(G389), .O(gate118inter8));
  nand2 gate3146(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate3147(.a(s_371), .b(gate118inter3), .O(gate118inter10));
  nor2  gate3148(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate3149(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate3150(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate673(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate674(.a(gate119inter0), .b(s_18), .O(gate119inter1));
  and2  gate675(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate676(.a(s_18), .O(gate119inter3));
  inv1  gate677(.a(s_19), .O(gate119inter4));
  nand2 gate678(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate679(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate680(.a(G390), .O(gate119inter7));
  inv1  gate681(.a(G391), .O(gate119inter8));
  nand2 gate682(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate683(.a(s_19), .b(gate119inter3), .O(gate119inter10));
  nor2  gate684(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate685(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate686(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2549(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2550(.a(gate122inter0), .b(s_286), .O(gate122inter1));
  and2  gate2551(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2552(.a(s_286), .O(gate122inter3));
  inv1  gate2553(.a(s_287), .O(gate122inter4));
  nand2 gate2554(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2555(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2556(.a(G396), .O(gate122inter7));
  inv1  gate2557(.a(G397), .O(gate122inter8));
  nand2 gate2558(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2559(.a(s_287), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2560(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2561(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2562(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1891(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1892(.a(gate124inter0), .b(s_192), .O(gate124inter1));
  and2  gate1893(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1894(.a(s_192), .O(gate124inter3));
  inv1  gate1895(.a(s_193), .O(gate124inter4));
  nand2 gate1896(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1897(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1898(.a(G400), .O(gate124inter7));
  inv1  gate1899(.a(G401), .O(gate124inter8));
  nand2 gate1900(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1901(.a(s_193), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1902(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1903(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1904(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate3291(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate3292(.a(gate125inter0), .b(s_392), .O(gate125inter1));
  and2  gate3293(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate3294(.a(s_392), .O(gate125inter3));
  inv1  gate3295(.a(s_393), .O(gate125inter4));
  nand2 gate3296(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate3297(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate3298(.a(G402), .O(gate125inter7));
  inv1  gate3299(.a(G403), .O(gate125inter8));
  nand2 gate3300(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate3301(.a(s_393), .b(gate125inter3), .O(gate125inter10));
  nor2  gate3302(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate3303(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate3304(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate561(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate562(.a(gate126inter0), .b(s_2), .O(gate126inter1));
  and2  gate563(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate564(.a(s_2), .O(gate126inter3));
  inv1  gate565(.a(s_3), .O(gate126inter4));
  nand2 gate566(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate567(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate568(.a(G404), .O(gate126inter7));
  inv1  gate569(.a(G405), .O(gate126inter8));
  nand2 gate570(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate571(.a(s_3), .b(gate126inter3), .O(gate126inter10));
  nor2  gate572(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate573(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate574(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1443(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1444(.a(gate128inter0), .b(s_128), .O(gate128inter1));
  and2  gate1445(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1446(.a(s_128), .O(gate128inter3));
  inv1  gate1447(.a(s_129), .O(gate128inter4));
  nand2 gate1448(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1449(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1450(.a(G408), .O(gate128inter7));
  inv1  gate1451(.a(G409), .O(gate128inter8));
  nand2 gate1452(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1453(.a(s_129), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1454(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1455(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1456(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate659(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate660(.a(gate129inter0), .b(s_16), .O(gate129inter1));
  and2  gate661(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate662(.a(s_16), .O(gate129inter3));
  inv1  gate663(.a(s_17), .O(gate129inter4));
  nand2 gate664(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate665(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate666(.a(G410), .O(gate129inter7));
  inv1  gate667(.a(G411), .O(gate129inter8));
  nand2 gate668(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate669(.a(s_17), .b(gate129inter3), .O(gate129inter10));
  nor2  gate670(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate671(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate672(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1037(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1038(.a(gate131inter0), .b(s_70), .O(gate131inter1));
  and2  gate1039(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1040(.a(s_70), .O(gate131inter3));
  inv1  gate1041(.a(s_71), .O(gate131inter4));
  nand2 gate1042(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1043(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1044(.a(G414), .O(gate131inter7));
  inv1  gate1045(.a(G415), .O(gate131inter8));
  nand2 gate1046(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1047(.a(s_71), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1048(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1049(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1050(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate645(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate646(.a(gate134inter0), .b(s_14), .O(gate134inter1));
  and2  gate647(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate648(.a(s_14), .O(gate134inter3));
  inv1  gate649(.a(s_15), .O(gate134inter4));
  nand2 gate650(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate651(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate652(.a(G420), .O(gate134inter7));
  inv1  gate653(.a(G421), .O(gate134inter8));
  nand2 gate654(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate655(.a(s_15), .b(gate134inter3), .O(gate134inter10));
  nor2  gate656(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate657(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate658(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2913(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2914(.a(gate137inter0), .b(s_338), .O(gate137inter1));
  and2  gate2915(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2916(.a(s_338), .O(gate137inter3));
  inv1  gate2917(.a(s_339), .O(gate137inter4));
  nand2 gate2918(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2919(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2920(.a(G426), .O(gate137inter7));
  inv1  gate2921(.a(G429), .O(gate137inter8));
  nand2 gate2922(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2923(.a(s_339), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2924(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2925(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2926(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate3053(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate3054(.a(gate138inter0), .b(s_358), .O(gate138inter1));
  and2  gate3055(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate3056(.a(s_358), .O(gate138inter3));
  inv1  gate3057(.a(s_359), .O(gate138inter4));
  nand2 gate3058(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate3059(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate3060(.a(G432), .O(gate138inter7));
  inv1  gate3061(.a(G435), .O(gate138inter8));
  nand2 gate3062(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate3063(.a(s_359), .b(gate138inter3), .O(gate138inter10));
  nor2  gate3064(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate3065(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate3066(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2227(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2228(.a(gate139inter0), .b(s_240), .O(gate139inter1));
  and2  gate2229(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2230(.a(s_240), .O(gate139inter3));
  inv1  gate2231(.a(s_241), .O(gate139inter4));
  nand2 gate2232(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2233(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2234(.a(G438), .O(gate139inter7));
  inv1  gate2235(.a(G441), .O(gate139inter8));
  nand2 gate2236(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2237(.a(s_241), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2238(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2239(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2240(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2745(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2746(.a(gate141inter0), .b(s_314), .O(gate141inter1));
  and2  gate2747(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2748(.a(s_314), .O(gate141inter3));
  inv1  gate2749(.a(s_315), .O(gate141inter4));
  nand2 gate2750(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2751(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2752(.a(G450), .O(gate141inter7));
  inv1  gate2753(.a(G453), .O(gate141inter8));
  nand2 gate2754(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2755(.a(s_315), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2756(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2757(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2758(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2157(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2158(.a(gate144inter0), .b(s_230), .O(gate144inter1));
  and2  gate2159(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2160(.a(s_230), .O(gate144inter3));
  inv1  gate2161(.a(s_231), .O(gate144inter4));
  nand2 gate2162(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2163(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2164(.a(G468), .O(gate144inter7));
  inv1  gate2165(.a(G471), .O(gate144inter8));
  nand2 gate2166(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2167(.a(s_231), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2168(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2169(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2170(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate3123(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate3124(.a(gate146inter0), .b(s_368), .O(gate146inter1));
  and2  gate3125(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate3126(.a(s_368), .O(gate146inter3));
  inv1  gate3127(.a(s_369), .O(gate146inter4));
  nand2 gate3128(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate3129(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate3130(.a(G480), .O(gate146inter7));
  inv1  gate3131(.a(G483), .O(gate146inter8));
  nand2 gate3132(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate3133(.a(s_369), .b(gate146inter3), .O(gate146inter10));
  nor2  gate3134(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate3135(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate3136(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate3235(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate3236(.a(gate147inter0), .b(s_384), .O(gate147inter1));
  and2  gate3237(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate3238(.a(s_384), .O(gate147inter3));
  inv1  gate3239(.a(s_385), .O(gate147inter4));
  nand2 gate3240(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate3241(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate3242(.a(G486), .O(gate147inter7));
  inv1  gate3243(.a(G489), .O(gate147inter8));
  nand2 gate3244(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate3245(.a(s_385), .b(gate147inter3), .O(gate147inter10));
  nor2  gate3246(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate3247(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate3248(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate687(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate688(.a(gate149inter0), .b(s_20), .O(gate149inter1));
  and2  gate689(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate690(.a(s_20), .O(gate149inter3));
  inv1  gate691(.a(s_21), .O(gate149inter4));
  nand2 gate692(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate693(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate694(.a(G498), .O(gate149inter7));
  inv1  gate695(.a(G501), .O(gate149inter8));
  nand2 gate696(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate697(.a(s_21), .b(gate149inter3), .O(gate149inter10));
  nor2  gate698(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate699(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate700(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2535(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2536(.a(gate153inter0), .b(s_284), .O(gate153inter1));
  and2  gate2537(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2538(.a(s_284), .O(gate153inter3));
  inv1  gate2539(.a(s_285), .O(gate153inter4));
  nand2 gate2540(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2541(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2542(.a(G426), .O(gate153inter7));
  inv1  gate2543(.a(G522), .O(gate153inter8));
  nand2 gate2544(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2545(.a(s_285), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2546(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2547(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2548(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1149(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1150(.a(gate158inter0), .b(s_86), .O(gate158inter1));
  and2  gate1151(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1152(.a(s_86), .O(gate158inter3));
  inv1  gate1153(.a(s_87), .O(gate158inter4));
  nand2 gate1154(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1155(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1156(.a(G441), .O(gate158inter7));
  inv1  gate1157(.a(G528), .O(gate158inter8));
  nand2 gate1158(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1159(.a(s_87), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1160(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1161(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1162(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1457(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1458(.a(gate159inter0), .b(s_130), .O(gate159inter1));
  and2  gate1459(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1460(.a(s_130), .O(gate159inter3));
  inv1  gate1461(.a(s_131), .O(gate159inter4));
  nand2 gate1462(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1463(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1464(.a(G444), .O(gate159inter7));
  inv1  gate1465(.a(G531), .O(gate159inter8));
  nand2 gate1466(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1467(.a(s_131), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1468(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1469(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1470(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2675(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2676(.a(gate160inter0), .b(s_304), .O(gate160inter1));
  and2  gate2677(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2678(.a(s_304), .O(gate160inter3));
  inv1  gate2679(.a(s_305), .O(gate160inter4));
  nand2 gate2680(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2681(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2682(.a(G447), .O(gate160inter7));
  inv1  gate2683(.a(G531), .O(gate160inter8));
  nand2 gate2684(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2685(.a(s_305), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2686(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2687(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2688(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1429(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1430(.a(gate161inter0), .b(s_126), .O(gate161inter1));
  and2  gate1431(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1432(.a(s_126), .O(gate161inter3));
  inv1  gate1433(.a(s_127), .O(gate161inter4));
  nand2 gate1434(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1435(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1436(.a(G450), .O(gate161inter7));
  inv1  gate1437(.a(G534), .O(gate161inter8));
  nand2 gate1438(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1439(.a(s_127), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1440(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1441(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1442(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1933(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1934(.a(gate163inter0), .b(s_198), .O(gate163inter1));
  and2  gate1935(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1936(.a(s_198), .O(gate163inter3));
  inv1  gate1937(.a(s_199), .O(gate163inter4));
  nand2 gate1938(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1939(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1940(.a(G456), .O(gate163inter7));
  inv1  gate1941(.a(G537), .O(gate163inter8));
  nand2 gate1942(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1943(.a(s_199), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1944(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1945(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1946(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2381(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2382(.a(gate174inter0), .b(s_262), .O(gate174inter1));
  and2  gate2383(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2384(.a(s_262), .O(gate174inter3));
  inv1  gate2385(.a(s_263), .O(gate174inter4));
  nand2 gate2386(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2387(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2388(.a(G489), .O(gate174inter7));
  inv1  gate2389(.a(G552), .O(gate174inter8));
  nand2 gate2390(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2391(.a(s_263), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2392(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2393(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2394(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate897(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate898(.a(gate179inter0), .b(s_50), .O(gate179inter1));
  and2  gate899(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate900(.a(s_50), .O(gate179inter3));
  inv1  gate901(.a(s_51), .O(gate179inter4));
  nand2 gate902(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate903(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate904(.a(G504), .O(gate179inter7));
  inv1  gate905(.a(G561), .O(gate179inter8));
  nand2 gate906(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate907(.a(s_51), .b(gate179inter3), .O(gate179inter10));
  nor2  gate908(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate909(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate910(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate3095(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate3096(.a(gate180inter0), .b(s_364), .O(gate180inter1));
  and2  gate3097(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate3098(.a(s_364), .O(gate180inter3));
  inv1  gate3099(.a(s_365), .O(gate180inter4));
  nand2 gate3100(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate3101(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate3102(.a(G507), .O(gate180inter7));
  inv1  gate3103(.a(G561), .O(gate180inter8));
  nand2 gate3104(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate3105(.a(s_365), .b(gate180inter3), .O(gate180inter10));
  nor2  gate3106(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate3107(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate3108(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate855(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate856(.a(gate181inter0), .b(s_44), .O(gate181inter1));
  and2  gate857(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate858(.a(s_44), .O(gate181inter3));
  inv1  gate859(.a(s_45), .O(gate181inter4));
  nand2 gate860(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate861(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate862(.a(G510), .O(gate181inter7));
  inv1  gate863(.a(G564), .O(gate181inter8));
  nand2 gate864(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate865(.a(s_45), .b(gate181inter3), .O(gate181inter10));
  nor2  gate866(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate867(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate868(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1415(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1416(.a(gate182inter0), .b(s_124), .O(gate182inter1));
  and2  gate1417(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1418(.a(s_124), .O(gate182inter3));
  inv1  gate1419(.a(s_125), .O(gate182inter4));
  nand2 gate1420(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1421(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1422(.a(G513), .O(gate182inter7));
  inv1  gate1423(.a(G564), .O(gate182inter8));
  nand2 gate1424(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1425(.a(s_125), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1426(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1427(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1428(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2857(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2858(.a(gate184inter0), .b(s_330), .O(gate184inter1));
  and2  gate2859(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2860(.a(s_330), .O(gate184inter3));
  inv1  gate2861(.a(s_331), .O(gate184inter4));
  nand2 gate2862(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2863(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2864(.a(G519), .O(gate184inter7));
  inv1  gate2865(.a(G567), .O(gate184inter8));
  nand2 gate2866(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2867(.a(s_331), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2868(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2869(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2870(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1779(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1780(.a(gate185inter0), .b(s_176), .O(gate185inter1));
  and2  gate1781(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1782(.a(s_176), .O(gate185inter3));
  inv1  gate1783(.a(s_177), .O(gate185inter4));
  nand2 gate1784(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1785(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1786(.a(G570), .O(gate185inter7));
  inv1  gate1787(.a(G571), .O(gate185inter8));
  nand2 gate1788(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1789(.a(s_177), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1790(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1791(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1792(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1177(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1178(.a(gate186inter0), .b(s_90), .O(gate186inter1));
  and2  gate1179(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1180(.a(s_90), .O(gate186inter3));
  inv1  gate1181(.a(s_91), .O(gate186inter4));
  nand2 gate1182(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1183(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1184(.a(G572), .O(gate186inter7));
  inv1  gate1185(.a(G573), .O(gate186inter8));
  nand2 gate1186(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1187(.a(s_91), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1188(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1189(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1190(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1919(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1920(.a(gate189inter0), .b(s_196), .O(gate189inter1));
  and2  gate1921(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1922(.a(s_196), .O(gate189inter3));
  inv1  gate1923(.a(s_197), .O(gate189inter4));
  nand2 gate1924(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1925(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1926(.a(G578), .O(gate189inter7));
  inv1  gate1927(.a(G579), .O(gate189inter8));
  nand2 gate1928(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1929(.a(s_197), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1930(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1931(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1932(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate939(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate940(.a(gate190inter0), .b(s_56), .O(gate190inter1));
  and2  gate941(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate942(.a(s_56), .O(gate190inter3));
  inv1  gate943(.a(s_57), .O(gate190inter4));
  nand2 gate944(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate945(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate946(.a(G580), .O(gate190inter7));
  inv1  gate947(.a(G581), .O(gate190inter8));
  nand2 gate948(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate949(.a(s_57), .b(gate190inter3), .O(gate190inter10));
  nor2  gate950(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate951(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate952(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate3249(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate3250(.a(gate191inter0), .b(s_386), .O(gate191inter1));
  and2  gate3251(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate3252(.a(s_386), .O(gate191inter3));
  inv1  gate3253(.a(s_387), .O(gate191inter4));
  nand2 gate3254(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate3255(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate3256(.a(G582), .O(gate191inter7));
  inv1  gate3257(.a(G583), .O(gate191inter8));
  nand2 gate3258(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate3259(.a(s_387), .b(gate191inter3), .O(gate191inter10));
  nor2  gate3260(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate3261(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate3262(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2101(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2102(.a(gate193inter0), .b(s_222), .O(gate193inter1));
  and2  gate2103(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2104(.a(s_222), .O(gate193inter3));
  inv1  gate2105(.a(s_223), .O(gate193inter4));
  nand2 gate2106(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2107(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2108(.a(G586), .O(gate193inter7));
  inv1  gate2109(.a(G587), .O(gate193inter8));
  nand2 gate2110(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2111(.a(s_223), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2112(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2113(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2114(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2129(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2130(.a(gate195inter0), .b(s_226), .O(gate195inter1));
  and2  gate2131(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2132(.a(s_226), .O(gate195inter3));
  inv1  gate2133(.a(s_227), .O(gate195inter4));
  nand2 gate2134(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2135(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2136(.a(G590), .O(gate195inter7));
  inv1  gate2137(.a(G591), .O(gate195inter8));
  nand2 gate2138(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2139(.a(s_227), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2140(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2141(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2142(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1485(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1486(.a(gate198inter0), .b(s_134), .O(gate198inter1));
  and2  gate1487(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1488(.a(s_134), .O(gate198inter3));
  inv1  gate1489(.a(s_135), .O(gate198inter4));
  nand2 gate1490(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1491(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1492(.a(G596), .O(gate198inter7));
  inv1  gate1493(.a(G597), .O(gate198inter8));
  nand2 gate1494(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1495(.a(s_135), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1496(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1497(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1498(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1667(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1668(.a(gate199inter0), .b(s_160), .O(gate199inter1));
  and2  gate1669(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1670(.a(s_160), .O(gate199inter3));
  inv1  gate1671(.a(s_161), .O(gate199inter4));
  nand2 gate1672(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1673(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1674(.a(G598), .O(gate199inter7));
  inv1  gate1675(.a(G599), .O(gate199inter8));
  nand2 gate1676(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1677(.a(s_161), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1678(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1679(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1680(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1317(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1318(.a(gate200inter0), .b(s_110), .O(gate200inter1));
  and2  gate1319(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1320(.a(s_110), .O(gate200inter3));
  inv1  gate1321(.a(s_111), .O(gate200inter4));
  nand2 gate1322(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1323(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1324(.a(G600), .O(gate200inter7));
  inv1  gate1325(.a(G601), .O(gate200inter8));
  nand2 gate1326(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1327(.a(s_111), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1328(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1329(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1330(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2703(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2704(.a(gate202inter0), .b(s_308), .O(gate202inter1));
  and2  gate2705(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2706(.a(s_308), .O(gate202inter3));
  inv1  gate2707(.a(s_309), .O(gate202inter4));
  nand2 gate2708(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2709(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2710(.a(G612), .O(gate202inter7));
  inv1  gate2711(.a(G617), .O(gate202inter8));
  nand2 gate2712(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2713(.a(s_309), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2714(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2715(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2716(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2451(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2452(.a(gate204inter0), .b(s_272), .O(gate204inter1));
  and2  gate2453(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2454(.a(s_272), .O(gate204inter3));
  inv1  gate2455(.a(s_273), .O(gate204inter4));
  nand2 gate2456(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2457(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2458(.a(G607), .O(gate204inter7));
  inv1  gate2459(.a(G617), .O(gate204inter8));
  nand2 gate2460(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2461(.a(s_273), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2462(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2463(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2464(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate911(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate912(.a(gate206inter0), .b(s_52), .O(gate206inter1));
  and2  gate913(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate914(.a(s_52), .O(gate206inter3));
  inv1  gate915(.a(s_53), .O(gate206inter4));
  nand2 gate916(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate917(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate918(.a(G632), .O(gate206inter7));
  inv1  gate919(.a(G637), .O(gate206inter8));
  nand2 gate920(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate921(.a(s_53), .b(gate206inter3), .O(gate206inter10));
  nor2  gate922(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate923(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate924(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate925(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate926(.a(gate207inter0), .b(s_54), .O(gate207inter1));
  and2  gate927(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate928(.a(s_54), .O(gate207inter3));
  inv1  gate929(.a(s_55), .O(gate207inter4));
  nand2 gate930(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate931(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate932(.a(G622), .O(gate207inter7));
  inv1  gate933(.a(G632), .O(gate207inter8));
  nand2 gate934(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate935(.a(s_55), .b(gate207inter3), .O(gate207inter10));
  nor2  gate936(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate937(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate938(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1009(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1010(.a(gate208inter0), .b(s_66), .O(gate208inter1));
  and2  gate1011(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1012(.a(s_66), .O(gate208inter3));
  inv1  gate1013(.a(s_67), .O(gate208inter4));
  nand2 gate1014(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1015(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1016(.a(G627), .O(gate208inter7));
  inv1  gate1017(.a(G637), .O(gate208inter8));
  nand2 gate1018(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1019(.a(s_67), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1020(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1021(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1022(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2311(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2312(.a(gate209inter0), .b(s_252), .O(gate209inter1));
  and2  gate2313(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2314(.a(s_252), .O(gate209inter3));
  inv1  gate2315(.a(s_253), .O(gate209inter4));
  nand2 gate2316(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2317(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2318(.a(G602), .O(gate209inter7));
  inv1  gate2319(.a(G666), .O(gate209inter8));
  nand2 gate2320(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2321(.a(s_253), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2322(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2323(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2324(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1947(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1948(.a(gate211inter0), .b(s_200), .O(gate211inter1));
  and2  gate1949(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1950(.a(s_200), .O(gate211inter3));
  inv1  gate1951(.a(s_201), .O(gate211inter4));
  nand2 gate1952(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1953(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1954(.a(G612), .O(gate211inter7));
  inv1  gate1955(.a(G669), .O(gate211inter8));
  nand2 gate1956(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1957(.a(s_201), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1958(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1959(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1960(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1261(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1262(.a(gate212inter0), .b(s_102), .O(gate212inter1));
  and2  gate1263(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1264(.a(s_102), .O(gate212inter3));
  inv1  gate1265(.a(s_103), .O(gate212inter4));
  nand2 gate1266(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1267(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1268(.a(G617), .O(gate212inter7));
  inv1  gate1269(.a(G669), .O(gate212inter8));
  nand2 gate1270(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1271(.a(s_103), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1272(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1273(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1274(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate785(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate786(.a(gate214inter0), .b(s_34), .O(gate214inter1));
  and2  gate787(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate788(.a(s_34), .O(gate214inter3));
  inv1  gate789(.a(s_35), .O(gate214inter4));
  nand2 gate790(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate791(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate792(.a(G612), .O(gate214inter7));
  inv1  gate793(.a(G672), .O(gate214inter8));
  nand2 gate794(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate795(.a(s_35), .b(gate214inter3), .O(gate214inter10));
  nor2  gate796(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate797(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate798(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate967(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate968(.a(gate215inter0), .b(s_60), .O(gate215inter1));
  and2  gate969(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate970(.a(s_60), .O(gate215inter3));
  inv1  gate971(.a(s_61), .O(gate215inter4));
  nand2 gate972(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate973(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate974(.a(G607), .O(gate215inter7));
  inv1  gate975(.a(G675), .O(gate215inter8));
  nand2 gate976(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate977(.a(s_61), .b(gate215inter3), .O(gate215inter10));
  nor2  gate978(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate979(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate980(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1303(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1304(.a(gate216inter0), .b(s_108), .O(gate216inter1));
  and2  gate1305(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1306(.a(s_108), .O(gate216inter3));
  inv1  gate1307(.a(s_109), .O(gate216inter4));
  nand2 gate1308(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1309(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1310(.a(G617), .O(gate216inter7));
  inv1  gate1311(.a(G675), .O(gate216inter8));
  nand2 gate1312(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1313(.a(s_109), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1314(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1315(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1316(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2479(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2480(.a(gate217inter0), .b(s_276), .O(gate217inter1));
  and2  gate2481(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2482(.a(s_276), .O(gate217inter3));
  inv1  gate2483(.a(s_277), .O(gate217inter4));
  nand2 gate2484(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2485(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2486(.a(G622), .O(gate217inter7));
  inv1  gate2487(.a(G678), .O(gate217inter8));
  nand2 gate2488(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2489(.a(s_277), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2490(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2491(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2492(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1555(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1556(.a(gate221inter0), .b(s_144), .O(gate221inter1));
  and2  gate1557(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1558(.a(s_144), .O(gate221inter3));
  inv1  gate1559(.a(s_145), .O(gate221inter4));
  nand2 gate1560(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1561(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1562(.a(G622), .O(gate221inter7));
  inv1  gate1563(.a(G684), .O(gate221inter8));
  nand2 gate1564(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1565(.a(s_145), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1566(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1567(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1568(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate2815(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2816(.a(gate222inter0), .b(s_324), .O(gate222inter1));
  and2  gate2817(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2818(.a(s_324), .O(gate222inter3));
  inv1  gate2819(.a(s_325), .O(gate222inter4));
  nand2 gate2820(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2821(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2822(.a(G632), .O(gate222inter7));
  inv1  gate2823(.a(G684), .O(gate222inter8));
  nand2 gate2824(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2825(.a(s_325), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2826(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2827(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2828(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate3179(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate3180(.a(gate223inter0), .b(s_376), .O(gate223inter1));
  and2  gate3181(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate3182(.a(s_376), .O(gate223inter3));
  inv1  gate3183(.a(s_377), .O(gate223inter4));
  nand2 gate3184(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate3185(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate3186(.a(G627), .O(gate223inter7));
  inv1  gate3187(.a(G687), .O(gate223inter8));
  nand2 gate3188(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate3189(.a(s_377), .b(gate223inter3), .O(gate223inter10));
  nor2  gate3190(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate3191(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate3192(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate729(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate730(.a(gate224inter0), .b(s_26), .O(gate224inter1));
  and2  gate731(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate732(.a(s_26), .O(gate224inter3));
  inv1  gate733(.a(s_27), .O(gate224inter4));
  nand2 gate734(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate735(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate736(.a(G637), .O(gate224inter7));
  inv1  gate737(.a(G687), .O(gate224inter8));
  nand2 gate738(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate739(.a(s_27), .b(gate224inter3), .O(gate224inter10));
  nor2  gate740(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate741(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate742(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate3109(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate3110(.a(gate225inter0), .b(s_366), .O(gate225inter1));
  and2  gate3111(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate3112(.a(s_366), .O(gate225inter3));
  inv1  gate3113(.a(s_367), .O(gate225inter4));
  nand2 gate3114(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate3115(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate3116(.a(G690), .O(gate225inter7));
  inv1  gate3117(.a(G691), .O(gate225inter8));
  nand2 gate3118(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate3119(.a(s_367), .b(gate225inter3), .O(gate225inter10));
  nor2  gate3120(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate3121(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate3122(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate3193(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate3194(.a(gate226inter0), .b(s_378), .O(gate226inter1));
  and2  gate3195(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate3196(.a(s_378), .O(gate226inter3));
  inv1  gate3197(.a(s_379), .O(gate226inter4));
  nand2 gate3198(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate3199(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate3200(.a(G692), .O(gate226inter7));
  inv1  gate3201(.a(G693), .O(gate226inter8));
  nand2 gate3202(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate3203(.a(s_379), .b(gate226inter3), .O(gate226inter10));
  nor2  gate3204(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate3205(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate3206(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1359(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1360(.a(gate228inter0), .b(s_116), .O(gate228inter1));
  and2  gate1361(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1362(.a(s_116), .O(gate228inter3));
  inv1  gate1363(.a(s_117), .O(gate228inter4));
  nand2 gate1364(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1365(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1366(.a(G696), .O(gate228inter7));
  inv1  gate1367(.a(G697), .O(gate228inter8));
  nand2 gate1368(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1369(.a(s_117), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1370(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1371(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1372(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1135(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1136(.a(gate230inter0), .b(s_84), .O(gate230inter1));
  and2  gate1137(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1138(.a(s_84), .O(gate230inter3));
  inv1  gate1139(.a(s_85), .O(gate230inter4));
  nand2 gate1140(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1141(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1142(.a(G700), .O(gate230inter7));
  inv1  gate1143(.a(G701), .O(gate230inter8));
  nand2 gate1144(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1145(.a(s_85), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1146(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1147(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1148(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1513(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1514(.a(gate234inter0), .b(s_138), .O(gate234inter1));
  and2  gate1515(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1516(.a(s_138), .O(gate234inter3));
  inv1  gate1517(.a(s_139), .O(gate234inter4));
  nand2 gate1518(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1519(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1520(.a(G245), .O(gate234inter7));
  inv1  gate1521(.a(G721), .O(gate234inter8));
  nand2 gate1522(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1523(.a(s_139), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1524(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1525(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1526(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1989(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1990(.a(gate235inter0), .b(s_206), .O(gate235inter1));
  and2  gate1991(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1992(.a(s_206), .O(gate235inter3));
  inv1  gate1993(.a(s_207), .O(gate235inter4));
  nand2 gate1994(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1995(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1996(.a(G248), .O(gate235inter7));
  inv1  gate1997(.a(G724), .O(gate235inter8));
  nand2 gate1998(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1999(.a(s_207), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2000(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2001(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2002(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1275(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1276(.a(gate237inter0), .b(s_104), .O(gate237inter1));
  and2  gate1277(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1278(.a(s_104), .O(gate237inter3));
  inv1  gate1279(.a(s_105), .O(gate237inter4));
  nand2 gate1280(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1281(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1282(.a(G254), .O(gate237inter7));
  inv1  gate1283(.a(G706), .O(gate237inter8));
  nand2 gate1284(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1285(.a(s_105), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1286(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1287(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1288(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1247(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1248(.a(gate238inter0), .b(s_100), .O(gate238inter1));
  and2  gate1249(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1250(.a(s_100), .O(gate238inter3));
  inv1  gate1251(.a(s_101), .O(gate238inter4));
  nand2 gate1252(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1253(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1254(.a(G257), .O(gate238inter7));
  inv1  gate1255(.a(G709), .O(gate238inter8));
  nand2 gate1256(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1257(.a(s_101), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1258(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1259(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1260(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate995(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate996(.a(gate239inter0), .b(s_64), .O(gate239inter1));
  and2  gate997(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate998(.a(s_64), .O(gate239inter3));
  inv1  gate999(.a(s_65), .O(gate239inter4));
  nand2 gate1000(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1001(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1002(.a(G260), .O(gate239inter7));
  inv1  gate1003(.a(G712), .O(gate239inter8));
  nand2 gate1004(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1005(.a(s_65), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1006(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1007(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1008(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1961(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1962(.a(gate241inter0), .b(s_202), .O(gate241inter1));
  and2  gate1963(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1964(.a(s_202), .O(gate241inter3));
  inv1  gate1965(.a(s_203), .O(gate241inter4));
  nand2 gate1966(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1967(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1968(.a(G242), .O(gate241inter7));
  inv1  gate1969(.a(G730), .O(gate241inter8));
  nand2 gate1970(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1971(.a(s_203), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1972(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1973(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1974(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2591(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2592(.a(gate243inter0), .b(s_292), .O(gate243inter1));
  and2  gate2593(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2594(.a(s_292), .O(gate243inter3));
  inv1  gate2595(.a(s_293), .O(gate243inter4));
  nand2 gate2596(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2597(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2598(.a(G245), .O(gate243inter7));
  inv1  gate2599(.a(G733), .O(gate243inter8));
  nand2 gate2600(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2601(.a(s_293), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2602(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2603(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2604(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1023(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1024(.a(gate246inter0), .b(s_68), .O(gate246inter1));
  and2  gate1025(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1026(.a(s_68), .O(gate246inter3));
  inv1  gate1027(.a(s_69), .O(gate246inter4));
  nand2 gate1028(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1029(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1030(.a(G724), .O(gate246inter7));
  inv1  gate1031(.a(G736), .O(gate246inter8));
  nand2 gate1032(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1033(.a(s_69), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1034(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1035(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1036(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate3221(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate3222(.a(gate251inter0), .b(s_382), .O(gate251inter1));
  and2  gate3223(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate3224(.a(s_382), .O(gate251inter3));
  inv1  gate3225(.a(s_383), .O(gate251inter4));
  nand2 gate3226(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate3227(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate3228(.a(G257), .O(gate251inter7));
  inv1  gate3229(.a(G745), .O(gate251inter8));
  nand2 gate3230(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate3231(.a(s_383), .b(gate251inter3), .O(gate251inter10));
  nor2  gate3232(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate3233(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate3234(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate2143(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2144(.a(gate252inter0), .b(s_228), .O(gate252inter1));
  and2  gate2145(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2146(.a(s_228), .O(gate252inter3));
  inv1  gate2147(.a(s_229), .O(gate252inter4));
  nand2 gate2148(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2149(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2150(.a(G709), .O(gate252inter7));
  inv1  gate2151(.a(G745), .O(gate252inter8));
  nand2 gate2152(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2153(.a(s_229), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2154(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2155(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2156(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2689(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2690(.a(gate256inter0), .b(s_306), .O(gate256inter1));
  and2  gate2691(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2692(.a(s_306), .O(gate256inter3));
  inv1  gate2693(.a(s_307), .O(gate256inter4));
  nand2 gate2694(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2695(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2696(.a(G715), .O(gate256inter7));
  inv1  gate2697(.a(G751), .O(gate256inter8));
  nand2 gate2698(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2699(.a(s_307), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2700(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2701(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2702(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1065(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1066(.a(gate257inter0), .b(s_74), .O(gate257inter1));
  and2  gate1067(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1068(.a(s_74), .O(gate257inter3));
  inv1  gate1069(.a(s_75), .O(gate257inter4));
  nand2 gate1070(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1071(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1072(.a(G754), .O(gate257inter7));
  inv1  gate1073(.a(G755), .O(gate257inter8));
  nand2 gate1074(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1075(.a(s_75), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1076(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1077(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1078(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate869(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate870(.a(gate260inter0), .b(s_46), .O(gate260inter1));
  and2  gate871(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate872(.a(s_46), .O(gate260inter3));
  inv1  gate873(.a(s_47), .O(gate260inter4));
  nand2 gate874(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate875(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate876(.a(G760), .O(gate260inter7));
  inv1  gate877(.a(G761), .O(gate260inter8));
  nand2 gate878(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate879(.a(s_47), .b(gate260inter3), .O(gate260inter10));
  nor2  gate880(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate881(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate882(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2171(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2172(.a(gate261inter0), .b(s_232), .O(gate261inter1));
  and2  gate2173(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2174(.a(s_232), .O(gate261inter3));
  inv1  gate2175(.a(s_233), .O(gate261inter4));
  nand2 gate2176(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2177(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2178(.a(G762), .O(gate261inter7));
  inv1  gate2179(.a(G763), .O(gate261inter8));
  nand2 gate2180(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2181(.a(s_233), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2182(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2183(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2184(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2899(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2900(.a(gate262inter0), .b(s_336), .O(gate262inter1));
  and2  gate2901(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2902(.a(s_336), .O(gate262inter3));
  inv1  gate2903(.a(s_337), .O(gate262inter4));
  nand2 gate2904(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2905(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2906(.a(G764), .O(gate262inter7));
  inv1  gate2907(.a(G765), .O(gate262inter8));
  nand2 gate2908(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2909(.a(s_337), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2910(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2911(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2912(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate743(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate744(.a(gate263inter0), .b(s_28), .O(gate263inter1));
  and2  gate745(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate746(.a(s_28), .O(gate263inter3));
  inv1  gate747(.a(s_29), .O(gate263inter4));
  nand2 gate748(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate749(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate750(.a(G766), .O(gate263inter7));
  inv1  gate751(.a(G767), .O(gate263inter8));
  nand2 gate752(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate753(.a(s_29), .b(gate263inter3), .O(gate263inter10));
  nor2  gate754(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate755(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate756(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1569(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1570(.a(gate265inter0), .b(s_146), .O(gate265inter1));
  and2  gate1571(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1572(.a(s_146), .O(gate265inter3));
  inv1  gate1573(.a(s_147), .O(gate265inter4));
  nand2 gate1574(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1575(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1576(.a(G642), .O(gate265inter7));
  inv1  gate1577(.a(G770), .O(gate265inter8));
  nand2 gate1578(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1579(.a(s_147), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1580(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1581(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1582(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1121(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1122(.a(gate266inter0), .b(s_82), .O(gate266inter1));
  and2  gate1123(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1124(.a(s_82), .O(gate266inter3));
  inv1  gate1125(.a(s_83), .O(gate266inter4));
  nand2 gate1126(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1127(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1128(.a(G645), .O(gate266inter7));
  inv1  gate1129(.a(G773), .O(gate266inter8));
  nand2 gate1130(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1131(.a(s_83), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1132(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1133(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1134(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1401(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1402(.a(gate267inter0), .b(s_122), .O(gate267inter1));
  and2  gate1403(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1404(.a(s_122), .O(gate267inter3));
  inv1  gate1405(.a(s_123), .O(gate267inter4));
  nand2 gate1406(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1407(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1408(.a(G648), .O(gate267inter7));
  inv1  gate1409(.a(G776), .O(gate267inter8));
  nand2 gate1410(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1411(.a(s_123), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1412(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1413(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1414(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1219(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1220(.a(gate269inter0), .b(s_96), .O(gate269inter1));
  and2  gate1221(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1222(.a(s_96), .O(gate269inter3));
  inv1  gate1223(.a(s_97), .O(gate269inter4));
  nand2 gate1224(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1225(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1226(.a(G654), .O(gate269inter7));
  inv1  gate1227(.a(G782), .O(gate269inter8));
  nand2 gate1228(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1229(.a(s_97), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1230(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1231(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1232(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate2787(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2788(.a(gate270inter0), .b(s_320), .O(gate270inter1));
  and2  gate2789(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2790(.a(s_320), .O(gate270inter3));
  inv1  gate2791(.a(s_321), .O(gate270inter4));
  nand2 gate2792(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2793(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2794(.a(G657), .O(gate270inter7));
  inv1  gate2795(.a(G785), .O(gate270inter8));
  nand2 gate2796(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2797(.a(s_321), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2798(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2799(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2800(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate757(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate758(.a(gate272inter0), .b(s_30), .O(gate272inter1));
  and2  gate759(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate760(.a(s_30), .O(gate272inter3));
  inv1  gate761(.a(s_31), .O(gate272inter4));
  nand2 gate762(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate763(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate764(.a(G663), .O(gate272inter7));
  inv1  gate765(.a(G791), .O(gate272inter8));
  nand2 gate766(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate767(.a(s_31), .b(gate272inter3), .O(gate272inter10));
  nor2  gate768(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate769(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate770(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1191(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1192(.a(gate273inter0), .b(s_92), .O(gate273inter1));
  and2  gate1193(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1194(.a(s_92), .O(gate273inter3));
  inv1  gate1195(.a(s_93), .O(gate273inter4));
  nand2 gate1196(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1197(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1198(.a(G642), .O(gate273inter7));
  inv1  gate1199(.a(G794), .O(gate273inter8));
  nand2 gate1200(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1201(.a(s_93), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1202(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1203(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1204(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1625(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1626(.a(gate275inter0), .b(s_154), .O(gate275inter1));
  and2  gate1627(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1628(.a(s_154), .O(gate275inter3));
  inv1  gate1629(.a(s_155), .O(gate275inter4));
  nand2 gate1630(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1631(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1632(.a(G645), .O(gate275inter7));
  inv1  gate1633(.a(G797), .O(gate275inter8));
  nand2 gate1634(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1635(.a(s_155), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1636(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1637(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1638(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2563(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2564(.a(gate278inter0), .b(s_288), .O(gate278inter1));
  and2  gate2565(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2566(.a(s_288), .O(gate278inter3));
  inv1  gate2567(.a(s_289), .O(gate278inter4));
  nand2 gate2568(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2569(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2570(.a(G776), .O(gate278inter7));
  inv1  gate2571(.a(G800), .O(gate278inter8));
  nand2 gate2572(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2573(.a(s_289), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2574(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2575(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2576(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2003(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2004(.a(gate285inter0), .b(s_208), .O(gate285inter1));
  and2  gate2005(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2006(.a(s_208), .O(gate285inter3));
  inv1  gate2007(.a(s_209), .O(gate285inter4));
  nand2 gate2008(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2009(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2010(.a(G660), .O(gate285inter7));
  inv1  gate2011(.a(G812), .O(gate285inter8));
  nand2 gate2012(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2013(.a(s_209), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2014(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2015(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2016(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2871(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2872(.a(gate286inter0), .b(s_332), .O(gate286inter1));
  and2  gate2873(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2874(.a(s_332), .O(gate286inter3));
  inv1  gate2875(.a(s_333), .O(gate286inter4));
  nand2 gate2876(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2877(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2878(.a(G788), .O(gate286inter7));
  inv1  gate2879(.a(G812), .O(gate286inter8));
  nand2 gate2880(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2881(.a(s_333), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2882(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2883(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2884(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate589(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate590(.a(gate287inter0), .b(s_6), .O(gate287inter1));
  and2  gate591(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate592(.a(s_6), .O(gate287inter3));
  inv1  gate593(.a(s_7), .O(gate287inter4));
  nand2 gate594(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate595(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate596(.a(G663), .O(gate287inter7));
  inv1  gate597(.a(G815), .O(gate287inter8));
  nand2 gate598(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate599(.a(s_7), .b(gate287inter3), .O(gate287inter10));
  nor2  gate600(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate601(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate602(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate953(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate954(.a(gate289inter0), .b(s_58), .O(gate289inter1));
  and2  gate955(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate956(.a(s_58), .O(gate289inter3));
  inv1  gate957(.a(s_59), .O(gate289inter4));
  nand2 gate958(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate959(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate960(.a(G818), .O(gate289inter7));
  inv1  gate961(.a(G819), .O(gate289inter8));
  nand2 gate962(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate963(.a(s_59), .b(gate289inter3), .O(gate289inter10));
  nor2  gate964(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate965(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate966(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1653(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1654(.a(gate292inter0), .b(s_158), .O(gate292inter1));
  and2  gate1655(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1656(.a(s_158), .O(gate292inter3));
  inv1  gate1657(.a(s_159), .O(gate292inter4));
  nand2 gate1658(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1659(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1660(.a(G824), .O(gate292inter7));
  inv1  gate1661(.a(G825), .O(gate292inter8));
  nand2 gate1662(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1663(.a(s_159), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1664(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1665(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1666(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2997(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2998(.a(gate294inter0), .b(s_350), .O(gate294inter1));
  and2  gate2999(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate3000(.a(s_350), .O(gate294inter3));
  inv1  gate3001(.a(s_351), .O(gate294inter4));
  nand2 gate3002(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate3003(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate3004(.a(G832), .O(gate294inter7));
  inv1  gate3005(.a(G833), .O(gate294inter8));
  nand2 gate3006(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate3007(.a(s_351), .b(gate294inter3), .O(gate294inter10));
  nor2  gate3008(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate3009(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate3010(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1877(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1878(.a(gate296inter0), .b(s_190), .O(gate296inter1));
  and2  gate1879(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1880(.a(s_190), .O(gate296inter3));
  inv1  gate1881(.a(s_191), .O(gate296inter4));
  nand2 gate1882(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1883(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1884(.a(G826), .O(gate296inter7));
  inv1  gate1885(.a(G827), .O(gate296inter8));
  nand2 gate1886(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1887(.a(s_191), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1888(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1889(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1890(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1975(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1976(.a(gate387inter0), .b(s_204), .O(gate387inter1));
  and2  gate1977(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1978(.a(s_204), .O(gate387inter3));
  inv1  gate1979(.a(s_205), .O(gate387inter4));
  nand2 gate1980(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1981(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1982(.a(G1), .O(gate387inter7));
  inv1  gate1983(.a(G1036), .O(gate387inter8));
  nand2 gate1984(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1985(.a(s_205), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1986(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1987(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1988(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate2941(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2942(.a(gate390inter0), .b(s_342), .O(gate390inter1));
  and2  gate2943(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2944(.a(s_342), .O(gate390inter3));
  inv1  gate2945(.a(s_343), .O(gate390inter4));
  nand2 gate2946(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2947(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2948(.a(G4), .O(gate390inter7));
  inv1  gate2949(.a(G1045), .O(gate390inter8));
  nand2 gate2950(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2951(.a(s_343), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2952(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2953(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2954(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1849(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1850(.a(gate391inter0), .b(s_186), .O(gate391inter1));
  and2  gate1851(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1852(.a(s_186), .O(gate391inter3));
  inv1  gate1853(.a(s_187), .O(gate391inter4));
  nand2 gate1854(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1855(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1856(.a(G5), .O(gate391inter7));
  inv1  gate1857(.a(G1048), .O(gate391inter8));
  nand2 gate1858(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1859(.a(s_187), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1860(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1861(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1862(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2633(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2634(.a(gate394inter0), .b(s_298), .O(gate394inter1));
  and2  gate2635(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2636(.a(s_298), .O(gate394inter3));
  inv1  gate2637(.a(s_299), .O(gate394inter4));
  nand2 gate2638(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2639(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2640(.a(G8), .O(gate394inter7));
  inv1  gate2641(.a(G1057), .O(gate394inter8));
  nand2 gate2642(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2643(.a(s_299), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2644(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2645(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2646(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1079(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1080(.a(gate395inter0), .b(s_76), .O(gate395inter1));
  and2  gate1081(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1082(.a(s_76), .O(gate395inter3));
  inv1  gate1083(.a(s_77), .O(gate395inter4));
  nand2 gate1084(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1085(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1086(.a(G9), .O(gate395inter7));
  inv1  gate1087(.a(G1060), .O(gate395inter8));
  nand2 gate1088(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1089(.a(s_77), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1090(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1091(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1092(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2283(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2284(.a(gate396inter0), .b(s_248), .O(gate396inter1));
  and2  gate2285(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2286(.a(s_248), .O(gate396inter3));
  inv1  gate2287(.a(s_249), .O(gate396inter4));
  nand2 gate2288(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2289(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2290(.a(G10), .O(gate396inter7));
  inv1  gate2291(.a(G1063), .O(gate396inter8));
  nand2 gate2292(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2293(.a(s_249), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2294(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2295(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2296(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate2465(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2466(.a(gate397inter0), .b(s_274), .O(gate397inter1));
  and2  gate2467(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2468(.a(s_274), .O(gate397inter3));
  inv1  gate2469(.a(s_275), .O(gate397inter4));
  nand2 gate2470(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2471(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2472(.a(G11), .O(gate397inter7));
  inv1  gate2473(.a(G1066), .O(gate397inter8));
  nand2 gate2474(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2475(.a(s_275), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2476(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2477(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2478(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2073(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2074(.a(gate398inter0), .b(s_218), .O(gate398inter1));
  and2  gate2075(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2076(.a(s_218), .O(gate398inter3));
  inv1  gate2077(.a(s_219), .O(gate398inter4));
  nand2 gate2078(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2079(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2080(.a(G12), .O(gate398inter7));
  inv1  gate2081(.a(G1069), .O(gate398inter8));
  nand2 gate2082(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2083(.a(s_219), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2084(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2085(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2086(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate2269(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2270(.a(gate399inter0), .b(s_246), .O(gate399inter1));
  and2  gate2271(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2272(.a(s_246), .O(gate399inter3));
  inv1  gate2273(.a(s_247), .O(gate399inter4));
  nand2 gate2274(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2275(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2276(.a(G13), .O(gate399inter7));
  inv1  gate2277(.a(G1072), .O(gate399inter8));
  nand2 gate2278(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2279(.a(s_247), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2280(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2281(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2282(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2829(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2830(.a(gate400inter0), .b(s_326), .O(gate400inter1));
  and2  gate2831(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2832(.a(s_326), .O(gate400inter3));
  inv1  gate2833(.a(s_327), .O(gate400inter4));
  nand2 gate2834(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2835(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2836(.a(G14), .O(gate400inter7));
  inv1  gate2837(.a(G1075), .O(gate400inter8));
  nand2 gate2838(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2839(.a(s_327), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2840(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2841(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2842(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2843(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2844(.a(gate401inter0), .b(s_328), .O(gate401inter1));
  and2  gate2845(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2846(.a(s_328), .O(gate401inter3));
  inv1  gate2847(.a(s_329), .O(gate401inter4));
  nand2 gate2848(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2849(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2850(.a(G15), .O(gate401inter7));
  inv1  gate2851(.a(G1078), .O(gate401inter8));
  nand2 gate2852(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2853(.a(s_329), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2854(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2855(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2856(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2661(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2662(.a(gate404inter0), .b(s_302), .O(gate404inter1));
  and2  gate2663(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2664(.a(s_302), .O(gate404inter3));
  inv1  gate2665(.a(s_303), .O(gate404inter4));
  nand2 gate2666(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2667(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2668(.a(G18), .O(gate404inter7));
  inv1  gate2669(.a(G1087), .O(gate404inter8));
  nand2 gate2670(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2671(.a(s_303), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2672(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2673(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2674(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate2185(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2186(.a(gate405inter0), .b(s_234), .O(gate405inter1));
  and2  gate2187(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2188(.a(s_234), .O(gate405inter3));
  inv1  gate2189(.a(s_235), .O(gate405inter4));
  nand2 gate2190(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2191(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2192(.a(G19), .O(gate405inter7));
  inv1  gate2193(.a(G1090), .O(gate405inter8));
  nand2 gate2194(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2195(.a(s_235), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2196(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2197(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2198(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1345(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1346(.a(gate406inter0), .b(s_114), .O(gate406inter1));
  and2  gate1347(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1348(.a(s_114), .O(gate406inter3));
  inv1  gate1349(.a(s_115), .O(gate406inter4));
  nand2 gate1350(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1351(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1352(.a(G20), .O(gate406inter7));
  inv1  gate1353(.a(G1093), .O(gate406inter8));
  nand2 gate1354(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1355(.a(s_115), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1356(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1357(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1358(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate827(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate828(.a(gate408inter0), .b(s_40), .O(gate408inter1));
  and2  gate829(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate830(.a(s_40), .O(gate408inter3));
  inv1  gate831(.a(s_41), .O(gate408inter4));
  nand2 gate832(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate833(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate834(.a(G22), .O(gate408inter7));
  inv1  gate835(.a(G1099), .O(gate408inter8));
  nand2 gate836(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate837(.a(s_41), .b(gate408inter3), .O(gate408inter10));
  nor2  gate838(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate839(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate840(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate2353(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2354(.a(gate409inter0), .b(s_258), .O(gate409inter1));
  and2  gate2355(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2356(.a(s_258), .O(gate409inter3));
  inv1  gate2357(.a(s_259), .O(gate409inter4));
  nand2 gate2358(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2359(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2360(.a(G23), .O(gate409inter7));
  inv1  gate2361(.a(G1102), .O(gate409inter8));
  nand2 gate2362(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2363(.a(s_259), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2364(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2365(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2366(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1387(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1388(.a(gate413inter0), .b(s_120), .O(gate413inter1));
  and2  gate1389(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1390(.a(s_120), .O(gate413inter3));
  inv1  gate1391(.a(s_121), .O(gate413inter4));
  nand2 gate1392(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1393(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1394(.a(G27), .O(gate413inter7));
  inv1  gate1395(.a(G1114), .O(gate413inter8));
  nand2 gate1396(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1397(.a(s_121), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1398(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1399(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1400(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1793(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1794(.a(gate415inter0), .b(s_178), .O(gate415inter1));
  and2  gate1795(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1796(.a(s_178), .O(gate415inter3));
  inv1  gate1797(.a(s_179), .O(gate415inter4));
  nand2 gate1798(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1799(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1800(.a(G29), .O(gate415inter7));
  inv1  gate1801(.a(G1120), .O(gate415inter8));
  nand2 gate1802(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1803(.a(s_179), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1804(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1805(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1806(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate2885(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2886(.a(gate416inter0), .b(s_334), .O(gate416inter1));
  and2  gate2887(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2888(.a(s_334), .O(gate416inter3));
  inv1  gate2889(.a(s_335), .O(gate416inter4));
  nand2 gate2890(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2891(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2892(.a(G30), .O(gate416inter7));
  inv1  gate2893(.a(G1123), .O(gate416inter8));
  nand2 gate2894(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2895(.a(s_335), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2896(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2897(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2898(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1737(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1738(.a(gate417inter0), .b(s_170), .O(gate417inter1));
  and2  gate1739(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1740(.a(s_170), .O(gate417inter3));
  inv1  gate1741(.a(s_171), .O(gate417inter4));
  nand2 gate1742(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1743(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1744(.a(G31), .O(gate417inter7));
  inv1  gate1745(.a(G1126), .O(gate417inter8));
  nand2 gate1746(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1747(.a(s_171), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1748(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1749(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1750(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate981(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate982(.a(gate418inter0), .b(s_62), .O(gate418inter1));
  and2  gate983(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate984(.a(s_62), .O(gate418inter3));
  inv1  gate985(.a(s_63), .O(gate418inter4));
  nand2 gate986(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate987(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate988(.a(G32), .O(gate418inter7));
  inv1  gate989(.a(G1129), .O(gate418inter8));
  nand2 gate990(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate991(.a(s_63), .b(gate418inter3), .O(gate418inter10));
  nor2  gate992(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate993(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate994(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2213(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2214(.a(gate419inter0), .b(s_238), .O(gate419inter1));
  and2  gate2215(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2216(.a(s_238), .O(gate419inter3));
  inv1  gate2217(.a(s_239), .O(gate419inter4));
  nand2 gate2218(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2219(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2220(.a(G1), .O(gate419inter7));
  inv1  gate2221(.a(G1132), .O(gate419inter8));
  nand2 gate2222(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2223(.a(s_239), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2224(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2225(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2226(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1051(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1052(.a(gate420inter0), .b(s_72), .O(gate420inter1));
  and2  gate1053(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1054(.a(s_72), .O(gate420inter3));
  inv1  gate1055(.a(s_73), .O(gate420inter4));
  nand2 gate1056(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1057(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1058(.a(G1036), .O(gate420inter7));
  inv1  gate1059(.a(G1132), .O(gate420inter8));
  nand2 gate1060(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1061(.a(s_73), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1062(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1063(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1064(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2031(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2032(.a(gate424inter0), .b(s_212), .O(gate424inter1));
  and2  gate2033(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2034(.a(s_212), .O(gate424inter3));
  inv1  gate2035(.a(s_213), .O(gate424inter4));
  nand2 gate2036(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2037(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2038(.a(G1042), .O(gate424inter7));
  inv1  gate2039(.a(G1138), .O(gate424inter8));
  nand2 gate2040(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2041(.a(s_213), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2042(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2043(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2044(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2059(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2060(.a(gate430inter0), .b(s_216), .O(gate430inter1));
  and2  gate2061(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2062(.a(s_216), .O(gate430inter3));
  inv1  gate2063(.a(s_217), .O(gate430inter4));
  nand2 gate2064(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2065(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2066(.a(G1051), .O(gate430inter7));
  inv1  gate2067(.a(G1147), .O(gate430inter8));
  nand2 gate2068(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2069(.a(s_217), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2070(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2071(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2072(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1233(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1234(.a(gate431inter0), .b(s_98), .O(gate431inter1));
  and2  gate1235(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1236(.a(s_98), .O(gate431inter3));
  inv1  gate1237(.a(s_99), .O(gate431inter4));
  nand2 gate1238(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1239(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1240(.a(G7), .O(gate431inter7));
  inv1  gate1241(.a(G1150), .O(gate431inter8));
  nand2 gate1242(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1243(.a(s_99), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1244(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1245(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1246(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate2521(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2522(.a(gate436inter0), .b(s_282), .O(gate436inter1));
  and2  gate2523(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2524(.a(s_282), .O(gate436inter3));
  inv1  gate2525(.a(s_283), .O(gate436inter4));
  nand2 gate2526(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2527(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2528(.a(G1060), .O(gate436inter7));
  inv1  gate2529(.a(G1156), .O(gate436inter8));
  nand2 gate2530(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2531(.a(s_283), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2532(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2533(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2534(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2409(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2410(.a(gate439inter0), .b(s_266), .O(gate439inter1));
  and2  gate2411(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2412(.a(s_266), .O(gate439inter3));
  inv1  gate2413(.a(s_267), .O(gate439inter4));
  nand2 gate2414(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2415(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2416(.a(G11), .O(gate439inter7));
  inv1  gate2417(.a(G1162), .O(gate439inter8));
  nand2 gate2418(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2419(.a(s_267), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2420(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2421(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2422(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2339(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2340(.a(gate442inter0), .b(s_256), .O(gate442inter1));
  and2  gate2341(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2342(.a(s_256), .O(gate442inter3));
  inv1  gate2343(.a(s_257), .O(gate442inter4));
  nand2 gate2344(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2345(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2346(.a(G1069), .O(gate442inter7));
  inv1  gate2347(.a(G1165), .O(gate442inter8));
  nand2 gate2348(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2349(.a(s_257), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2350(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2351(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2352(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1471(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1472(.a(gate444inter0), .b(s_132), .O(gate444inter1));
  and2  gate1473(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1474(.a(s_132), .O(gate444inter3));
  inv1  gate1475(.a(s_133), .O(gate444inter4));
  nand2 gate1476(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1477(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1478(.a(G1072), .O(gate444inter7));
  inv1  gate1479(.a(G1168), .O(gate444inter8));
  nand2 gate1480(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1481(.a(s_133), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1482(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1483(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1484(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate3347(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate3348(.a(gate445inter0), .b(s_400), .O(gate445inter1));
  and2  gate3349(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate3350(.a(s_400), .O(gate445inter3));
  inv1  gate3351(.a(s_401), .O(gate445inter4));
  nand2 gate3352(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate3353(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate3354(.a(G14), .O(gate445inter7));
  inv1  gate3355(.a(G1171), .O(gate445inter8));
  nand2 gate3356(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate3357(.a(s_401), .b(gate445inter3), .O(gate445inter10));
  nor2  gate3358(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate3359(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate3360(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1205(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1206(.a(gate446inter0), .b(s_94), .O(gate446inter1));
  and2  gate1207(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1208(.a(s_94), .O(gate446inter3));
  inv1  gate1209(.a(s_95), .O(gate446inter4));
  nand2 gate1210(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1211(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1212(.a(G1075), .O(gate446inter7));
  inv1  gate1213(.a(G1171), .O(gate446inter8));
  nand2 gate1214(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1215(.a(s_95), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1216(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1217(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1218(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2241(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2242(.a(gate448inter0), .b(s_242), .O(gate448inter1));
  and2  gate2243(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2244(.a(s_242), .O(gate448inter3));
  inv1  gate2245(.a(s_243), .O(gate448inter4));
  nand2 gate2246(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2247(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2248(.a(G1078), .O(gate448inter7));
  inv1  gate2249(.a(G1174), .O(gate448inter8));
  nand2 gate2250(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2251(.a(s_243), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2252(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2253(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2254(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate3263(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate3264(.a(gate449inter0), .b(s_388), .O(gate449inter1));
  and2  gate3265(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate3266(.a(s_388), .O(gate449inter3));
  inv1  gate3267(.a(s_389), .O(gate449inter4));
  nand2 gate3268(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate3269(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate3270(.a(G16), .O(gate449inter7));
  inv1  gate3271(.a(G1177), .O(gate449inter8));
  nand2 gate3272(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate3273(.a(s_389), .b(gate449inter3), .O(gate449inter10));
  nor2  gate3274(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate3275(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate3276(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1695(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1696(.a(gate454inter0), .b(s_164), .O(gate454inter1));
  and2  gate1697(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1698(.a(s_164), .O(gate454inter3));
  inv1  gate1699(.a(s_165), .O(gate454inter4));
  nand2 gate1700(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1701(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1702(.a(G1087), .O(gate454inter7));
  inv1  gate1703(.a(G1183), .O(gate454inter8));
  nand2 gate1704(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1705(.a(s_165), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1706(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1707(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1708(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1835(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1836(.a(gate459inter0), .b(s_184), .O(gate459inter1));
  and2  gate1837(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1838(.a(s_184), .O(gate459inter3));
  inv1  gate1839(.a(s_185), .O(gate459inter4));
  nand2 gate1840(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1841(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1842(.a(G21), .O(gate459inter7));
  inv1  gate1843(.a(G1192), .O(gate459inter8));
  nand2 gate1844(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1845(.a(s_185), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1846(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1847(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1848(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2647(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2648(.a(gate462inter0), .b(s_300), .O(gate462inter1));
  and2  gate2649(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2650(.a(s_300), .O(gate462inter3));
  inv1  gate2651(.a(s_301), .O(gate462inter4));
  nand2 gate2652(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2653(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2654(.a(G1099), .O(gate462inter7));
  inv1  gate2655(.a(G1195), .O(gate462inter8));
  nand2 gate2656(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2657(.a(s_301), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2658(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2659(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2660(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1723(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1724(.a(gate463inter0), .b(s_168), .O(gate463inter1));
  and2  gate1725(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1726(.a(s_168), .O(gate463inter3));
  inv1  gate1727(.a(s_169), .O(gate463inter4));
  nand2 gate1728(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1729(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1730(.a(G23), .O(gate463inter7));
  inv1  gate1731(.a(G1198), .O(gate463inter8));
  nand2 gate1732(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1733(.a(s_169), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1734(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1735(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1736(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate3333(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate3334(.a(gate467inter0), .b(s_398), .O(gate467inter1));
  and2  gate3335(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate3336(.a(s_398), .O(gate467inter3));
  inv1  gate3337(.a(s_399), .O(gate467inter4));
  nand2 gate3338(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate3339(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate3340(.a(G25), .O(gate467inter7));
  inv1  gate3341(.a(G1204), .O(gate467inter8));
  nand2 gate3342(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate3343(.a(s_399), .b(gate467inter3), .O(gate467inter10));
  nor2  gate3344(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate3345(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate3346(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1639(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1640(.a(gate471inter0), .b(s_156), .O(gate471inter1));
  and2  gate1641(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1642(.a(s_156), .O(gate471inter3));
  inv1  gate1643(.a(s_157), .O(gate471inter4));
  nand2 gate1644(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1645(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1646(.a(G27), .O(gate471inter7));
  inv1  gate1647(.a(G1210), .O(gate471inter8));
  nand2 gate1648(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1649(.a(s_157), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1650(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1651(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1652(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate3165(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate3166(.a(gate473inter0), .b(s_374), .O(gate473inter1));
  and2  gate3167(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate3168(.a(s_374), .O(gate473inter3));
  inv1  gate3169(.a(s_375), .O(gate473inter4));
  nand2 gate3170(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate3171(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate3172(.a(G28), .O(gate473inter7));
  inv1  gate3173(.a(G1213), .O(gate473inter8));
  nand2 gate3174(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate3175(.a(s_375), .b(gate473inter3), .O(gate473inter10));
  nor2  gate3176(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate3177(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate3178(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2199(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2200(.a(gate475inter0), .b(s_236), .O(gate475inter1));
  and2  gate2201(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2202(.a(s_236), .O(gate475inter3));
  inv1  gate2203(.a(s_237), .O(gate475inter4));
  nand2 gate2204(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2205(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2206(.a(G29), .O(gate475inter7));
  inv1  gate2207(.a(G1216), .O(gate475inter8));
  nand2 gate2208(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2209(.a(s_237), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2210(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2211(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2212(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2045(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2046(.a(gate477inter0), .b(s_214), .O(gate477inter1));
  and2  gate2047(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2048(.a(s_214), .O(gate477inter3));
  inv1  gate2049(.a(s_215), .O(gate477inter4));
  nand2 gate2050(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2051(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2052(.a(G30), .O(gate477inter7));
  inv1  gate2053(.a(G1219), .O(gate477inter8));
  nand2 gate2054(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2055(.a(s_215), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2056(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2057(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2058(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate3207(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate3208(.a(gate478inter0), .b(s_380), .O(gate478inter1));
  and2  gate3209(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate3210(.a(s_380), .O(gate478inter3));
  inv1  gate3211(.a(s_381), .O(gate478inter4));
  nand2 gate3212(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate3213(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate3214(.a(G1123), .O(gate478inter7));
  inv1  gate3215(.a(G1219), .O(gate478inter8));
  nand2 gate3216(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate3217(.a(s_381), .b(gate478inter3), .O(gate478inter10));
  nor2  gate3218(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate3219(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate3220(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate3067(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate3068(.a(gate480inter0), .b(s_360), .O(gate480inter1));
  and2  gate3069(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate3070(.a(s_360), .O(gate480inter3));
  inv1  gate3071(.a(s_361), .O(gate480inter4));
  nand2 gate3072(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate3073(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate3074(.a(G1126), .O(gate480inter7));
  inv1  gate3075(.a(G1222), .O(gate480inter8));
  nand2 gate3076(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate3077(.a(s_361), .b(gate480inter3), .O(gate480inter10));
  nor2  gate3078(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate3079(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate3080(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate3277(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate3278(.a(gate484inter0), .b(s_390), .O(gate484inter1));
  and2  gate3279(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate3280(.a(s_390), .O(gate484inter3));
  inv1  gate3281(.a(s_391), .O(gate484inter4));
  nand2 gate3282(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate3283(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate3284(.a(G1230), .O(gate484inter7));
  inv1  gate3285(.a(G1231), .O(gate484inter8));
  nand2 gate3286(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate3287(.a(s_391), .b(gate484inter3), .O(gate484inter10));
  nor2  gate3288(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate3289(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate3290(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate603(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate604(.a(gate487inter0), .b(s_8), .O(gate487inter1));
  and2  gate605(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate606(.a(s_8), .O(gate487inter3));
  inv1  gate607(.a(s_9), .O(gate487inter4));
  nand2 gate608(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate609(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate610(.a(G1236), .O(gate487inter7));
  inv1  gate611(.a(G1237), .O(gate487inter8));
  nand2 gate612(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate613(.a(s_9), .b(gate487inter3), .O(gate487inter10));
  nor2  gate614(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate615(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate616(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1807(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1808(.a(gate489inter0), .b(s_180), .O(gate489inter1));
  and2  gate1809(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1810(.a(s_180), .O(gate489inter3));
  inv1  gate1811(.a(s_181), .O(gate489inter4));
  nand2 gate1812(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1813(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1814(.a(G1240), .O(gate489inter7));
  inv1  gate1815(.a(G1241), .O(gate489inter8));
  nand2 gate1816(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1817(.a(s_181), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1818(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1819(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1820(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2619(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2620(.a(gate493inter0), .b(s_296), .O(gate493inter1));
  and2  gate2621(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2622(.a(s_296), .O(gate493inter3));
  inv1  gate2623(.a(s_297), .O(gate493inter4));
  nand2 gate2624(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2625(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2626(.a(G1248), .O(gate493inter7));
  inv1  gate2627(.a(G1249), .O(gate493inter8));
  nand2 gate2628(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2629(.a(s_297), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2630(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2631(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2632(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate3319(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate3320(.a(gate494inter0), .b(s_396), .O(gate494inter1));
  and2  gate3321(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate3322(.a(s_396), .O(gate494inter3));
  inv1  gate3323(.a(s_397), .O(gate494inter4));
  nand2 gate3324(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate3325(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate3326(.a(G1250), .O(gate494inter7));
  inv1  gate3327(.a(G1251), .O(gate494inter8));
  nand2 gate3328(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate3329(.a(s_397), .b(gate494inter3), .O(gate494inter10));
  nor2  gate3330(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate3331(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate3332(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate2087(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2088(.a(gate498inter0), .b(s_220), .O(gate498inter1));
  and2  gate2089(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2090(.a(s_220), .O(gate498inter3));
  inv1  gate2091(.a(s_221), .O(gate498inter4));
  nand2 gate2092(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2093(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2094(.a(G1258), .O(gate498inter7));
  inv1  gate2095(.a(G1259), .O(gate498inter8));
  nand2 gate2096(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2097(.a(s_221), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2098(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2099(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2100(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate3025(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate3026(.a(gate501inter0), .b(s_354), .O(gate501inter1));
  and2  gate3027(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate3028(.a(s_354), .O(gate501inter3));
  inv1  gate3029(.a(s_355), .O(gate501inter4));
  nand2 gate3030(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate3031(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate3032(.a(G1264), .O(gate501inter7));
  inv1  gate3033(.a(G1265), .O(gate501inter8));
  nand2 gate3034(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate3035(.a(s_355), .b(gate501inter3), .O(gate501inter10));
  nor2  gate3036(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate3037(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate3038(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate813(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate814(.a(gate502inter0), .b(s_38), .O(gate502inter1));
  and2  gate815(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate816(.a(s_38), .O(gate502inter3));
  inv1  gate817(.a(s_39), .O(gate502inter4));
  nand2 gate818(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate819(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate820(.a(G1266), .O(gate502inter7));
  inv1  gate821(.a(G1267), .O(gate502inter8));
  nand2 gate822(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate823(.a(s_39), .b(gate502inter3), .O(gate502inter10));
  nor2  gate824(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate825(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate826(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1163(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1164(.a(gate504inter0), .b(s_88), .O(gate504inter1));
  and2  gate1165(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1166(.a(s_88), .O(gate504inter3));
  inv1  gate1167(.a(s_89), .O(gate504inter4));
  nand2 gate1168(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1169(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1170(.a(G1270), .O(gate504inter7));
  inv1  gate1171(.a(G1271), .O(gate504inter8));
  nand2 gate1172(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1173(.a(s_89), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1174(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1175(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1176(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate3011(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate3012(.a(gate506inter0), .b(s_352), .O(gate506inter1));
  and2  gate3013(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate3014(.a(s_352), .O(gate506inter3));
  inv1  gate3015(.a(s_353), .O(gate506inter4));
  nand2 gate3016(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate3017(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate3018(.a(G1274), .O(gate506inter7));
  inv1  gate3019(.a(G1275), .O(gate506inter8));
  nand2 gate3020(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate3021(.a(s_353), .b(gate506inter3), .O(gate506inter10));
  nor2  gate3022(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate3023(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate3024(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2801(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2802(.a(gate509inter0), .b(s_322), .O(gate509inter1));
  and2  gate2803(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2804(.a(s_322), .O(gate509inter3));
  inv1  gate2805(.a(s_323), .O(gate509inter4));
  nand2 gate2806(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2807(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2808(.a(G1280), .O(gate509inter7));
  inv1  gate2809(.a(G1281), .O(gate509inter8));
  nand2 gate2810(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2811(.a(s_323), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2812(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2813(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2814(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1583(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1584(.a(gate512inter0), .b(s_148), .O(gate512inter1));
  and2  gate1585(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1586(.a(s_148), .O(gate512inter3));
  inv1  gate1587(.a(s_149), .O(gate512inter4));
  nand2 gate1588(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1589(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1590(.a(G1286), .O(gate512inter7));
  inv1  gate1591(.a(G1287), .O(gate512inter8));
  nand2 gate1592(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1593(.a(s_149), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1594(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1595(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1596(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2955(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2956(.a(gate514inter0), .b(s_344), .O(gate514inter1));
  and2  gate2957(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2958(.a(s_344), .O(gate514inter3));
  inv1  gate2959(.a(s_345), .O(gate514inter4));
  nand2 gate2960(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2961(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2962(.a(G1290), .O(gate514inter7));
  inv1  gate2963(.a(G1291), .O(gate514inter8));
  nand2 gate2964(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2965(.a(s_345), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2966(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2967(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2968(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule