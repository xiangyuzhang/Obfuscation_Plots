module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate701(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate702(.a(gate14inter0), .b(s_22), .O(gate14inter1));
  and2  gate703(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate704(.a(s_22), .O(gate14inter3));
  inv1  gate705(.a(s_23), .O(gate14inter4));
  nand2 gate706(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate707(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate708(.a(G11), .O(gate14inter7));
  inv1  gate709(.a(G12), .O(gate14inter8));
  nand2 gate710(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate711(.a(s_23), .b(gate14inter3), .O(gate14inter10));
  nor2  gate712(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate713(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate714(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate897(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate898(.a(gate16inter0), .b(s_50), .O(gate16inter1));
  and2  gate899(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate900(.a(s_50), .O(gate16inter3));
  inv1  gate901(.a(s_51), .O(gate16inter4));
  nand2 gate902(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate903(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate904(.a(G15), .O(gate16inter7));
  inv1  gate905(.a(G16), .O(gate16inter8));
  nand2 gate906(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate907(.a(s_51), .b(gate16inter3), .O(gate16inter10));
  nor2  gate908(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate909(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate910(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1163(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1164(.a(gate17inter0), .b(s_88), .O(gate17inter1));
  and2  gate1165(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1166(.a(s_88), .O(gate17inter3));
  inv1  gate1167(.a(s_89), .O(gate17inter4));
  nand2 gate1168(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1169(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1170(.a(G17), .O(gate17inter7));
  inv1  gate1171(.a(G18), .O(gate17inter8));
  nand2 gate1172(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1173(.a(s_89), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1174(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1175(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1176(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1219(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1220(.a(gate25inter0), .b(s_96), .O(gate25inter1));
  and2  gate1221(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1222(.a(s_96), .O(gate25inter3));
  inv1  gate1223(.a(s_97), .O(gate25inter4));
  nand2 gate1224(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1225(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1226(.a(G1), .O(gate25inter7));
  inv1  gate1227(.a(G5), .O(gate25inter8));
  nand2 gate1228(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1229(.a(s_97), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1230(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1231(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1232(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate659(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate660(.a(gate27inter0), .b(s_16), .O(gate27inter1));
  and2  gate661(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate662(.a(s_16), .O(gate27inter3));
  inv1  gate663(.a(s_17), .O(gate27inter4));
  nand2 gate664(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate665(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate666(.a(G2), .O(gate27inter7));
  inv1  gate667(.a(G6), .O(gate27inter8));
  nand2 gate668(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate669(.a(s_17), .b(gate27inter3), .O(gate27inter10));
  nor2  gate670(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate671(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate672(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate561(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate562(.a(gate29inter0), .b(s_2), .O(gate29inter1));
  and2  gate563(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate564(.a(s_2), .O(gate29inter3));
  inv1  gate565(.a(s_3), .O(gate29inter4));
  nand2 gate566(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate567(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate568(.a(G3), .O(gate29inter7));
  inv1  gate569(.a(G7), .O(gate29inter8));
  nand2 gate570(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate571(.a(s_3), .b(gate29inter3), .O(gate29inter10));
  nor2  gate572(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate573(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate574(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1639(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1640(.a(gate31inter0), .b(s_156), .O(gate31inter1));
  and2  gate1641(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1642(.a(s_156), .O(gate31inter3));
  inv1  gate1643(.a(s_157), .O(gate31inter4));
  nand2 gate1644(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1645(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1646(.a(G4), .O(gate31inter7));
  inv1  gate1647(.a(G8), .O(gate31inter8));
  nand2 gate1648(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1649(.a(s_157), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1650(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1651(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1652(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate953(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate954(.a(gate41inter0), .b(s_58), .O(gate41inter1));
  and2  gate955(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate956(.a(s_58), .O(gate41inter3));
  inv1  gate957(.a(s_59), .O(gate41inter4));
  nand2 gate958(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate959(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate960(.a(G1), .O(gate41inter7));
  inv1  gate961(.a(G266), .O(gate41inter8));
  nand2 gate962(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate963(.a(s_59), .b(gate41inter3), .O(gate41inter10));
  nor2  gate964(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate965(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate966(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1863(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1864(.a(gate44inter0), .b(s_188), .O(gate44inter1));
  and2  gate1865(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1866(.a(s_188), .O(gate44inter3));
  inv1  gate1867(.a(s_189), .O(gate44inter4));
  nand2 gate1868(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1869(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1870(.a(G4), .O(gate44inter7));
  inv1  gate1871(.a(G269), .O(gate44inter8));
  nand2 gate1872(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1873(.a(s_189), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1874(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1875(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1876(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1289(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1290(.a(gate55inter0), .b(s_106), .O(gate55inter1));
  and2  gate1291(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1292(.a(s_106), .O(gate55inter3));
  inv1  gate1293(.a(s_107), .O(gate55inter4));
  nand2 gate1294(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1295(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1296(.a(G15), .O(gate55inter7));
  inv1  gate1297(.a(G287), .O(gate55inter8));
  nand2 gate1298(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1299(.a(s_107), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1300(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1301(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1302(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate911(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate912(.a(gate56inter0), .b(s_52), .O(gate56inter1));
  and2  gate913(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate914(.a(s_52), .O(gate56inter3));
  inv1  gate915(.a(s_53), .O(gate56inter4));
  nand2 gate916(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate917(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate918(.a(G16), .O(gate56inter7));
  inv1  gate919(.a(G287), .O(gate56inter8));
  nand2 gate920(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate921(.a(s_53), .b(gate56inter3), .O(gate56inter10));
  nor2  gate922(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate923(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate924(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1023(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1024(.a(gate59inter0), .b(s_68), .O(gate59inter1));
  and2  gate1025(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1026(.a(s_68), .O(gate59inter3));
  inv1  gate1027(.a(s_69), .O(gate59inter4));
  nand2 gate1028(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1029(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1030(.a(G19), .O(gate59inter7));
  inv1  gate1031(.a(G293), .O(gate59inter8));
  nand2 gate1032(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1033(.a(s_69), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1034(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1035(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1036(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1527(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1528(.a(gate61inter0), .b(s_140), .O(gate61inter1));
  and2  gate1529(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1530(.a(s_140), .O(gate61inter3));
  inv1  gate1531(.a(s_141), .O(gate61inter4));
  nand2 gate1532(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1533(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1534(.a(G21), .O(gate61inter7));
  inv1  gate1535(.a(G296), .O(gate61inter8));
  nand2 gate1536(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1537(.a(s_141), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1538(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1539(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1540(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate855(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate856(.a(gate63inter0), .b(s_44), .O(gate63inter1));
  and2  gate857(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate858(.a(s_44), .O(gate63inter3));
  inv1  gate859(.a(s_45), .O(gate63inter4));
  nand2 gate860(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate861(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate862(.a(G23), .O(gate63inter7));
  inv1  gate863(.a(G299), .O(gate63inter8));
  nand2 gate864(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate865(.a(s_45), .b(gate63inter3), .O(gate63inter10));
  nor2  gate866(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate867(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate868(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate645(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate646(.a(gate65inter0), .b(s_14), .O(gate65inter1));
  and2  gate647(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate648(.a(s_14), .O(gate65inter3));
  inv1  gate649(.a(s_15), .O(gate65inter4));
  nand2 gate650(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate651(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate652(.a(G25), .O(gate65inter7));
  inv1  gate653(.a(G302), .O(gate65inter8));
  nand2 gate654(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate655(.a(s_15), .b(gate65inter3), .O(gate65inter10));
  nor2  gate656(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate657(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate658(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1037(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1038(.a(gate67inter0), .b(s_70), .O(gate67inter1));
  and2  gate1039(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1040(.a(s_70), .O(gate67inter3));
  inv1  gate1041(.a(s_71), .O(gate67inter4));
  nand2 gate1042(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1043(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1044(.a(G27), .O(gate67inter7));
  inv1  gate1045(.a(G305), .O(gate67inter8));
  nand2 gate1046(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1047(.a(s_71), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1048(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1049(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1050(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1415(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1416(.a(gate69inter0), .b(s_124), .O(gate69inter1));
  and2  gate1417(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1418(.a(s_124), .O(gate69inter3));
  inv1  gate1419(.a(s_125), .O(gate69inter4));
  nand2 gate1420(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1421(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1422(.a(G29), .O(gate69inter7));
  inv1  gate1423(.a(G308), .O(gate69inter8));
  nand2 gate1424(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1425(.a(s_125), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1426(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1427(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1428(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate631(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate632(.a(gate75inter0), .b(s_12), .O(gate75inter1));
  and2  gate633(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate634(.a(s_12), .O(gate75inter3));
  inv1  gate635(.a(s_13), .O(gate75inter4));
  nand2 gate636(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate637(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate638(.a(G9), .O(gate75inter7));
  inv1  gate639(.a(G317), .O(gate75inter8));
  nand2 gate640(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate641(.a(s_13), .b(gate75inter3), .O(gate75inter10));
  nor2  gate642(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate643(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate644(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1471(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1472(.a(gate81inter0), .b(s_132), .O(gate81inter1));
  and2  gate1473(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1474(.a(s_132), .O(gate81inter3));
  inv1  gate1475(.a(s_133), .O(gate81inter4));
  nand2 gate1476(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1477(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1478(.a(G3), .O(gate81inter7));
  inv1  gate1479(.a(G326), .O(gate81inter8));
  nand2 gate1480(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1481(.a(s_133), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1482(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1483(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1484(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1807(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1808(.a(gate83inter0), .b(s_180), .O(gate83inter1));
  and2  gate1809(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1810(.a(s_180), .O(gate83inter3));
  inv1  gate1811(.a(s_181), .O(gate83inter4));
  nand2 gate1812(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1813(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1814(.a(G11), .O(gate83inter7));
  inv1  gate1815(.a(G329), .O(gate83inter8));
  nand2 gate1816(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1817(.a(s_181), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1818(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1819(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1820(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1359(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1360(.a(gate93inter0), .b(s_116), .O(gate93inter1));
  and2  gate1361(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1362(.a(s_116), .O(gate93inter3));
  inv1  gate1363(.a(s_117), .O(gate93inter4));
  nand2 gate1364(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1365(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1366(.a(G18), .O(gate93inter7));
  inv1  gate1367(.a(G344), .O(gate93inter8));
  nand2 gate1368(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1369(.a(s_117), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1370(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1371(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1372(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1009(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1010(.a(gate95inter0), .b(s_66), .O(gate95inter1));
  and2  gate1011(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1012(.a(s_66), .O(gate95inter3));
  inv1  gate1013(.a(s_67), .O(gate95inter4));
  nand2 gate1014(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1015(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1016(.a(G26), .O(gate95inter7));
  inv1  gate1017(.a(G347), .O(gate95inter8));
  nand2 gate1018(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1019(.a(s_67), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1020(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1021(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1022(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate925(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate926(.a(gate98inter0), .b(s_54), .O(gate98inter1));
  and2  gate927(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate928(.a(s_54), .O(gate98inter3));
  inv1  gate929(.a(s_55), .O(gate98inter4));
  nand2 gate930(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate931(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate932(.a(G23), .O(gate98inter7));
  inv1  gate933(.a(G350), .O(gate98inter8));
  nand2 gate934(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate935(.a(s_55), .b(gate98inter3), .O(gate98inter10));
  nor2  gate936(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate937(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate938(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1513(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1514(.a(gate100inter0), .b(s_138), .O(gate100inter1));
  and2  gate1515(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1516(.a(s_138), .O(gate100inter3));
  inv1  gate1517(.a(s_139), .O(gate100inter4));
  nand2 gate1518(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1519(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1520(.a(G31), .O(gate100inter7));
  inv1  gate1521(.a(G353), .O(gate100inter8));
  nand2 gate1522(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1523(.a(s_139), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1524(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1525(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1526(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1681(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1682(.a(gate107inter0), .b(s_162), .O(gate107inter1));
  and2  gate1683(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1684(.a(s_162), .O(gate107inter3));
  inv1  gate1685(.a(s_163), .O(gate107inter4));
  nand2 gate1686(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1687(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1688(.a(G366), .O(gate107inter7));
  inv1  gate1689(.a(G367), .O(gate107inter8));
  nand2 gate1690(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1691(.a(s_163), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1692(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1693(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1694(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate785(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate786(.a(gate109inter0), .b(s_34), .O(gate109inter1));
  and2  gate787(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate788(.a(s_34), .O(gate109inter3));
  inv1  gate789(.a(s_35), .O(gate109inter4));
  nand2 gate790(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate791(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate792(.a(G370), .O(gate109inter7));
  inv1  gate793(.a(G371), .O(gate109inter8));
  nand2 gate794(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate795(.a(s_35), .b(gate109inter3), .O(gate109inter10));
  nor2  gate796(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate797(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate798(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1177(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1178(.a(gate118inter0), .b(s_90), .O(gate118inter1));
  and2  gate1179(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1180(.a(s_90), .O(gate118inter3));
  inv1  gate1181(.a(s_91), .O(gate118inter4));
  nand2 gate1182(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1183(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1184(.a(G388), .O(gate118inter7));
  inv1  gate1185(.a(G389), .O(gate118inter8));
  nand2 gate1186(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1187(.a(s_91), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1188(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1189(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1190(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1093(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1094(.a(gate121inter0), .b(s_78), .O(gate121inter1));
  and2  gate1095(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1096(.a(s_78), .O(gate121inter3));
  inv1  gate1097(.a(s_79), .O(gate121inter4));
  nand2 gate1098(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1099(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1100(.a(G394), .O(gate121inter7));
  inv1  gate1101(.a(G395), .O(gate121inter8));
  nand2 gate1102(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1103(.a(s_79), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1104(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1105(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1106(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1303(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1304(.a(gate128inter0), .b(s_108), .O(gate128inter1));
  and2  gate1305(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1306(.a(s_108), .O(gate128inter3));
  inv1  gate1307(.a(s_109), .O(gate128inter4));
  nand2 gate1308(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1309(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1310(.a(G408), .O(gate128inter7));
  inv1  gate1311(.a(G409), .O(gate128inter8));
  nand2 gate1312(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1313(.a(s_109), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1314(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1315(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1316(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1135(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1136(.a(gate136inter0), .b(s_84), .O(gate136inter1));
  and2  gate1137(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1138(.a(s_84), .O(gate136inter3));
  inv1  gate1139(.a(s_85), .O(gate136inter4));
  nand2 gate1140(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1141(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1142(.a(G424), .O(gate136inter7));
  inv1  gate1143(.a(G425), .O(gate136inter8));
  nand2 gate1144(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1145(.a(s_85), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1146(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1147(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1148(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1107(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1108(.a(gate137inter0), .b(s_80), .O(gate137inter1));
  and2  gate1109(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1110(.a(s_80), .O(gate137inter3));
  inv1  gate1111(.a(s_81), .O(gate137inter4));
  nand2 gate1112(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1113(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1114(.a(G426), .O(gate137inter7));
  inv1  gate1115(.a(G429), .O(gate137inter8));
  nand2 gate1116(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1117(.a(s_81), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1118(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1119(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1120(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1191(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1192(.a(gate139inter0), .b(s_92), .O(gate139inter1));
  and2  gate1193(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1194(.a(s_92), .O(gate139inter3));
  inv1  gate1195(.a(s_93), .O(gate139inter4));
  nand2 gate1196(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1197(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1198(.a(G438), .O(gate139inter7));
  inv1  gate1199(.a(G441), .O(gate139inter8));
  nand2 gate1200(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1201(.a(s_93), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1202(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1203(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1204(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1149(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1150(.a(gate142inter0), .b(s_86), .O(gate142inter1));
  and2  gate1151(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1152(.a(s_86), .O(gate142inter3));
  inv1  gate1153(.a(s_87), .O(gate142inter4));
  nand2 gate1154(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1155(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1156(.a(G456), .O(gate142inter7));
  inv1  gate1157(.a(G459), .O(gate142inter8));
  nand2 gate1158(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1159(.a(s_87), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1160(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1161(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1162(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1457(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1458(.a(gate147inter0), .b(s_130), .O(gate147inter1));
  and2  gate1459(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1460(.a(s_130), .O(gate147inter3));
  inv1  gate1461(.a(s_131), .O(gate147inter4));
  nand2 gate1462(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1463(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1464(.a(G486), .O(gate147inter7));
  inv1  gate1465(.a(G489), .O(gate147inter8));
  nand2 gate1466(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1467(.a(s_131), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1468(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1469(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1470(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1723(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1724(.a(gate149inter0), .b(s_168), .O(gate149inter1));
  and2  gate1725(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1726(.a(s_168), .O(gate149inter3));
  inv1  gate1727(.a(s_169), .O(gate149inter4));
  nand2 gate1728(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1729(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1730(.a(G498), .O(gate149inter7));
  inv1  gate1731(.a(G501), .O(gate149inter8));
  nand2 gate1732(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1733(.a(s_169), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1734(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1735(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1736(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1779(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1780(.a(gate150inter0), .b(s_176), .O(gate150inter1));
  and2  gate1781(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1782(.a(s_176), .O(gate150inter3));
  inv1  gate1783(.a(s_177), .O(gate150inter4));
  nand2 gate1784(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1785(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1786(.a(G504), .O(gate150inter7));
  inv1  gate1787(.a(G507), .O(gate150inter8));
  nand2 gate1788(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1789(.a(s_177), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1790(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1791(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1792(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1205(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1206(.a(gate151inter0), .b(s_94), .O(gate151inter1));
  and2  gate1207(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1208(.a(s_94), .O(gate151inter3));
  inv1  gate1209(.a(s_95), .O(gate151inter4));
  nand2 gate1210(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1211(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1212(.a(G510), .O(gate151inter7));
  inv1  gate1213(.a(G513), .O(gate151inter8));
  nand2 gate1214(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1215(.a(s_95), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1216(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1217(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1218(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate981(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate982(.a(gate152inter0), .b(s_62), .O(gate152inter1));
  and2  gate983(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate984(.a(s_62), .O(gate152inter3));
  inv1  gate985(.a(s_63), .O(gate152inter4));
  nand2 gate986(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate987(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate988(.a(G516), .O(gate152inter7));
  inv1  gate989(.a(G519), .O(gate152inter8));
  nand2 gate990(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate991(.a(s_63), .b(gate152inter3), .O(gate152inter10));
  nor2  gate992(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate993(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate994(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1387(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1388(.a(gate160inter0), .b(s_120), .O(gate160inter1));
  and2  gate1389(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1390(.a(s_120), .O(gate160inter3));
  inv1  gate1391(.a(s_121), .O(gate160inter4));
  nand2 gate1392(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1393(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1394(.a(G447), .O(gate160inter7));
  inv1  gate1395(.a(G531), .O(gate160inter8));
  nand2 gate1396(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1397(.a(s_121), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1398(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1399(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1400(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate575(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate576(.a(gate163inter0), .b(s_4), .O(gate163inter1));
  and2  gate577(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate578(.a(s_4), .O(gate163inter3));
  inv1  gate579(.a(s_5), .O(gate163inter4));
  nand2 gate580(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate581(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate582(.a(G456), .O(gate163inter7));
  inv1  gate583(.a(G537), .O(gate163inter8));
  nand2 gate584(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate585(.a(s_5), .b(gate163inter3), .O(gate163inter10));
  nor2  gate586(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate587(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate588(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1275(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1276(.a(gate166inter0), .b(s_104), .O(gate166inter1));
  and2  gate1277(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1278(.a(s_104), .O(gate166inter3));
  inv1  gate1279(.a(s_105), .O(gate166inter4));
  nand2 gate1280(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1281(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1282(.a(G465), .O(gate166inter7));
  inv1  gate1283(.a(G540), .O(gate166inter8));
  nand2 gate1284(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1285(.a(s_105), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1286(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1287(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1288(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1695(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1696(.a(gate175inter0), .b(s_164), .O(gate175inter1));
  and2  gate1697(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1698(.a(s_164), .O(gate175inter3));
  inv1  gate1699(.a(s_165), .O(gate175inter4));
  nand2 gate1700(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1701(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1702(.a(G492), .O(gate175inter7));
  inv1  gate1703(.a(G555), .O(gate175inter8));
  nand2 gate1704(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1705(.a(s_165), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1706(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1707(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1708(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1345(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1346(.a(gate179inter0), .b(s_114), .O(gate179inter1));
  and2  gate1347(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1348(.a(s_114), .O(gate179inter3));
  inv1  gate1349(.a(s_115), .O(gate179inter4));
  nand2 gate1350(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1351(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1352(.a(G504), .O(gate179inter7));
  inv1  gate1353(.a(G561), .O(gate179inter8));
  nand2 gate1354(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1355(.a(s_115), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1356(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1357(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1358(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate687(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate688(.a(gate181inter0), .b(s_20), .O(gate181inter1));
  and2  gate689(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate690(.a(s_20), .O(gate181inter3));
  inv1  gate691(.a(s_21), .O(gate181inter4));
  nand2 gate692(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate693(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate694(.a(G510), .O(gate181inter7));
  inv1  gate695(.a(G564), .O(gate181inter8));
  nand2 gate696(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate697(.a(s_21), .b(gate181inter3), .O(gate181inter10));
  nor2  gate698(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate699(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate700(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate813(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate814(.a(gate182inter0), .b(s_38), .O(gate182inter1));
  and2  gate815(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate816(.a(s_38), .O(gate182inter3));
  inv1  gate817(.a(s_39), .O(gate182inter4));
  nand2 gate818(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate819(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate820(.a(G513), .O(gate182inter7));
  inv1  gate821(.a(G564), .O(gate182inter8));
  nand2 gate822(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate823(.a(s_39), .b(gate182inter3), .O(gate182inter10));
  nor2  gate824(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate825(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate826(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1877(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1878(.a(gate199inter0), .b(s_190), .O(gate199inter1));
  and2  gate1879(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1880(.a(s_190), .O(gate199inter3));
  inv1  gate1881(.a(s_191), .O(gate199inter4));
  nand2 gate1882(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1883(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1884(.a(G598), .O(gate199inter7));
  inv1  gate1885(.a(G599), .O(gate199inter8));
  nand2 gate1886(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1887(.a(s_191), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1888(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1889(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1890(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1611(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1612(.a(gate202inter0), .b(s_152), .O(gate202inter1));
  and2  gate1613(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1614(.a(s_152), .O(gate202inter3));
  inv1  gate1615(.a(s_153), .O(gate202inter4));
  nand2 gate1616(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1617(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1618(.a(G612), .O(gate202inter7));
  inv1  gate1619(.a(G617), .O(gate202inter8));
  nand2 gate1620(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1621(.a(s_153), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1622(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1623(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1624(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate617(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate618(.a(gate203inter0), .b(s_10), .O(gate203inter1));
  and2  gate619(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate620(.a(s_10), .O(gate203inter3));
  inv1  gate621(.a(s_11), .O(gate203inter4));
  nand2 gate622(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate623(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate624(.a(G602), .O(gate203inter7));
  inv1  gate625(.a(G612), .O(gate203inter8));
  nand2 gate626(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate627(.a(s_11), .b(gate203inter3), .O(gate203inter10));
  nor2  gate628(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate629(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate630(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate939(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate940(.a(gate210inter0), .b(s_56), .O(gate210inter1));
  and2  gate941(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate942(.a(s_56), .O(gate210inter3));
  inv1  gate943(.a(s_57), .O(gate210inter4));
  nand2 gate944(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate945(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate946(.a(G607), .O(gate210inter7));
  inv1  gate947(.a(G666), .O(gate210inter8));
  nand2 gate948(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate949(.a(s_57), .b(gate210inter3), .O(gate210inter10));
  nor2  gate950(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate951(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate952(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1429(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1430(.a(gate213inter0), .b(s_126), .O(gate213inter1));
  and2  gate1431(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1432(.a(s_126), .O(gate213inter3));
  inv1  gate1433(.a(s_127), .O(gate213inter4));
  nand2 gate1434(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1435(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1436(.a(G602), .O(gate213inter7));
  inv1  gate1437(.a(G672), .O(gate213inter8));
  nand2 gate1438(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1439(.a(s_127), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1440(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1441(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1442(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate995(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate996(.a(gate214inter0), .b(s_64), .O(gate214inter1));
  and2  gate997(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate998(.a(s_64), .O(gate214inter3));
  inv1  gate999(.a(s_65), .O(gate214inter4));
  nand2 gate1000(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1001(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1002(.a(G612), .O(gate214inter7));
  inv1  gate1003(.a(G672), .O(gate214inter8));
  nand2 gate1004(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1005(.a(s_65), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1006(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1007(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1008(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1821(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1822(.a(gate219inter0), .b(s_182), .O(gate219inter1));
  and2  gate1823(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1824(.a(s_182), .O(gate219inter3));
  inv1  gate1825(.a(s_183), .O(gate219inter4));
  nand2 gate1826(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1827(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1828(.a(G632), .O(gate219inter7));
  inv1  gate1829(.a(G681), .O(gate219inter8));
  nand2 gate1830(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1831(.a(s_183), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1832(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1833(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1834(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate715(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate716(.a(gate220inter0), .b(s_24), .O(gate220inter1));
  and2  gate717(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate718(.a(s_24), .O(gate220inter3));
  inv1  gate719(.a(s_25), .O(gate220inter4));
  nand2 gate720(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate721(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate722(.a(G637), .O(gate220inter7));
  inv1  gate723(.a(G681), .O(gate220inter8));
  nand2 gate724(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate725(.a(s_25), .b(gate220inter3), .O(gate220inter10));
  nor2  gate726(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate727(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate728(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1401(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1402(.a(gate223inter0), .b(s_122), .O(gate223inter1));
  and2  gate1403(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1404(.a(s_122), .O(gate223inter3));
  inv1  gate1405(.a(s_123), .O(gate223inter4));
  nand2 gate1406(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1407(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1408(.a(G627), .O(gate223inter7));
  inv1  gate1409(.a(G687), .O(gate223inter8));
  nand2 gate1410(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1411(.a(s_123), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1412(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1413(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1414(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1065(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1066(.a(gate225inter0), .b(s_74), .O(gate225inter1));
  and2  gate1067(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1068(.a(s_74), .O(gate225inter3));
  inv1  gate1069(.a(s_75), .O(gate225inter4));
  nand2 gate1070(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1071(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1072(.a(G690), .O(gate225inter7));
  inv1  gate1073(.a(G691), .O(gate225inter8));
  nand2 gate1074(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1075(.a(s_75), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1076(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1077(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1078(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1653(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1654(.a(gate233inter0), .b(s_158), .O(gate233inter1));
  and2  gate1655(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1656(.a(s_158), .O(gate233inter3));
  inv1  gate1657(.a(s_159), .O(gate233inter4));
  nand2 gate1658(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1659(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1660(.a(G242), .O(gate233inter7));
  inv1  gate1661(.a(G718), .O(gate233inter8));
  nand2 gate1662(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1663(.a(s_159), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1664(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1665(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1666(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1793(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1794(.a(gate234inter0), .b(s_178), .O(gate234inter1));
  and2  gate1795(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1796(.a(s_178), .O(gate234inter3));
  inv1  gate1797(.a(s_179), .O(gate234inter4));
  nand2 gate1798(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1799(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1800(.a(G245), .O(gate234inter7));
  inv1  gate1801(.a(G721), .O(gate234inter8));
  nand2 gate1802(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1803(.a(s_179), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1804(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1805(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1806(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1849(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1850(.a(gate241inter0), .b(s_186), .O(gate241inter1));
  and2  gate1851(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1852(.a(s_186), .O(gate241inter3));
  inv1  gate1853(.a(s_187), .O(gate241inter4));
  nand2 gate1854(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1855(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1856(.a(G242), .O(gate241inter7));
  inv1  gate1857(.a(G730), .O(gate241inter8));
  nand2 gate1858(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1859(.a(s_187), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1860(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1861(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1862(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1835(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1836(.a(gate249inter0), .b(s_184), .O(gate249inter1));
  and2  gate1837(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1838(.a(s_184), .O(gate249inter3));
  inv1  gate1839(.a(s_185), .O(gate249inter4));
  nand2 gate1840(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1841(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1842(.a(G254), .O(gate249inter7));
  inv1  gate1843(.a(G742), .O(gate249inter8));
  nand2 gate1844(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1845(.a(s_185), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1846(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1847(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1848(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1121(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1122(.a(gate256inter0), .b(s_82), .O(gate256inter1));
  and2  gate1123(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1124(.a(s_82), .O(gate256inter3));
  inv1  gate1125(.a(s_83), .O(gate256inter4));
  nand2 gate1126(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1127(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1128(.a(G715), .O(gate256inter7));
  inv1  gate1129(.a(G751), .O(gate256inter8));
  nand2 gate1130(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1131(.a(s_83), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1132(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1133(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1134(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1051(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1052(.a(gate257inter0), .b(s_72), .O(gate257inter1));
  and2  gate1053(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1054(.a(s_72), .O(gate257inter3));
  inv1  gate1055(.a(s_73), .O(gate257inter4));
  nand2 gate1056(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1057(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1058(.a(G754), .O(gate257inter7));
  inv1  gate1059(.a(G755), .O(gate257inter8));
  nand2 gate1060(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1061(.a(s_73), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1062(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1063(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1064(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1331(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1332(.a(gate259inter0), .b(s_112), .O(gate259inter1));
  and2  gate1333(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1334(.a(s_112), .O(gate259inter3));
  inv1  gate1335(.a(s_113), .O(gate259inter4));
  nand2 gate1336(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1337(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1338(.a(G758), .O(gate259inter7));
  inv1  gate1339(.a(G759), .O(gate259inter8));
  nand2 gate1340(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1341(.a(s_113), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1342(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1343(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1344(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1597(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1598(.a(gate260inter0), .b(s_150), .O(gate260inter1));
  and2  gate1599(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1600(.a(s_150), .O(gate260inter3));
  inv1  gate1601(.a(s_151), .O(gate260inter4));
  nand2 gate1602(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1603(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1604(.a(G760), .O(gate260inter7));
  inv1  gate1605(.a(G761), .O(gate260inter8));
  nand2 gate1606(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1607(.a(s_151), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1608(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1609(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1610(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1443(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1444(.a(gate267inter0), .b(s_128), .O(gate267inter1));
  and2  gate1445(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1446(.a(s_128), .O(gate267inter3));
  inv1  gate1447(.a(s_129), .O(gate267inter4));
  nand2 gate1448(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1449(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1450(.a(G648), .O(gate267inter7));
  inv1  gate1451(.a(G776), .O(gate267inter8));
  nand2 gate1452(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1453(.a(s_129), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1454(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1455(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1456(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1541(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1542(.a(gate280inter0), .b(s_142), .O(gate280inter1));
  and2  gate1543(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1544(.a(s_142), .O(gate280inter3));
  inv1  gate1545(.a(s_143), .O(gate280inter4));
  nand2 gate1546(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1547(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1548(.a(G779), .O(gate280inter7));
  inv1  gate1549(.a(G803), .O(gate280inter8));
  nand2 gate1550(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1551(.a(s_143), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1552(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1553(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1554(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1737(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1738(.a(gate288inter0), .b(s_170), .O(gate288inter1));
  and2  gate1739(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1740(.a(s_170), .O(gate288inter3));
  inv1  gate1741(.a(s_171), .O(gate288inter4));
  nand2 gate1742(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1743(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1744(.a(G791), .O(gate288inter7));
  inv1  gate1745(.a(G815), .O(gate288inter8));
  nand2 gate1746(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1747(.a(s_171), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1748(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1749(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1750(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1247(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1248(.a(gate292inter0), .b(s_100), .O(gate292inter1));
  and2  gate1249(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1250(.a(s_100), .O(gate292inter3));
  inv1  gate1251(.a(s_101), .O(gate292inter4));
  nand2 gate1252(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1253(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1254(.a(G824), .O(gate292inter7));
  inv1  gate1255(.a(G825), .O(gate292inter8));
  nand2 gate1256(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1257(.a(s_101), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1258(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1259(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1260(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate547(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate548(.a(gate293inter0), .b(s_0), .O(gate293inter1));
  and2  gate549(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate550(.a(s_0), .O(gate293inter3));
  inv1  gate551(.a(s_1), .O(gate293inter4));
  nand2 gate552(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate553(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate554(.a(G828), .O(gate293inter7));
  inv1  gate555(.a(G829), .O(gate293inter8));
  nand2 gate556(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate557(.a(s_1), .b(gate293inter3), .O(gate293inter10));
  nor2  gate558(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate559(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate560(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate841(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate842(.a(gate296inter0), .b(s_42), .O(gate296inter1));
  and2  gate843(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate844(.a(s_42), .O(gate296inter3));
  inv1  gate845(.a(s_43), .O(gate296inter4));
  nand2 gate846(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate847(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate848(.a(G826), .O(gate296inter7));
  inv1  gate849(.a(G827), .O(gate296inter8));
  nand2 gate850(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate851(.a(s_43), .b(gate296inter3), .O(gate296inter10));
  nor2  gate852(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate853(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate854(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1555(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1556(.a(gate390inter0), .b(s_144), .O(gate390inter1));
  and2  gate1557(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1558(.a(s_144), .O(gate390inter3));
  inv1  gate1559(.a(s_145), .O(gate390inter4));
  nand2 gate1560(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1561(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1562(.a(G4), .O(gate390inter7));
  inv1  gate1563(.a(G1045), .O(gate390inter8));
  nand2 gate1564(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1565(.a(s_145), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1566(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1567(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1568(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1625(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1626(.a(gate395inter0), .b(s_154), .O(gate395inter1));
  and2  gate1627(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1628(.a(s_154), .O(gate395inter3));
  inv1  gate1629(.a(s_155), .O(gate395inter4));
  nand2 gate1630(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1631(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1632(.a(G9), .O(gate395inter7));
  inv1  gate1633(.a(G1060), .O(gate395inter8));
  nand2 gate1634(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1635(.a(s_155), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1636(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1637(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1638(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate967(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate968(.a(gate397inter0), .b(s_60), .O(gate397inter1));
  and2  gate969(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate970(.a(s_60), .O(gate397inter3));
  inv1  gate971(.a(s_61), .O(gate397inter4));
  nand2 gate972(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate973(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate974(.a(G11), .O(gate397inter7));
  inv1  gate975(.a(G1066), .O(gate397inter8));
  nand2 gate976(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate977(.a(s_61), .b(gate397inter3), .O(gate397inter10));
  nor2  gate978(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate979(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate980(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1317(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1318(.a(gate402inter0), .b(s_110), .O(gate402inter1));
  and2  gate1319(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1320(.a(s_110), .O(gate402inter3));
  inv1  gate1321(.a(s_111), .O(gate402inter4));
  nand2 gate1322(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1323(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1324(.a(G16), .O(gate402inter7));
  inv1  gate1325(.a(G1081), .O(gate402inter8));
  nand2 gate1326(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1327(.a(s_111), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1328(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1329(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1330(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate673(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate674(.a(gate407inter0), .b(s_18), .O(gate407inter1));
  and2  gate675(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate676(.a(s_18), .O(gate407inter3));
  inv1  gate677(.a(s_19), .O(gate407inter4));
  nand2 gate678(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate679(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate680(.a(G21), .O(gate407inter7));
  inv1  gate681(.a(G1096), .O(gate407inter8));
  nand2 gate682(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate683(.a(s_19), .b(gate407inter3), .O(gate407inter10));
  nor2  gate684(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate685(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate686(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1233(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1234(.a(gate411inter0), .b(s_98), .O(gate411inter1));
  and2  gate1235(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1236(.a(s_98), .O(gate411inter3));
  inv1  gate1237(.a(s_99), .O(gate411inter4));
  nand2 gate1238(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1239(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1240(.a(G25), .O(gate411inter7));
  inv1  gate1241(.a(G1108), .O(gate411inter8));
  nand2 gate1242(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1243(.a(s_99), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1244(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1245(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1246(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1583(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1584(.a(gate415inter0), .b(s_148), .O(gate415inter1));
  and2  gate1585(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1586(.a(s_148), .O(gate415inter3));
  inv1  gate1587(.a(s_149), .O(gate415inter4));
  nand2 gate1588(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1589(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1590(.a(G29), .O(gate415inter7));
  inv1  gate1591(.a(G1120), .O(gate415inter8));
  nand2 gate1592(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1593(.a(s_149), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1594(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1595(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1596(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1667(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1668(.a(gate424inter0), .b(s_160), .O(gate424inter1));
  and2  gate1669(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1670(.a(s_160), .O(gate424inter3));
  inv1  gate1671(.a(s_161), .O(gate424inter4));
  nand2 gate1672(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1673(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1674(.a(G1042), .O(gate424inter7));
  inv1  gate1675(.a(G1138), .O(gate424inter8));
  nand2 gate1676(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1677(.a(s_161), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1678(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1679(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1680(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1485(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1486(.a(gate426inter0), .b(s_134), .O(gate426inter1));
  and2  gate1487(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1488(.a(s_134), .O(gate426inter3));
  inv1  gate1489(.a(s_135), .O(gate426inter4));
  nand2 gate1490(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1491(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1492(.a(G1045), .O(gate426inter7));
  inv1  gate1493(.a(G1141), .O(gate426inter8));
  nand2 gate1494(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1495(.a(s_135), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1496(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1497(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1498(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1765(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1766(.a(gate428inter0), .b(s_174), .O(gate428inter1));
  and2  gate1767(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1768(.a(s_174), .O(gate428inter3));
  inv1  gate1769(.a(s_175), .O(gate428inter4));
  nand2 gate1770(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1771(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1772(.a(G1048), .O(gate428inter7));
  inv1  gate1773(.a(G1144), .O(gate428inter8));
  nand2 gate1774(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1775(.a(s_175), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1776(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1777(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1778(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate883(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate884(.a(gate447inter0), .b(s_48), .O(gate447inter1));
  and2  gate885(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate886(.a(s_48), .O(gate447inter3));
  inv1  gate887(.a(s_49), .O(gate447inter4));
  nand2 gate888(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate889(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate890(.a(G15), .O(gate447inter7));
  inv1  gate891(.a(G1174), .O(gate447inter8));
  nand2 gate892(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate893(.a(s_49), .b(gate447inter3), .O(gate447inter10));
  nor2  gate894(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate895(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate896(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate799(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate800(.a(gate452inter0), .b(s_36), .O(gate452inter1));
  and2  gate801(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate802(.a(s_36), .O(gate452inter3));
  inv1  gate803(.a(s_37), .O(gate452inter4));
  nand2 gate804(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate805(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate806(.a(G1084), .O(gate452inter7));
  inv1  gate807(.a(G1180), .O(gate452inter8));
  nand2 gate808(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate809(.a(s_37), .b(gate452inter3), .O(gate452inter10));
  nor2  gate810(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate811(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate812(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1499(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1500(.a(gate455inter0), .b(s_136), .O(gate455inter1));
  and2  gate1501(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1502(.a(s_136), .O(gate455inter3));
  inv1  gate1503(.a(s_137), .O(gate455inter4));
  nand2 gate1504(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1505(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1506(.a(G19), .O(gate455inter7));
  inv1  gate1507(.a(G1186), .O(gate455inter8));
  nand2 gate1508(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1509(.a(s_137), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1510(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1511(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1512(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate589(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate590(.a(gate461inter0), .b(s_6), .O(gate461inter1));
  and2  gate591(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate592(.a(s_6), .O(gate461inter3));
  inv1  gate593(.a(s_7), .O(gate461inter4));
  nand2 gate594(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate595(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate596(.a(G22), .O(gate461inter7));
  inv1  gate597(.a(G1195), .O(gate461inter8));
  nand2 gate598(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate599(.a(s_7), .b(gate461inter3), .O(gate461inter10));
  nor2  gate600(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate601(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate602(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate729(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate730(.a(gate470inter0), .b(s_26), .O(gate470inter1));
  and2  gate731(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate732(.a(s_26), .O(gate470inter3));
  inv1  gate733(.a(s_27), .O(gate470inter4));
  nand2 gate734(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate735(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate736(.a(G1111), .O(gate470inter7));
  inv1  gate737(.a(G1207), .O(gate470inter8));
  nand2 gate738(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate739(.a(s_27), .b(gate470inter3), .O(gate470inter10));
  nor2  gate740(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate741(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate742(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1079(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1080(.a(gate471inter0), .b(s_76), .O(gate471inter1));
  and2  gate1081(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1082(.a(s_76), .O(gate471inter3));
  inv1  gate1083(.a(s_77), .O(gate471inter4));
  nand2 gate1084(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1085(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1086(.a(G27), .O(gate471inter7));
  inv1  gate1087(.a(G1210), .O(gate471inter8));
  nand2 gate1088(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1089(.a(s_77), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1090(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1091(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1092(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1709(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1710(.a(gate475inter0), .b(s_166), .O(gate475inter1));
  and2  gate1711(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1712(.a(s_166), .O(gate475inter3));
  inv1  gate1713(.a(s_167), .O(gate475inter4));
  nand2 gate1714(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1715(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1716(.a(G29), .O(gate475inter7));
  inv1  gate1717(.a(G1216), .O(gate475inter8));
  nand2 gate1718(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1719(.a(s_167), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1720(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1721(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1722(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1751(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1752(.a(gate477inter0), .b(s_172), .O(gate477inter1));
  and2  gate1753(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1754(.a(s_172), .O(gate477inter3));
  inv1  gate1755(.a(s_173), .O(gate477inter4));
  nand2 gate1756(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1757(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1758(.a(G30), .O(gate477inter7));
  inv1  gate1759(.a(G1219), .O(gate477inter8));
  nand2 gate1760(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1761(.a(s_173), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1762(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1763(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1764(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate771(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate772(.a(gate478inter0), .b(s_32), .O(gate478inter1));
  and2  gate773(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate774(.a(s_32), .O(gate478inter3));
  inv1  gate775(.a(s_33), .O(gate478inter4));
  nand2 gate776(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate777(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate778(.a(G1123), .O(gate478inter7));
  inv1  gate779(.a(G1219), .O(gate478inter8));
  nand2 gate780(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate781(.a(s_33), .b(gate478inter3), .O(gate478inter10));
  nor2  gate782(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate783(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate784(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1261(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1262(.a(gate479inter0), .b(s_102), .O(gate479inter1));
  and2  gate1263(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1264(.a(s_102), .O(gate479inter3));
  inv1  gate1265(.a(s_103), .O(gate479inter4));
  nand2 gate1266(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1267(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1268(.a(G31), .O(gate479inter7));
  inv1  gate1269(.a(G1222), .O(gate479inter8));
  nand2 gate1270(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1271(.a(s_103), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1272(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1273(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1274(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1373(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1374(.a(gate485inter0), .b(s_118), .O(gate485inter1));
  and2  gate1375(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1376(.a(s_118), .O(gate485inter3));
  inv1  gate1377(.a(s_119), .O(gate485inter4));
  nand2 gate1378(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1379(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1380(.a(G1232), .O(gate485inter7));
  inv1  gate1381(.a(G1233), .O(gate485inter8));
  nand2 gate1382(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1383(.a(s_119), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1384(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1385(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1386(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate757(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate758(.a(gate489inter0), .b(s_30), .O(gate489inter1));
  and2  gate759(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate760(.a(s_30), .O(gate489inter3));
  inv1  gate761(.a(s_31), .O(gate489inter4));
  nand2 gate762(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate763(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate764(.a(G1240), .O(gate489inter7));
  inv1  gate765(.a(G1241), .O(gate489inter8));
  nand2 gate766(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate767(.a(s_31), .b(gate489inter3), .O(gate489inter10));
  nor2  gate768(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate769(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate770(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1569(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1570(.a(gate492inter0), .b(s_146), .O(gate492inter1));
  and2  gate1571(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1572(.a(s_146), .O(gate492inter3));
  inv1  gate1573(.a(s_147), .O(gate492inter4));
  nand2 gate1574(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1575(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1576(.a(G1246), .O(gate492inter7));
  inv1  gate1577(.a(G1247), .O(gate492inter8));
  nand2 gate1578(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1579(.a(s_147), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1580(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1581(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1582(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate827(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate828(.a(gate500inter0), .b(s_40), .O(gate500inter1));
  and2  gate829(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate830(.a(s_40), .O(gate500inter3));
  inv1  gate831(.a(s_41), .O(gate500inter4));
  nand2 gate832(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate833(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate834(.a(G1262), .O(gate500inter7));
  inv1  gate835(.a(G1263), .O(gate500inter8));
  nand2 gate836(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate837(.a(s_41), .b(gate500inter3), .O(gate500inter10));
  nor2  gate838(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate839(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate840(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate603(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate604(.a(gate508inter0), .b(s_8), .O(gate508inter1));
  and2  gate605(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate606(.a(s_8), .O(gate508inter3));
  inv1  gate607(.a(s_9), .O(gate508inter4));
  nand2 gate608(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate609(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate610(.a(G1278), .O(gate508inter7));
  inv1  gate611(.a(G1279), .O(gate508inter8));
  nand2 gate612(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate613(.a(s_9), .b(gate508inter3), .O(gate508inter10));
  nor2  gate614(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate615(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate616(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate869(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate870(.a(gate510inter0), .b(s_46), .O(gate510inter1));
  and2  gate871(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate872(.a(s_46), .O(gate510inter3));
  inv1  gate873(.a(s_47), .O(gate510inter4));
  nand2 gate874(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate875(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate876(.a(G1282), .O(gate510inter7));
  inv1  gate877(.a(G1283), .O(gate510inter8));
  nand2 gate878(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate879(.a(s_47), .b(gate510inter3), .O(gate510inter10));
  nor2  gate880(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate881(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate882(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate743(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate744(.a(gate511inter0), .b(s_28), .O(gate511inter1));
  and2  gate745(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate746(.a(s_28), .O(gate511inter3));
  inv1  gate747(.a(s_29), .O(gate511inter4));
  nand2 gate748(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate749(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate750(.a(G1284), .O(gate511inter7));
  inv1  gate751(.a(G1285), .O(gate511inter8));
  nand2 gate752(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate753(.a(s_29), .b(gate511inter3), .O(gate511inter10));
  nor2  gate754(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate755(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate756(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule