module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate673(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate674(.a(gate11inter0), .b(s_18), .O(gate11inter1));
  and2  gate675(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate676(.a(s_18), .O(gate11inter3));
  inv1  gate677(.a(s_19), .O(gate11inter4));
  nand2 gate678(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate679(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate680(.a(G5), .O(gate11inter7));
  inv1  gate681(.a(G6), .O(gate11inter8));
  nand2 gate682(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate683(.a(s_19), .b(gate11inter3), .O(gate11inter10));
  nor2  gate684(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate685(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate686(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1401(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1402(.a(gate15inter0), .b(s_122), .O(gate15inter1));
  and2  gate1403(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1404(.a(s_122), .O(gate15inter3));
  inv1  gate1405(.a(s_123), .O(gate15inter4));
  nand2 gate1406(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1407(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1408(.a(G13), .O(gate15inter7));
  inv1  gate1409(.a(G14), .O(gate15inter8));
  nand2 gate1410(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1411(.a(s_123), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1412(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1413(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1414(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate575(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate576(.a(gate16inter0), .b(s_4), .O(gate16inter1));
  and2  gate577(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate578(.a(s_4), .O(gate16inter3));
  inv1  gate579(.a(s_5), .O(gate16inter4));
  nand2 gate580(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate581(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate582(.a(G15), .O(gate16inter7));
  inv1  gate583(.a(G16), .O(gate16inter8));
  nand2 gate584(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate585(.a(s_5), .b(gate16inter3), .O(gate16inter10));
  nor2  gate586(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate587(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate588(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2563(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2564(.a(gate19inter0), .b(s_288), .O(gate19inter1));
  and2  gate2565(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2566(.a(s_288), .O(gate19inter3));
  inv1  gate2567(.a(s_289), .O(gate19inter4));
  nand2 gate2568(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2569(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2570(.a(G21), .O(gate19inter7));
  inv1  gate2571(.a(G22), .O(gate19inter8));
  nand2 gate2572(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2573(.a(s_289), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2574(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2575(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2576(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1429(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1430(.a(gate23inter0), .b(s_126), .O(gate23inter1));
  and2  gate1431(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1432(.a(s_126), .O(gate23inter3));
  inv1  gate1433(.a(s_127), .O(gate23inter4));
  nand2 gate1434(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1435(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1436(.a(G29), .O(gate23inter7));
  inv1  gate1437(.a(G30), .O(gate23inter8));
  nand2 gate1438(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1439(.a(s_127), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1440(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1441(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1442(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1597(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1598(.a(gate25inter0), .b(s_150), .O(gate25inter1));
  and2  gate1599(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1600(.a(s_150), .O(gate25inter3));
  inv1  gate1601(.a(s_151), .O(gate25inter4));
  nand2 gate1602(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1603(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1604(.a(G1), .O(gate25inter7));
  inv1  gate1605(.a(G5), .O(gate25inter8));
  nand2 gate1606(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1607(.a(s_151), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1608(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1609(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1610(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate701(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate702(.a(gate27inter0), .b(s_22), .O(gate27inter1));
  and2  gate703(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate704(.a(s_22), .O(gate27inter3));
  inv1  gate705(.a(s_23), .O(gate27inter4));
  nand2 gate706(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate707(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate708(.a(G2), .O(gate27inter7));
  inv1  gate709(.a(G6), .O(gate27inter8));
  nand2 gate710(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate711(.a(s_23), .b(gate27inter3), .O(gate27inter10));
  nor2  gate712(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate713(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate714(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1443(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1444(.a(gate29inter0), .b(s_128), .O(gate29inter1));
  and2  gate1445(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1446(.a(s_128), .O(gate29inter3));
  inv1  gate1447(.a(s_129), .O(gate29inter4));
  nand2 gate1448(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1449(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1450(.a(G3), .O(gate29inter7));
  inv1  gate1451(.a(G7), .O(gate29inter8));
  nand2 gate1452(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1453(.a(s_129), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1454(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1455(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1456(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate841(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate842(.a(gate31inter0), .b(s_42), .O(gate31inter1));
  and2  gate843(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate844(.a(s_42), .O(gate31inter3));
  inv1  gate845(.a(s_43), .O(gate31inter4));
  nand2 gate846(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate847(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate848(.a(G4), .O(gate31inter7));
  inv1  gate849(.a(G8), .O(gate31inter8));
  nand2 gate850(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate851(.a(s_43), .b(gate31inter3), .O(gate31inter10));
  nor2  gate852(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate853(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate854(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate799(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate800(.a(gate41inter0), .b(s_36), .O(gate41inter1));
  and2  gate801(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate802(.a(s_36), .O(gate41inter3));
  inv1  gate803(.a(s_37), .O(gate41inter4));
  nand2 gate804(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate805(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate806(.a(G1), .O(gate41inter7));
  inv1  gate807(.a(G266), .O(gate41inter8));
  nand2 gate808(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate809(.a(s_37), .b(gate41inter3), .O(gate41inter10));
  nor2  gate810(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate811(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate812(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1653(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1654(.a(gate45inter0), .b(s_158), .O(gate45inter1));
  and2  gate1655(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1656(.a(s_158), .O(gate45inter3));
  inv1  gate1657(.a(s_159), .O(gate45inter4));
  nand2 gate1658(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1659(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1660(.a(G5), .O(gate45inter7));
  inv1  gate1661(.a(G272), .O(gate45inter8));
  nand2 gate1662(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1663(.a(s_159), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1664(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1665(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1666(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2549(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2550(.a(gate47inter0), .b(s_286), .O(gate47inter1));
  and2  gate2551(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2552(.a(s_286), .O(gate47inter3));
  inv1  gate2553(.a(s_287), .O(gate47inter4));
  nand2 gate2554(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2555(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2556(.a(G7), .O(gate47inter7));
  inv1  gate2557(.a(G275), .O(gate47inter8));
  nand2 gate2558(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2559(.a(s_287), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2560(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2561(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2562(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1933(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1934(.a(gate49inter0), .b(s_198), .O(gate49inter1));
  and2  gate1935(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1936(.a(s_198), .O(gate49inter3));
  inv1  gate1937(.a(s_199), .O(gate49inter4));
  nand2 gate1938(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1939(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1940(.a(G9), .O(gate49inter7));
  inv1  gate1941(.a(G278), .O(gate49inter8));
  nand2 gate1942(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1943(.a(s_199), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1944(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1945(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1946(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1303(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1304(.a(gate53inter0), .b(s_108), .O(gate53inter1));
  and2  gate1305(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1306(.a(s_108), .O(gate53inter3));
  inv1  gate1307(.a(s_109), .O(gate53inter4));
  nand2 gate1308(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1309(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1310(.a(G13), .O(gate53inter7));
  inv1  gate1311(.a(G284), .O(gate53inter8));
  nand2 gate1312(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1313(.a(s_109), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1314(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1315(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1316(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate827(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate828(.a(gate54inter0), .b(s_40), .O(gate54inter1));
  and2  gate829(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate830(.a(s_40), .O(gate54inter3));
  inv1  gate831(.a(s_41), .O(gate54inter4));
  nand2 gate832(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate833(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate834(.a(G14), .O(gate54inter7));
  inv1  gate835(.a(G284), .O(gate54inter8));
  nand2 gate836(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate837(.a(s_41), .b(gate54inter3), .O(gate54inter10));
  nor2  gate838(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate839(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate840(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1751(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1752(.a(gate57inter0), .b(s_172), .O(gate57inter1));
  and2  gate1753(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1754(.a(s_172), .O(gate57inter3));
  inv1  gate1755(.a(s_173), .O(gate57inter4));
  nand2 gate1756(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1757(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1758(.a(G17), .O(gate57inter7));
  inv1  gate1759(.a(G290), .O(gate57inter8));
  nand2 gate1760(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1761(.a(s_173), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1762(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1763(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1764(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1247(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1248(.a(gate59inter0), .b(s_100), .O(gate59inter1));
  and2  gate1249(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1250(.a(s_100), .O(gate59inter3));
  inv1  gate1251(.a(s_101), .O(gate59inter4));
  nand2 gate1252(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1253(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1254(.a(G19), .O(gate59inter7));
  inv1  gate1255(.a(G293), .O(gate59inter8));
  nand2 gate1256(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1257(.a(s_101), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1258(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1259(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1260(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1709(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1710(.a(gate60inter0), .b(s_166), .O(gate60inter1));
  and2  gate1711(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1712(.a(s_166), .O(gate60inter3));
  inv1  gate1713(.a(s_167), .O(gate60inter4));
  nand2 gate1714(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1715(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1716(.a(G20), .O(gate60inter7));
  inv1  gate1717(.a(G293), .O(gate60inter8));
  nand2 gate1718(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1719(.a(s_167), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1720(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1721(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1722(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2521(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2522(.a(gate61inter0), .b(s_282), .O(gate61inter1));
  and2  gate2523(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2524(.a(s_282), .O(gate61inter3));
  inv1  gate2525(.a(s_283), .O(gate61inter4));
  nand2 gate2526(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2527(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2528(.a(G21), .O(gate61inter7));
  inv1  gate2529(.a(G296), .O(gate61inter8));
  nand2 gate2530(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2531(.a(s_283), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2532(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2533(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2534(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate645(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate646(.a(gate64inter0), .b(s_14), .O(gate64inter1));
  and2  gate647(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate648(.a(s_14), .O(gate64inter3));
  inv1  gate649(.a(s_15), .O(gate64inter4));
  nand2 gate650(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate651(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate652(.a(G24), .O(gate64inter7));
  inv1  gate653(.a(G299), .O(gate64inter8));
  nand2 gate654(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate655(.a(s_15), .b(gate64inter3), .O(gate64inter10));
  nor2  gate656(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate657(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate658(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate547(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate548(.a(gate65inter0), .b(s_0), .O(gate65inter1));
  and2  gate549(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate550(.a(s_0), .O(gate65inter3));
  inv1  gate551(.a(s_1), .O(gate65inter4));
  nand2 gate552(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate553(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate554(.a(G25), .O(gate65inter7));
  inv1  gate555(.a(G302), .O(gate65inter8));
  nand2 gate556(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate557(.a(s_1), .b(gate65inter3), .O(gate65inter10));
  nor2  gate558(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate559(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate560(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1779(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1780(.a(gate69inter0), .b(s_176), .O(gate69inter1));
  and2  gate1781(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1782(.a(s_176), .O(gate69inter3));
  inv1  gate1783(.a(s_177), .O(gate69inter4));
  nand2 gate1784(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1785(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1786(.a(G29), .O(gate69inter7));
  inv1  gate1787(.a(G308), .O(gate69inter8));
  nand2 gate1788(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1789(.a(s_177), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1790(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1791(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1792(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2507(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2508(.a(gate70inter0), .b(s_280), .O(gate70inter1));
  and2  gate2509(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2510(.a(s_280), .O(gate70inter3));
  inv1  gate2511(.a(s_281), .O(gate70inter4));
  nand2 gate2512(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2513(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2514(.a(G30), .O(gate70inter7));
  inv1  gate2515(.a(G308), .O(gate70inter8));
  nand2 gate2516(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2517(.a(s_281), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2518(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2519(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2520(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1499(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1500(.a(gate71inter0), .b(s_136), .O(gate71inter1));
  and2  gate1501(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1502(.a(s_136), .O(gate71inter3));
  inv1  gate1503(.a(s_137), .O(gate71inter4));
  nand2 gate1504(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1505(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1506(.a(G31), .O(gate71inter7));
  inv1  gate1507(.a(G311), .O(gate71inter8));
  nand2 gate1508(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1509(.a(s_137), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1510(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1511(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1512(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1905(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1906(.a(gate73inter0), .b(s_194), .O(gate73inter1));
  and2  gate1907(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1908(.a(s_194), .O(gate73inter3));
  inv1  gate1909(.a(s_195), .O(gate73inter4));
  nand2 gate1910(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1911(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1912(.a(G1), .O(gate73inter7));
  inv1  gate1913(.a(G314), .O(gate73inter8));
  nand2 gate1914(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1915(.a(s_195), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1916(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1917(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1918(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1527(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1528(.a(gate75inter0), .b(s_140), .O(gate75inter1));
  and2  gate1529(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1530(.a(s_140), .O(gate75inter3));
  inv1  gate1531(.a(s_141), .O(gate75inter4));
  nand2 gate1532(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1533(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1534(.a(G9), .O(gate75inter7));
  inv1  gate1535(.a(G317), .O(gate75inter8));
  nand2 gate1536(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1537(.a(s_141), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1538(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1539(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1540(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1205(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1206(.a(gate76inter0), .b(s_94), .O(gate76inter1));
  and2  gate1207(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1208(.a(s_94), .O(gate76inter3));
  inv1  gate1209(.a(s_95), .O(gate76inter4));
  nand2 gate1210(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1211(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1212(.a(G13), .O(gate76inter7));
  inv1  gate1213(.a(G317), .O(gate76inter8));
  nand2 gate1214(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1215(.a(s_95), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1216(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1217(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1218(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2367(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2368(.a(gate78inter0), .b(s_260), .O(gate78inter1));
  and2  gate2369(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2370(.a(s_260), .O(gate78inter3));
  inv1  gate2371(.a(s_261), .O(gate78inter4));
  nand2 gate2372(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2373(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2374(.a(G6), .O(gate78inter7));
  inv1  gate2375(.a(G320), .O(gate78inter8));
  nand2 gate2376(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2377(.a(s_261), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2378(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2379(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2380(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1149(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1150(.a(gate82inter0), .b(s_86), .O(gate82inter1));
  and2  gate1151(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1152(.a(s_86), .O(gate82inter3));
  inv1  gate1153(.a(s_87), .O(gate82inter4));
  nand2 gate1154(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1155(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1156(.a(G7), .O(gate82inter7));
  inv1  gate1157(.a(G326), .O(gate82inter8));
  nand2 gate1158(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1159(.a(s_87), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1160(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1161(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1162(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate589(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate590(.a(gate84inter0), .b(s_6), .O(gate84inter1));
  and2  gate591(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate592(.a(s_6), .O(gate84inter3));
  inv1  gate593(.a(s_7), .O(gate84inter4));
  nand2 gate594(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate595(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate596(.a(G15), .O(gate84inter7));
  inv1  gate597(.a(G329), .O(gate84inter8));
  nand2 gate598(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate599(.a(s_7), .b(gate84inter3), .O(gate84inter10));
  nor2  gate600(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate601(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate602(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2633(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2634(.a(gate89inter0), .b(s_298), .O(gate89inter1));
  and2  gate2635(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2636(.a(s_298), .O(gate89inter3));
  inv1  gate2637(.a(s_299), .O(gate89inter4));
  nand2 gate2638(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2639(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2640(.a(G17), .O(gate89inter7));
  inv1  gate2641(.a(G338), .O(gate89inter8));
  nand2 gate2642(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2643(.a(s_299), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2644(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2645(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2646(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1177(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1178(.a(gate91inter0), .b(s_90), .O(gate91inter1));
  and2  gate1179(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1180(.a(s_90), .O(gate91inter3));
  inv1  gate1181(.a(s_91), .O(gate91inter4));
  nand2 gate1182(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1183(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1184(.a(G25), .O(gate91inter7));
  inv1  gate1185(.a(G341), .O(gate91inter8));
  nand2 gate1186(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1187(.a(s_91), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1188(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1189(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1190(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate561(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate562(.a(gate93inter0), .b(s_2), .O(gate93inter1));
  and2  gate563(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate564(.a(s_2), .O(gate93inter3));
  inv1  gate565(.a(s_3), .O(gate93inter4));
  nand2 gate566(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate567(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate568(.a(G18), .O(gate93inter7));
  inv1  gate569(.a(G344), .O(gate93inter8));
  nand2 gate570(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate571(.a(s_3), .b(gate93inter3), .O(gate93inter10));
  nor2  gate572(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate573(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate574(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2717(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2718(.a(gate98inter0), .b(s_310), .O(gate98inter1));
  and2  gate2719(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2720(.a(s_310), .O(gate98inter3));
  inv1  gate2721(.a(s_311), .O(gate98inter4));
  nand2 gate2722(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2723(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2724(.a(G23), .O(gate98inter7));
  inv1  gate2725(.a(G350), .O(gate98inter8));
  nand2 gate2726(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2727(.a(s_311), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2728(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2729(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2730(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2437(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2438(.a(gate100inter0), .b(s_270), .O(gate100inter1));
  and2  gate2439(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2440(.a(s_270), .O(gate100inter3));
  inv1  gate2441(.a(s_271), .O(gate100inter4));
  nand2 gate2442(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2443(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2444(.a(G31), .O(gate100inter7));
  inv1  gate2445(.a(G353), .O(gate100inter8));
  nand2 gate2446(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2447(.a(s_271), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2448(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2449(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2450(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1121(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1122(.a(gate103inter0), .b(s_82), .O(gate103inter1));
  and2  gate1123(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1124(.a(s_82), .O(gate103inter3));
  inv1  gate1125(.a(s_83), .O(gate103inter4));
  nand2 gate1126(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1127(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1128(.a(G28), .O(gate103inter7));
  inv1  gate1129(.a(G359), .O(gate103inter8));
  nand2 gate1130(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1131(.a(s_83), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1132(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1133(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1134(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1877(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1878(.a(gate104inter0), .b(s_190), .O(gate104inter1));
  and2  gate1879(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1880(.a(s_190), .O(gate104inter3));
  inv1  gate1881(.a(s_191), .O(gate104inter4));
  nand2 gate1882(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1883(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1884(.a(G32), .O(gate104inter7));
  inv1  gate1885(.a(G359), .O(gate104inter8));
  nand2 gate1886(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1887(.a(s_191), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1888(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1889(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1890(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2297(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2298(.a(gate106inter0), .b(s_250), .O(gate106inter1));
  and2  gate2299(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2300(.a(s_250), .O(gate106inter3));
  inv1  gate2301(.a(s_251), .O(gate106inter4));
  nand2 gate2302(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2303(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2304(.a(G364), .O(gate106inter7));
  inv1  gate2305(.a(G365), .O(gate106inter8));
  nand2 gate2306(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2307(.a(s_251), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2308(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2309(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2310(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2269(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2270(.a(gate111inter0), .b(s_246), .O(gate111inter1));
  and2  gate2271(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2272(.a(s_246), .O(gate111inter3));
  inv1  gate2273(.a(s_247), .O(gate111inter4));
  nand2 gate2274(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2275(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2276(.a(G374), .O(gate111inter7));
  inv1  gate2277(.a(G375), .O(gate111inter8));
  nand2 gate2278(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2279(.a(s_247), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2280(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2281(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2282(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1583(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1584(.a(gate114inter0), .b(s_148), .O(gate114inter1));
  and2  gate1585(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1586(.a(s_148), .O(gate114inter3));
  inv1  gate1587(.a(s_149), .O(gate114inter4));
  nand2 gate1588(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1589(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1590(.a(G380), .O(gate114inter7));
  inv1  gate1591(.a(G381), .O(gate114inter8));
  nand2 gate1592(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1593(.a(s_149), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1594(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1595(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1596(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate869(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate870(.a(gate115inter0), .b(s_46), .O(gate115inter1));
  and2  gate871(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate872(.a(s_46), .O(gate115inter3));
  inv1  gate873(.a(s_47), .O(gate115inter4));
  nand2 gate874(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate875(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate876(.a(G382), .O(gate115inter7));
  inv1  gate877(.a(G383), .O(gate115inter8));
  nand2 gate878(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate879(.a(s_47), .b(gate115inter3), .O(gate115inter10));
  nor2  gate880(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate881(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate882(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1695(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1696(.a(gate117inter0), .b(s_164), .O(gate117inter1));
  and2  gate1697(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1698(.a(s_164), .O(gate117inter3));
  inv1  gate1699(.a(s_165), .O(gate117inter4));
  nand2 gate1700(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1701(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1702(.a(G386), .O(gate117inter7));
  inv1  gate1703(.a(G387), .O(gate117inter8));
  nand2 gate1704(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1705(.a(s_165), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1706(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1707(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1708(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2017(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2018(.a(gate119inter0), .b(s_210), .O(gate119inter1));
  and2  gate2019(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2020(.a(s_210), .O(gate119inter3));
  inv1  gate2021(.a(s_211), .O(gate119inter4));
  nand2 gate2022(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2023(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2024(.a(G390), .O(gate119inter7));
  inv1  gate2025(.a(G391), .O(gate119inter8));
  nand2 gate2026(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2027(.a(s_211), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2028(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2029(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2030(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1051(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1052(.a(gate120inter0), .b(s_72), .O(gate120inter1));
  and2  gate1053(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1054(.a(s_72), .O(gate120inter3));
  inv1  gate1055(.a(s_73), .O(gate120inter4));
  nand2 gate1056(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1057(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1058(.a(G392), .O(gate120inter7));
  inv1  gate1059(.a(G393), .O(gate120inter8));
  nand2 gate1060(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1061(.a(s_73), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1062(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1063(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1064(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1359(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1360(.a(gate122inter0), .b(s_116), .O(gate122inter1));
  and2  gate1361(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1362(.a(s_116), .O(gate122inter3));
  inv1  gate1363(.a(s_117), .O(gate122inter4));
  nand2 gate1364(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1365(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1366(.a(G396), .O(gate122inter7));
  inv1  gate1367(.a(G397), .O(gate122inter8));
  nand2 gate1368(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1369(.a(s_117), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1370(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1371(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1372(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2101(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2102(.a(gate136inter0), .b(s_222), .O(gate136inter1));
  and2  gate2103(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2104(.a(s_222), .O(gate136inter3));
  inv1  gate2105(.a(s_223), .O(gate136inter4));
  nand2 gate2106(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2107(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2108(.a(G424), .O(gate136inter7));
  inv1  gate2109(.a(G425), .O(gate136inter8));
  nand2 gate2110(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2111(.a(s_223), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2112(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2113(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2114(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1723(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1724(.a(gate137inter0), .b(s_168), .O(gate137inter1));
  and2  gate1725(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1726(.a(s_168), .O(gate137inter3));
  inv1  gate1727(.a(s_169), .O(gate137inter4));
  nand2 gate1728(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1729(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1730(.a(G426), .O(gate137inter7));
  inv1  gate1731(.a(G429), .O(gate137inter8));
  nand2 gate1732(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1733(.a(s_169), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1734(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1735(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1736(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1807(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1808(.a(gate139inter0), .b(s_180), .O(gate139inter1));
  and2  gate1809(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1810(.a(s_180), .O(gate139inter3));
  inv1  gate1811(.a(s_181), .O(gate139inter4));
  nand2 gate1812(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1813(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1814(.a(G438), .O(gate139inter7));
  inv1  gate1815(.a(G441), .O(gate139inter8));
  nand2 gate1816(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1817(.a(s_181), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1818(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1819(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1820(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2059(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2060(.a(gate140inter0), .b(s_216), .O(gate140inter1));
  and2  gate2061(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2062(.a(s_216), .O(gate140inter3));
  inv1  gate2063(.a(s_217), .O(gate140inter4));
  nand2 gate2064(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2065(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2066(.a(G444), .O(gate140inter7));
  inv1  gate2067(.a(G447), .O(gate140inter8));
  nand2 gate2068(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2069(.a(s_217), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2070(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2071(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2072(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2003(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2004(.a(gate142inter0), .b(s_208), .O(gate142inter1));
  and2  gate2005(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2006(.a(s_208), .O(gate142inter3));
  inv1  gate2007(.a(s_209), .O(gate142inter4));
  nand2 gate2008(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2009(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2010(.a(G456), .O(gate142inter7));
  inv1  gate2011(.a(G459), .O(gate142inter8));
  nand2 gate2012(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2013(.a(s_209), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2014(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2015(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2016(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2451(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2452(.a(gate146inter0), .b(s_272), .O(gate146inter1));
  and2  gate2453(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2454(.a(s_272), .O(gate146inter3));
  inv1  gate2455(.a(s_273), .O(gate146inter4));
  nand2 gate2456(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2457(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2458(.a(G480), .O(gate146inter7));
  inv1  gate2459(.a(G483), .O(gate146inter8));
  nand2 gate2460(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2461(.a(s_273), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2462(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2463(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2464(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate743(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate744(.a(gate148inter0), .b(s_28), .O(gate148inter1));
  and2  gate745(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate746(.a(s_28), .O(gate148inter3));
  inv1  gate747(.a(s_29), .O(gate148inter4));
  nand2 gate748(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate749(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate750(.a(G492), .O(gate148inter7));
  inv1  gate751(.a(G495), .O(gate148inter8));
  nand2 gate752(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate753(.a(s_29), .b(gate148inter3), .O(gate148inter10));
  nor2  gate754(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate755(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate756(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2255(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2256(.a(gate151inter0), .b(s_244), .O(gate151inter1));
  and2  gate2257(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2258(.a(s_244), .O(gate151inter3));
  inv1  gate2259(.a(s_245), .O(gate151inter4));
  nand2 gate2260(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2261(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2262(.a(G510), .O(gate151inter7));
  inv1  gate2263(.a(G513), .O(gate151inter8));
  nand2 gate2264(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2265(.a(s_245), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2266(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2267(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2268(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate687(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate688(.a(gate153inter0), .b(s_20), .O(gate153inter1));
  and2  gate689(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate690(.a(s_20), .O(gate153inter3));
  inv1  gate691(.a(s_21), .O(gate153inter4));
  nand2 gate692(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate693(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate694(.a(G426), .O(gate153inter7));
  inv1  gate695(.a(G522), .O(gate153inter8));
  nand2 gate696(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate697(.a(s_21), .b(gate153inter3), .O(gate153inter10));
  nor2  gate698(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate699(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate700(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2703(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2704(.a(gate156inter0), .b(s_308), .O(gate156inter1));
  and2  gate2705(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2706(.a(s_308), .O(gate156inter3));
  inv1  gate2707(.a(s_309), .O(gate156inter4));
  nand2 gate2708(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2709(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2710(.a(G435), .O(gate156inter7));
  inv1  gate2711(.a(G525), .O(gate156inter8));
  nand2 gate2712(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2713(.a(s_309), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2714(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2715(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2716(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1023(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1024(.a(gate158inter0), .b(s_68), .O(gate158inter1));
  and2  gate1025(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1026(.a(s_68), .O(gate158inter3));
  inv1  gate1027(.a(s_69), .O(gate158inter4));
  nand2 gate1028(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1029(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1030(.a(G441), .O(gate158inter7));
  inv1  gate1031(.a(G528), .O(gate158inter8));
  nand2 gate1032(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1033(.a(s_69), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1034(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1035(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1036(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1191(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1192(.a(gate159inter0), .b(s_92), .O(gate159inter1));
  and2  gate1193(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1194(.a(s_92), .O(gate159inter3));
  inv1  gate1195(.a(s_93), .O(gate159inter4));
  nand2 gate1196(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1197(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1198(.a(G444), .O(gate159inter7));
  inv1  gate1199(.a(G531), .O(gate159inter8));
  nand2 gate1200(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1201(.a(s_93), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1202(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1203(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1204(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1863(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1864(.a(gate160inter0), .b(s_188), .O(gate160inter1));
  and2  gate1865(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1866(.a(s_188), .O(gate160inter3));
  inv1  gate1867(.a(s_189), .O(gate160inter4));
  nand2 gate1868(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1869(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1870(.a(G447), .O(gate160inter7));
  inv1  gate1871(.a(G531), .O(gate160inter8));
  nand2 gate1872(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1873(.a(s_189), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1874(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1875(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1876(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate2577(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2578(.a(gate163inter0), .b(s_290), .O(gate163inter1));
  and2  gate2579(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2580(.a(s_290), .O(gate163inter3));
  inv1  gate2581(.a(s_291), .O(gate163inter4));
  nand2 gate2582(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2583(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2584(.a(G456), .O(gate163inter7));
  inv1  gate2585(.a(G537), .O(gate163inter8));
  nand2 gate2586(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2587(.a(s_291), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2588(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2589(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2590(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2395(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2396(.a(gate165inter0), .b(s_264), .O(gate165inter1));
  and2  gate2397(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2398(.a(s_264), .O(gate165inter3));
  inv1  gate2399(.a(s_265), .O(gate165inter4));
  nand2 gate2400(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2401(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2402(.a(G462), .O(gate165inter7));
  inv1  gate2403(.a(G540), .O(gate165inter8));
  nand2 gate2404(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2405(.a(s_265), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2406(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2407(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2408(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate939(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate940(.a(gate172inter0), .b(s_56), .O(gate172inter1));
  and2  gate941(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate942(.a(s_56), .O(gate172inter3));
  inv1  gate943(.a(s_57), .O(gate172inter4));
  nand2 gate944(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate945(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate946(.a(G483), .O(gate172inter7));
  inv1  gate947(.a(G549), .O(gate172inter8));
  nand2 gate948(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate949(.a(s_57), .b(gate172inter3), .O(gate172inter10));
  nor2  gate950(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate951(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate952(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1793(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1794(.a(gate173inter0), .b(s_178), .O(gate173inter1));
  and2  gate1795(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1796(.a(s_178), .O(gate173inter3));
  inv1  gate1797(.a(s_179), .O(gate173inter4));
  nand2 gate1798(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1799(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1800(.a(G486), .O(gate173inter7));
  inv1  gate1801(.a(G552), .O(gate173inter8));
  nand2 gate1802(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1803(.a(s_179), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1804(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1805(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1806(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate883(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate884(.a(gate177inter0), .b(s_48), .O(gate177inter1));
  and2  gate885(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate886(.a(s_48), .O(gate177inter3));
  inv1  gate887(.a(s_49), .O(gate177inter4));
  nand2 gate888(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate889(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate890(.a(G498), .O(gate177inter7));
  inv1  gate891(.a(G558), .O(gate177inter8));
  nand2 gate892(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate893(.a(s_49), .b(gate177inter3), .O(gate177inter10));
  nor2  gate894(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate895(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate896(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate2689(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2690(.a(gate178inter0), .b(s_306), .O(gate178inter1));
  and2  gate2691(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2692(.a(s_306), .O(gate178inter3));
  inv1  gate2693(.a(s_307), .O(gate178inter4));
  nand2 gate2694(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2695(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2696(.a(G501), .O(gate178inter7));
  inv1  gate2697(.a(G558), .O(gate178inter8));
  nand2 gate2698(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2699(.a(s_307), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2700(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2701(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2702(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1541(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1542(.a(gate186inter0), .b(s_142), .O(gate186inter1));
  and2  gate1543(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1544(.a(s_142), .O(gate186inter3));
  inv1  gate1545(.a(s_143), .O(gate186inter4));
  nand2 gate1546(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1547(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1548(.a(G572), .O(gate186inter7));
  inv1  gate1549(.a(G573), .O(gate186inter8));
  nand2 gate1550(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1551(.a(s_143), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1552(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1553(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1554(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate603(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate604(.a(gate188inter0), .b(s_8), .O(gate188inter1));
  and2  gate605(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate606(.a(s_8), .O(gate188inter3));
  inv1  gate607(.a(s_9), .O(gate188inter4));
  nand2 gate608(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate609(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate610(.a(G576), .O(gate188inter7));
  inv1  gate611(.a(G577), .O(gate188inter8));
  nand2 gate612(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate613(.a(s_9), .b(gate188inter3), .O(gate188inter10));
  nor2  gate614(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate615(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate616(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1639(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1640(.a(gate190inter0), .b(s_156), .O(gate190inter1));
  and2  gate1641(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1642(.a(s_156), .O(gate190inter3));
  inv1  gate1643(.a(s_157), .O(gate190inter4));
  nand2 gate1644(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1645(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1646(.a(G580), .O(gate190inter7));
  inv1  gate1647(.a(G581), .O(gate190inter8));
  nand2 gate1648(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1649(.a(s_157), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1650(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1651(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1652(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate995(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate996(.a(gate192inter0), .b(s_64), .O(gate192inter1));
  and2  gate997(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate998(.a(s_64), .O(gate192inter3));
  inv1  gate999(.a(s_65), .O(gate192inter4));
  nand2 gate1000(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1001(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1002(.a(G584), .O(gate192inter7));
  inv1  gate1003(.a(G585), .O(gate192inter8));
  nand2 gate1004(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1005(.a(s_65), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1006(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1007(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1008(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2605(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2606(.a(gate193inter0), .b(s_294), .O(gate193inter1));
  and2  gate2607(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2608(.a(s_294), .O(gate193inter3));
  inv1  gate2609(.a(s_295), .O(gate193inter4));
  nand2 gate2610(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2611(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2612(.a(G586), .O(gate193inter7));
  inv1  gate2613(.a(G587), .O(gate193inter8));
  nand2 gate2614(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2615(.a(s_295), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2616(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2617(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2618(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1387(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1388(.a(gate194inter0), .b(s_120), .O(gate194inter1));
  and2  gate1389(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1390(.a(s_120), .O(gate194inter3));
  inv1  gate1391(.a(s_121), .O(gate194inter4));
  nand2 gate1392(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1393(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1394(.a(G588), .O(gate194inter7));
  inv1  gate1395(.a(G589), .O(gate194inter8));
  nand2 gate1396(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1397(.a(s_121), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1398(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1399(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1400(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2423(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2424(.a(gate195inter0), .b(s_268), .O(gate195inter1));
  and2  gate2425(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2426(.a(s_268), .O(gate195inter3));
  inv1  gate2427(.a(s_269), .O(gate195inter4));
  nand2 gate2428(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2429(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2430(.a(G590), .O(gate195inter7));
  inv1  gate2431(.a(G591), .O(gate195inter8));
  nand2 gate2432(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2433(.a(s_269), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2434(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2435(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2436(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2185(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2186(.a(gate198inter0), .b(s_234), .O(gate198inter1));
  and2  gate2187(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2188(.a(s_234), .O(gate198inter3));
  inv1  gate2189(.a(s_235), .O(gate198inter4));
  nand2 gate2190(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2191(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2192(.a(G596), .O(gate198inter7));
  inv1  gate2193(.a(G597), .O(gate198inter8));
  nand2 gate2194(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2195(.a(s_235), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2196(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2197(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2198(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2227(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2228(.a(gate202inter0), .b(s_240), .O(gate202inter1));
  and2  gate2229(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2230(.a(s_240), .O(gate202inter3));
  inv1  gate2231(.a(s_241), .O(gate202inter4));
  nand2 gate2232(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2233(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2234(.a(G612), .O(gate202inter7));
  inv1  gate2235(.a(G617), .O(gate202inter8));
  nand2 gate2236(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2237(.a(s_241), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2238(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2239(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2240(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2115(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2116(.a(gate206inter0), .b(s_224), .O(gate206inter1));
  and2  gate2117(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2118(.a(s_224), .O(gate206inter3));
  inv1  gate2119(.a(s_225), .O(gate206inter4));
  nand2 gate2120(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2121(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2122(.a(G632), .O(gate206inter7));
  inv1  gate2123(.a(G637), .O(gate206inter8));
  nand2 gate2124(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2125(.a(s_225), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2126(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2127(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2128(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate729(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate730(.a(gate207inter0), .b(s_26), .O(gate207inter1));
  and2  gate731(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate732(.a(s_26), .O(gate207inter3));
  inv1  gate733(.a(s_27), .O(gate207inter4));
  nand2 gate734(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate735(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate736(.a(G622), .O(gate207inter7));
  inv1  gate737(.a(G632), .O(gate207inter8));
  nand2 gate738(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate739(.a(s_27), .b(gate207inter3), .O(gate207inter10));
  nor2  gate740(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate741(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate742(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1555(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1556(.a(gate212inter0), .b(s_144), .O(gate212inter1));
  and2  gate1557(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1558(.a(s_144), .O(gate212inter3));
  inv1  gate1559(.a(s_145), .O(gate212inter4));
  nand2 gate1560(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1561(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1562(.a(G617), .O(gate212inter7));
  inv1  gate1563(.a(G669), .O(gate212inter8));
  nand2 gate1564(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1565(.a(s_145), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1566(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1567(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1568(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate855(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate856(.a(gate213inter0), .b(s_44), .O(gate213inter1));
  and2  gate857(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate858(.a(s_44), .O(gate213inter3));
  inv1  gate859(.a(s_45), .O(gate213inter4));
  nand2 gate860(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate861(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate862(.a(G602), .O(gate213inter7));
  inv1  gate863(.a(G672), .O(gate213inter8));
  nand2 gate864(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate865(.a(s_45), .b(gate213inter3), .O(gate213inter10));
  nor2  gate866(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate867(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate868(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1513(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1514(.a(gate217inter0), .b(s_138), .O(gate217inter1));
  and2  gate1515(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1516(.a(s_138), .O(gate217inter3));
  inv1  gate1517(.a(s_139), .O(gate217inter4));
  nand2 gate1518(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1519(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1520(.a(G622), .O(gate217inter7));
  inv1  gate1521(.a(G678), .O(gate217inter8));
  nand2 gate1522(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1523(.a(s_139), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1524(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1525(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1526(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2213(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2214(.a(gate220inter0), .b(s_238), .O(gate220inter1));
  and2  gate2215(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2216(.a(s_238), .O(gate220inter3));
  inv1  gate2217(.a(s_239), .O(gate220inter4));
  nand2 gate2218(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2219(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2220(.a(G637), .O(gate220inter7));
  inv1  gate2221(.a(G681), .O(gate220inter8));
  nand2 gate2222(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2223(.a(s_239), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2224(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2225(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2226(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1331(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1332(.a(gate227inter0), .b(s_112), .O(gate227inter1));
  and2  gate1333(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1334(.a(s_112), .O(gate227inter3));
  inv1  gate1335(.a(s_113), .O(gate227inter4));
  nand2 gate1336(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1337(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1338(.a(G694), .O(gate227inter7));
  inv1  gate1339(.a(G695), .O(gate227inter8));
  nand2 gate1340(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1341(.a(s_113), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1342(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1343(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1344(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1485(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1486(.a(gate229inter0), .b(s_134), .O(gate229inter1));
  and2  gate1487(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1488(.a(s_134), .O(gate229inter3));
  inv1  gate1489(.a(s_135), .O(gate229inter4));
  nand2 gate1490(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1491(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1492(.a(G698), .O(gate229inter7));
  inv1  gate1493(.a(G699), .O(gate229inter8));
  nand2 gate1494(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1495(.a(s_135), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1496(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1497(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1498(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1835(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1836(.a(gate231inter0), .b(s_184), .O(gate231inter1));
  and2  gate1837(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1838(.a(s_184), .O(gate231inter3));
  inv1  gate1839(.a(s_185), .O(gate231inter4));
  nand2 gate1840(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1841(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1842(.a(G702), .O(gate231inter7));
  inv1  gate1843(.a(G703), .O(gate231inter8));
  nand2 gate1844(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1845(.a(s_185), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1846(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1847(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1848(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate631(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate632(.a(gate235inter0), .b(s_12), .O(gate235inter1));
  and2  gate633(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate634(.a(s_12), .O(gate235inter3));
  inv1  gate635(.a(s_13), .O(gate235inter4));
  nand2 gate636(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate637(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate638(.a(G248), .O(gate235inter7));
  inv1  gate639(.a(G724), .O(gate235inter8));
  nand2 gate640(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate641(.a(s_13), .b(gate235inter3), .O(gate235inter10));
  nor2  gate642(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate643(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate644(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2283(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2284(.a(gate240inter0), .b(s_248), .O(gate240inter1));
  and2  gate2285(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2286(.a(s_248), .O(gate240inter3));
  inv1  gate2287(.a(s_249), .O(gate240inter4));
  nand2 gate2288(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2289(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2290(.a(G263), .O(gate240inter7));
  inv1  gate2291(.a(G715), .O(gate240inter8));
  nand2 gate2292(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2293(.a(s_249), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2294(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2295(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2296(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2045(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2046(.a(gate242inter0), .b(s_214), .O(gate242inter1));
  and2  gate2047(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2048(.a(s_214), .O(gate242inter3));
  inv1  gate2049(.a(s_215), .O(gate242inter4));
  nand2 gate2050(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2051(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2052(.a(G718), .O(gate242inter7));
  inv1  gate2053(.a(G730), .O(gate242inter8));
  nand2 gate2054(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2055(.a(s_215), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2056(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2057(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2058(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1065(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1066(.a(gate243inter0), .b(s_74), .O(gate243inter1));
  and2  gate1067(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1068(.a(s_74), .O(gate243inter3));
  inv1  gate1069(.a(s_75), .O(gate243inter4));
  nand2 gate1070(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1071(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1072(.a(G245), .O(gate243inter7));
  inv1  gate1073(.a(G733), .O(gate243inter8));
  nand2 gate1074(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1075(.a(s_75), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1076(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1077(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1078(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1009(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1010(.a(gate244inter0), .b(s_66), .O(gate244inter1));
  and2  gate1011(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1012(.a(s_66), .O(gate244inter3));
  inv1  gate1013(.a(s_67), .O(gate244inter4));
  nand2 gate1014(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1015(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1016(.a(G721), .O(gate244inter7));
  inv1  gate1017(.a(G733), .O(gate244inter8));
  nand2 gate1018(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1019(.a(s_67), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1020(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1021(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1022(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate967(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate968(.a(gate245inter0), .b(s_60), .O(gate245inter1));
  and2  gate969(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate970(.a(s_60), .O(gate245inter3));
  inv1  gate971(.a(s_61), .O(gate245inter4));
  nand2 gate972(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate973(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate974(.a(G248), .O(gate245inter7));
  inv1  gate975(.a(G736), .O(gate245inter8));
  nand2 gate976(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate977(.a(s_61), .b(gate245inter3), .O(gate245inter10));
  nor2  gate978(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate979(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate980(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1667(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1668(.a(gate246inter0), .b(s_160), .O(gate246inter1));
  and2  gate1669(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1670(.a(s_160), .O(gate246inter3));
  inv1  gate1671(.a(s_161), .O(gate246inter4));
  nand2 gate1672(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1673(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1674(.a(G724), .O(gate246inter7));
  inv1  gate1675(.a(G736), .O(gate246inter8));
  nand2 gate1676(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1677(.a(s_161), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1678(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1679(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1680(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1233(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1234(.a(gate247inter0), .b(s_98), .O(gate247inter1));
  and2  gate1235(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1236(.a(s_98), .O(gate247inter3));
  inv1  gate1237(.a(s_99), .O(gate247inter4));
  nand2 gate1238(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1239(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1240(.a(G251), .O(gate247inter7));
  inv1  gate1241(.a(G739), .O(gate247inter8));
  nand2 gate1242(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1243(.a(s_99), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1244(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1245(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1246(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate715(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate716(.a(gate248inter0), .b(s_24), .O(gate248inter1));
  and2  gate717(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate718(.a(s_24), .O(gate248inter3));
  inv1  gate719(.a(s_25), .O(gate248inter4));
  nand2 gate720(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate721(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate722(.a(G727), .O(gate248inter7));
  inv1  gate723(.a(G739), .O(gate248inter8));
  nand2 gate724(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate725(.a(s_25), .b(gate248inter3), .O(gate248inter10));
  nor2  gate726(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate727(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate728(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1275(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1276(.a(gate249inter0), .b(s_104), .O(gate249inter1));
  and2  gate1277(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1278(.a(s_104), .O(gate249inter3));
  inv1  gate1279(.a(s_105), .O(gate249inter4));
  nand2 gate1280(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1281(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1282(.a(G254), .O(gate249inter7));
  inv1  gate1283(.a(G742), .O(gate249inter8));
  nand2 gate1284(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1285(.a(s_105), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1286(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1287(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1288(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2619(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2620(.a(gate252inter0), .b(s_296), .O(gate252inter1));
  and2  gate2621(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2622(.a(s_296), .O(gate252inter3));
  inv1  gate2623(.a(s_297), .O(gate252inter4));
  nand2 gate2624(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2625(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2626(.a(G709), .O(gate252inter7));
  inv1  gate2627(.a(G745), .O(gate252inter8));
  nand2 gate2628(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2629(.a(s_297), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2630(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2631(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2632(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate1989(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1990(.a(gate253inter0), .b(s_206), .O(gate253inter1));
  and2  gate1991(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1992(.a(s_206), .O(gate253inter3));
  inv1  gate1993(.a(s_207), .O(gate253inter4));
  nand2 gate1994(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1995(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1996(.a(G260), .O(gate253inter7));
  inv1  gate1997(.a(G748), .O(gate253inter8));
  nand2 gate1998(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1999(.a(s_207), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2000(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2001(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2002(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1737(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1738(.a(gate255inter0), .b(s_170), .O(gate255inter1));
  and2  gate1739(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1740(.a(s_170), .O(gate255inter3));
  inv1  gate1741(.a(s_171), .O(gate255inter4));
  nand2 gate1742(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1743(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1744(.a(G263), .O(gate255inter7));
  inv1  gate1745(.a(G751), .O(gate255inter8));
  nand2 gate1746(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1747(.a(s_171), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1748(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1749(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1750(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1107(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1108(.a(gate256inter0), .b(s_80), .O(gate256inter1));
  and2  gate1109(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1110(.a(s_80), .O(gate256inter3));
  inv1  gate1111(.a(s_81), .O(gate256inter4));
  nand2 gate1112(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1113(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1114(.a(G715), .O(gate256inter7));
  inv1  gate1115(.a(G751), .O(gate256inter8));
  nand2 gate1116(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1117(.a(s_81), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1118(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1119(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1120(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1975(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1976(.a(gate259inter0), .b(s_204), .O(gate259inter1));
  and2  gate1977(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1978(.a(s_204), .O(gate259inter3));
  inv1  gate1979(.a(s_205), .O(gate259inter4));
  nand2 gate1980(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1981(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1982(.a(G758), .O(gate259inter7));
  inv1  gate1983(.a(G759), .O(gate259inter8));
  nand2 gate1984(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1985(.a(s_205), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1986(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1987(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1988(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1037(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1038(.a(gate262inter0), .b(s_70), .O(gate262inter1));
  and2  gate1039(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1040(.a(s_70), .O(gate262inter3));
  inv1  gate1041(.a(s_71), .O(gate262inter4));
  nand2 gate1042(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1043(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1044(.a(G764), .O(gate262inter7));
  inv1  gate1045(.a(G765), .O(gate262inter8));
  nand2 gate1046(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1047(.a(s_71), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1048(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1049(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1050(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2325(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2326(.a(gate263inter0), .b(s_254), .O(gate263inter1));
  and2  gate2327(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2328(.a(s_254), .O(gate263inter3));
  inv1  gate2329(.a(s_255), .O(gate263inter4));
  nand2 gate2330(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2331(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2332(.a(G766), .O(gate263inter7));
  inv1  gate2333(.a(G767), .O(gate263inter8));
  nand2 gate2334(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2335(.a(s_255), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2336(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2337(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2338(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2129(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2130(.a(gate264inter0), .b(s_226), .O(gate264inter1));
  and2  gate2131(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2132(.a(s_226), .O(gate264inter3));
  inv1  gate2133(.a(s_227), .O(gate264inter4));
  nand2 gate2134(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2135(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2136(.a(G768), .O(gate264inter7));
  inv1  gate2137(.a(G769), .O(gate264inter8));
  nand2 gate2138(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2139(.a(s_227), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2140(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2141(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2142(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate2381(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2382(.a(gate265inter0), .b(s_262), .O(gate265inter1));
  and2  gate2383(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2384(.a(s_262), .O(gate265inter3));
  inv1  gate2385(.a(s_263), .O(gate265inter4));
  nand2 gate2386(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2387(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2388(.a(G642), .O(gate265inter7));
  inv1  gate2389(.a(G770), .O(gate265inter8));
  nand2 gate2390(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2391(.a(s_263), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2392(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2393(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2394(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate785(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate786(.a(gate266inter0), .b(s_34), .O(gate266inter1));
  and2  gate787(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate788(.a(s_34), .O(gate266inter3));
  inv1  gate789(.a(s_35), .O(gate266inter4));
  nand2 gate790(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate791(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate792(.a(G645), .O(gate266inter7));
  inv1  gate793(.a(G773), .O(gate266inter8));
  nand2 gate794(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate795(.a(s_35), .b(gate266inter3), .O(gate266inter10));
  nor2  gate796(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate797(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate798(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1681(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1682(.a(gate268inter0), .b(s_162), .O(gate268inter1));
  and2  gate1683(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1684(.a(s_162), .O(gate268inter3));
  inv1  gate1685(.a(s_163), .O(gate268inter4));
  nand2 gate1686(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1687(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1688(.a(G651), .O(gate268inter7));
  inv1  gate1689(.a(G779), .O(gate268inter8));
  nand2 gate1690(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1691(.a(s_163), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1692(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1693(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1694(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1373(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1374(.a(gate269inter0), .b(s_118), .O(gate269inter1));
  and2  gate1375(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1376(.a(s_118), .O(gate269inter3));
  inv1  gate1377(.a(s_119), .O(gate269inter4));
  nand2 gate1378(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1379(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1380(.a(G654), .O(gate269inter7));
  inv1  gate1381(.a(G782), .O(gate269inter8));
  nand2 gate1382(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1383(.a(s_119), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1384(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1385(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1386(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate2675(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2676(.a(gate270inter0), .b(s_304), .O(gate270inter1));
  and2  gate2677(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2678(.a(s_304), .O(gate270inter3));
  inv1  gate2679(.a(s_305), .O(gate270inter4));
  nand2 gate2680(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2681(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2682(.a(G657), .O(gate270inter7));
  inv1  gate2683(.a(G785), .O(gate270inter8));
  nand2 gate2684(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2685(.a(s_305), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2686(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2687(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2688(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2143(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2144(.a(gate271inter0), .b(s_228), .O(gate271inter1));
  and2  gate2145(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2146(.a(s_228), .O(gate271inter3));
  inv1  gate2147(.a(s_229), .O(gate271inter4));
  nand2 gate2148(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2149(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2150(.a(G660), .O(gate271inter7));
  inv1  gate2151(.a(G788), .O(gate271inter8));
  nand2 gate2152(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2153(.a(s_229), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2154(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2155(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2156(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2339(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2340(.a(gate272inter0), .b(s_256), .O(gate272inter1));
  and2  gate2341(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2342(.a(s_256), .O(gate272inter3));
  inv1  gate2343(.a(s_257), .O(gate272inter4));
  nand2 gate2344(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2345(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2346(.a(G663), .O(gate272inter7));
  inv1  gate2347(.a(G791), .O(gate272inter8));
  nand2 gate2348(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2349(.a(s_257), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2350(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2351(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2352(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate813(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate814(.a(gate273inter0), .b(s_38), .O(gate273inter1));
  and2  gate815(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate816(.a(s_38), .O(gate273inter3));
  inv1  gate817(.a(s_39), .O(gate273inter4));
  nand2 gate818(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate819(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate820(.a(G642), .O(gate273inter7));
  inv1  gate821(.a(G794), .O(gate273inter8));
  nand2 gate822(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate823(.a(s_39), .b(gate273inter3), .O(gate273inter10));
  nor2  gate824(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate825(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate826(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2073(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2074(.a(gate282inter0), .b(s_218), .O(gate282inter1));
  and2  gate2075(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2076(.a(s_218), .O(gate282inter3));
  inv1  gate2077(.a(s_219), .O(gate282inter4));
  nand2 gate2078(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2079(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2080(.a(G782), .O(gate282inter7));
  inv1  gate2081(.a(G806), .O(gate282inter8));
  nand2 gate2082(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2083(.a(s_219), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2084(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2085(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2086(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1919(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1920(.a(gate283inter0), .b(s_196), .O(gate283inter1));
  and2  gate1921(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1922(.a(s_196), .O(gate283inter3));
  inv1  gate1923(.a(s_197), .O(gate283inter4));
  nand2 gate1924(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1925(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1926(.a(G657), .O(gate283inter7));
  inv1  gate1927(.a(G809), .O(gate283inter8));
  nand2 gate1928(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1929(.a(s_197), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1930(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1931(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1932(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2171(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2172(.a(gate291inter0), .b(s_232), .O(gate291inter1));
  and2  gate2173(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2174(.a(s_232), .O(gate291inter3));
  inv1  gate2175(.a(s_233), .O(gate291inter4));
  nand2 gate2176(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2177(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2178(.a(G822), .O(gate291inter7));
  inv1  gate2179(.a(G823), .O(gate291inter8));
  nand2 gate2180(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2181(.a(s_233), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2182(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2183(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2184(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1415(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1416(.a(gate389inter0), .b(s_124), .O(gate389inter1));
  and2  gate1417(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1418(.a(s_124), .O(gate389inter3));
  inv1  gate1419(.a(s_125), .O(gate389inter4));
  nand2 gate1420(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1421(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1422(.a(G3), .O(gate389inter7));
  inv1  gate1423(.a(G1042), .O(gate389inter8));
  nand2 gate1424(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1425(.a(s_125), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1426(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1427(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1428(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1765(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1766(.a(gate391inter0), .b(s_174), .O(gate391inter1));
  and2  gate1767(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1768(.a(s_174), .O(gate391inter3));
  inv1  gate1769(.a(s_175), .O(gate391inter4));
  nand2 gate1770(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1771(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1772(.a(G5), .O(gate391inter7));
  inv1  gate1773(.a(G1048), .O(gate391inter8));
  nand2 gate1774(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1775(.a(s_175), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1776(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1777(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1778(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1947(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1948(.a(gate394inter0), .b(s_200), .O(gate394inter1));
  and2  gate1949(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1950(.a(s_200), .O(gate394inter3));
  inv1  gate1951(.a(s_201), .O(gate394inter4));
  nand2 gate1952(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1953(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1954(.a(G8), .O(gate394inter7));
  inv1  gate1955(.a(G1057), .O(gate394inter8));
  nand2 gate1956(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1957(.a(s_201), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1958(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1959(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1960(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1135(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1136(.a(gate396inter0), .b(s_84), .O(gate396inter1));
  and2  gate1137(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1138(.a(s_84), .O(gate396inter3));
  inv1  gate1139(.a(s_85), .O(gate396inter4));
  nand2 gate1140(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1141(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1142(.a(G10), .O(gate396inter7));
  inv1  gate1143(.a(G1063), .O(gate396inter8));
  nand2 gate1144(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1145(.a(s_85), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1146(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1147(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1148(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2591(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2592(.a(gate400inter0), .b(s_292), .O(gate400inter1));
  and2  gate2593(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2594(.a(s_292), .O(gate400inter3));
  inv1  gate2595(.a(s_293), .O(gate400inter4));
  nand2 gate2596(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2597(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2598(.a(G14), .O(gate400inter7));
  inv1  gate2599(.a(G1075), .O(gate400inter8));
  nand2 gate2600(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2601(.a(s_293), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2602(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2603(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2604(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate925(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate926(.a(gate402inter0), .b(s_54), .O(gate402inter1));
  and2  gate927(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate928(.a(s_54), .O(gate402inter3));
  inv1  gate929(.a(s_55), .O(gate402inter4));
  nand2 gate930(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate931(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate932(.a(G16), .O(gate402inter7));
  inv1  gate933(.a(G1081), .O(gate402inter8));
  nand2 gate934(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate935(.a(s_55), .b(gate402inter3), .O(gate402inter10));
  nor2  gate936(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate937(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate938(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate659(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate660(.a(gate403inter0), .b(s_16), .O(gate403inter1));
  and2  gate661(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate662(.a(s_16), .O(gate403inter3));
  inv1  gate663(.a(s_17), .O(gate403inter4));
  nand2 gate664(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate665(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate666(.a(G17), .O(gate403inter7));
  inv1  gate667(.a(G1084), .O(gate403inter8));
  nand2 gate668(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate669(.a(s_17), .b(gate403inter3), .O(gate403inter10));
  nor2  gate670(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate671(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate672(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate2031(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2032(.a(gate404inter0), .b(s_212), .O(gate404inter1));
  and2  gate2033(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2034(.a(s_212), .O(gate404inter3));
  inv1  gate2035(.a(s_213), .O(gate404inter4));
  nand2 gate2036(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2037(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2038(.a(G18), .O(gate404inter7));
  inv1  gate2039(.a(G1087), .O(gate404inter8));
  nand2 gate2040(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2041(.a(s_213), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2042(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2043(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2044(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate953(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate954(.a(gate405inter0), .b(s_58), .O(gate405inter1));
  and2  gate955(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate956(.a(s_58), .O(gate405inter3));
  inv1  gate957(.a(s_59), .O(gate405inter4));
  nand2 gate958(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate959(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate960(.a(G19), .O(gate405inter7));
  inv1  gate961(.a(G1090), .O(gate405inter8));
  nand2 gate962(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate963(.a(s_59), .b(gate405inter3), .O(gate405inter10));
  nor2  gate964(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate965(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate966(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1317(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1318(.a(gate407inter0), .b(s_110), .O(gate407inter1));
  and2  gate1319(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1320(.a(s_110), .O(gate407inter3));
  inv1  gate1321(.a(s_111), .O(gate407inter4));
  nand2 gate1322(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1323(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1324(.a(G21), .O(gate407inter7));
  inv1  gate1325(.a(G1096), .O(gate407inter8));
  nand2 gate1326(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1327(.a(s_111), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1328(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1329(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1330(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2661(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2662(.a(gate409inter0), .b(s_302), .O(gate409inter1));
  and2  gate2663(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2664(.a(s_302), .O(gate409inter3));
  inv1  gate2665(.a(s_303), .O(gate409inter4));
  nand2 gate2666(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2667(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2668(.a(G23), .O(gate409inter7));
  inv1  gate2669(.a(G1102), .O(gate409inter8));
  nand2 gate2670(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2671(.a(s_303), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2672(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2673(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2674(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate911(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate912(.a(gate416inter0), .b(s_52), .O(gate416inter1));
  and2  gate913(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate914(.a(s_52), .O(gate416inter3));
  inv1  gate915(.a(s_53), .O(gate416inter4));
  nand2 gate916(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate917(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate918(.a(G30), .O(gate416inter7));
  inv1  gate919(.a(G1123), .O(gate416inter8));
  nand2 gate920(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate921(.a(s_53), .b(gate416inter3), .O(gate416inter10));
  nor2  gate922(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate923(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate924(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2535(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2536(.a(gate417inter0), .b(s_284), .O(gate417inter1));
  and2  gate2537(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2538(.a(s_284), .O(gate417inter3));
  inv1  gate2539(.a(s_285), .O(gate417inter4));
  nand2 gate2540(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2541(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2542(.a(G31), .O(gate417inter7));
  inv1  gate2543(.a(G1126), .O(gate417inter8));
  nand2 gate2544(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2545(.a(s_285), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2546(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2547(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2548(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1961(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1962(.a(gate419inter0), .b(s_202), .O(gate419inter1));
  and2  gate1963(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1964(.a(s_202), .O(gate419inter3));
  inv1  gate1965(.a(s_203), .O(gate419inter4));
  nand2 gate1966(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1967(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1968(.a(G1), .O(gate419inter7));
  inv1  gate1969(.a(G1132), .O(gate419inter8));
  nand2 gate1970(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1971(.a(s_203), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1972(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1973(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1974(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2465(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2466(.a(gate429inter0), .b(s_274), .O(gate429inter1));
  and2  gate2467(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2468(.a(s_274), .O(gate429inter3));
  inv1  gate2469(.a(s_275), .O(gate429inter4));
  nand2 gate2470(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2471(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2472(.a(G6), .O(gate429inter7));
  inv1  gate2473(.a(G1147), .O(gate429inter8));
  nand2 gate2474(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2475(.a(s_275), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2476(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2477(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2478(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2241(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2242(.a(gate431inter0), .b(s_242), .O(gate431inter1));
  and2  gate2243(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2244(.a(s_242), .O(gate431inter3));
  inv1  gate2245(.a(s_243), .O(gate431inter4));
  nand2 gate2246(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2247(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2248(.a(G7), .O(gate431inter7));
  inv1  gate2249(.a(G1150), .O(gate431inter8));
  nand2 gate2250(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2251(.a(s_243), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2252(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2253(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2254(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate897(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate898(.a(gate435inter0), .b(s_50), .O(gate435inter1));
  and2  gate899(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate900(.a(s_50), .O(gate435inter3));
  inv1  gate901(.a(s_51), .O(gate435inter4));
  nand2 gate902(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate903(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate904(.a(G9), .O(gate435inter7));
  inv1  gate905(.a(G1156), .O(gate435inter8));
  nand2 gate906(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate907(.a(s_51), .b(gate435inter3), .O(gate435inter10));
  nor2  gate908(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate909(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate910(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate757(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate758(.a(gate436inter0), .b(s_30), .O(gate436inter1));
  and2  gate759(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate760(.a(s_30), .O(gate436inter3));
  inv1  gate761(.a(s_31), .O(gate436inter4));
  nand2 gate762(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate763(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate764(.a(G1060), .O(gate436inter7));
  inv1  gate765(.a(G1156), .O(gate436inter8));
  nand2 gate766(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate767(.a(s_31), .b(gate436inter3), .O(gate436inter10));
  nor2  gate768(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate769(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate770(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1079(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1080(.a(gate438inter0), .b(s_76), .O(gate438inter1));
  and2  gate1081(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1082(.a(s_76), .O(gate438inter3));
  inv1  gate1083(.a(s_77), .O(gate438inter4));
  nand2 gate1084(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1085(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1086(.a(G1063), .O(gate438inter7));
  inv1  gate1087(.a(G1159), .O(gate438inter8));
  nand2 gate1088(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1089(.a(s_77), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1090(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1091(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1092(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1289(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1290(.a(gate440inter0), .b(s_106), .O(gate440inter1));
  and2  gate1291(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1292(.a(s_106), .O(gate440inter3));
  inv1  gate1293(.a(s_107), .O(gate440inter4));
  nand2 gate1294(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1295(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1296(.a(G1066), .O(gate440inter7));
  inv1  gate1297(.a(G1162), .O(gate440inter8));
  nand2 gate1298(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1299(.a(s_107), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1300(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1301(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1302(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1261(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1262(.a(gate443inter0), .b(s_102), .O(gate443inter1));
  and2  gate1263(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1264(.a(s_102), .O(gate443inter3));
  inv1  gate1265(.a(s_103), .O(gate443inter4));
  nand2 gate1266(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1267(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1268(.a(G13), .O(gate443inter7));
  inv1  gate1269(.a(G1168), .O(gate443inter8));
  nand2 gate1270(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1271(.a(s_103), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1272(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1273(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1274(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1163(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1164(.a(gate447inter0), .b(s_88), .O(gate447inter1));
  and2  gate1165(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1166(.a(s_88), .O(gate447inter3));
  inv1  gate1167(.a(s_89), .O(gate447inter4));
  nand2 gate1168(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1169(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1170(.a(G15), .O(gate447inter7));
  inv1  gate1171(.a(G1174), .O(gate447inter8));
  nand2 gate1172(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1173(.a(s_89), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1174(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1175(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1176(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1471(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1472(.a(gate448inter0), .b(s_132), .O(gate448inter1));
  and2  gate1473(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1474(.a(s_132), .O(gate448inter3));
  inv1  gate1475(.a(s_133), .O(gate448inter4));
  nand2 gate1476(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1477(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1478(.a(G1078), .O(gate448inter7));
  inv1  gate1479(.a(G1174), .O(gate448inter8));
  nand2 gate1480(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1481(.a(s_133), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1482(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1483(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1484(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1093(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1094(.a(gate451inter0), .b(s_78), .O(gate451inter1));
  and2  gate1095(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1096(.a(s_78), .O(gate451inter3));
  inv1  gate1097(.a(s_79), .O(gate451inter4));
  nand2 gate1098(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1099(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1100(.a(G17), .O(gate451inter7));
  inv1  gate1101(.a(G1180), .O(gate451inter8));
  nand2 gate1102(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1103(.a(s_79), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1104(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1105(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1106(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate981(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate982(.a(gate452inter0), .b(s_62), .O(gate452inter1));
  and2  gate983(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate984(.a(s_62), .O(gate452inter3));
  inv1  gate985(.a(s_63), .O(gate452inter4));
  nand2 gate986(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate987(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate988(.a(G1084), .O(gate452inter7));
  inv1  gate989(.a(G1180), .O(gate452inter8));
  nand2 gate990(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate991(.a(s_63), .b(gate452inter3), .O(gate452inter10));
  nor2  gate992(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate993(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate994(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2311(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2312(.a(gate456inter0), .b(s_252), .O(gate456inter1));
  and2  gate2313(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2314(.a(s_252), .O(gate456inter3));
  inv1  gate2315(.a(s_253), .O(gate456inter4));
  nand2 gate2316(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2317(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2318(.a(G1090), .O(gate456inter7));
  inv1  gate2319(.a(G1186), .O(gate456inter8));
  nand2 gate2320(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2321(.a(s_253), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2322(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2323(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2324(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2199(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2200(.a(gate463inter0), .b(s_236), .O(gate463inter1));
  and2  gate2201(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2202(.a(s_236), .O(gate463inter3));
  inv1  gate2203(.a(s_237), .O(gate463inter4));
  nand2 gate2204(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2205(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2206(.a(G23), .O(gate463inter7));
  inv1  gate2207(.a(G1198), .O(gate463inter8));
  nand2 gate2208(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2209(.a(s_237), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2210(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2211(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2212(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1625(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1626(.a(gate464inter0), .b(s_154), .O(gate464inter1));
  and2  gate1627(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1628(.a(s_154), .O(gate464inter3));
  inv1  gate1629(.a(s_155), .O(gate464inter4));
  nand2 gate1630(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1631(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1632(.a(G1102), .O(gate464inter7));
  inv1  gate1633(.a(G1198), .O(gate464inter8));
  nand2 gate1634(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1635(.a(s_155), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1636(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1637(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1638(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1569(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1570(.a(gate468inter0), .b(s_146), .O(gate468inter1));
  and2  gate1571(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1572(.a(s_146), .O(gate468inter3));
  inv1  gate1573(.a(s_147), .O(gate468inter4));
  nand2 gate1574(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1575(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1576(.a(G1108), .O(gate468inter7));
  inv1  gate1577(.a(G1204), .O(gate468inter8));
  nand2 gate1578(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1579(.a(s_147), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1580(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1581(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1582(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate617(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate618(.a(gate472inter0), .b(s_10), .O(gate472inter1));
  and2  gate619(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate620(.a(s_10), .O(gate472inter3));
  inv1  gate621(.a(s_11), .O(gate472inter4));
  nand2 gate622(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate623(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate624(.a(G1114), .O(gate472inter7));
  inv1  gate625(.a(G1210), .O(gate472inter8));
  nand2 gate626(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate627(.a(s_11), .b(gate472inter3), .O(gate472inter10));
  nor2  gate628(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate629(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate630(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2647(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2648(.a(gate476inter0), .b(s_300), .O(gate476inter1));
  and2  gate2649(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2650(.a(s_300), .O(gate476inter3));
  inv1  gate2651(.a(s_301), .O(gate476inter4));
  nand2 gate2652(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2653(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2654(.a(G1120), .O(gate476inter7));
  inv1  gate2655(.a(G1216), .O(gate476inter8));
  nand2 gate2656(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2657(.a(s_301), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2658(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2659(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2660(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate771(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate772(.a(gate477inter0), .b(s_32), .O(gate477inter1));
  and2  gate773(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate774(.a(s_32), .O(gate477inter3));
  inv1  gate775(.a(s_33), .O(gate477inter4));
  nand2 gate776(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate777(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate778(.a(G30), .O(gate477inter7));
  inv1  gate779(.a(G1219), .O(gate477inter8));
  nand2 gate780(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate781(.a(s_33), .b(gate477inter3), .O(gate477inter10));
  nor2  gate782(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate783(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate784(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1891(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1892(.a(gate478inter0), .b(s_192), .O(gate478inter1));
  and2  gate1893(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1894(.a(s_192), .O(gate478inter3));
  inv1  gate1895(.a(s_193), .O(gate478inter4));
  nand2 gate1896(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1897(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1898(.a(G1123), .O(gate478inter7));
  inv1  gate1899(.a(G1219), .O(gate478inter8));
  nand2 gate1900(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1901(.a(s_193), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1902(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1903(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1904(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1345(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1346(.a(gate482inter0), .b(s_114), .O(gate482inter1));
  and2  gate1347(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1348(.a(s_114), .O(gate482inter3));
  inv1  gate1349(.a(s_115), .O(gate482inter4));
  nand2 gate1350(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1351(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1352(.a(G1129), .O(gate482inter7));
  inv1  gate1353(.a(G1225), .O(gate482inter8));
  nand2 gate1354(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1355(.a(s_115), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1356(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1357(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1358(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1219(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1220(.a(gate486inter0), .b(s_96), .O(gate486inter1));
  and2  gate1221(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1222(.a(s_96), .O(gate486inter3));
  inv1  gate1223(.a(s_97), .O(gate486inter4));
  nand2 gate1224(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1225(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1226(.a(G1234), .O(gate486inter7));
  inv1  gate1227(.a(G1235), .O(gate486inter8));
  nand2 gate1228(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1229(.a(s_97), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1230(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1231(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1232(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2409(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2410(.a(gate488inter0), .b(s_266), .O(gate488inter1));
  and2  gate2411(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2412(.a(s_266), .O(gate488inter3));
  inv1  gate2413(.a(s_267), .O(gate488inter4));
  nand2 gate2414(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2415(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2416(.a(G1238), .O(gate488inter7));
  inv1  gate2417(.a(G1239), .O(gate488inter8));
  nand2 gate2418(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2419(.a(s_267), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2420(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2421(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2422(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2087(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2088(.a(gate492inter0), .b(s_220), .O(gate492inter1));
  and2  gate2089(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2090(.a(s_220), .O(gate492inter3));
  inv1  gate2091(.a(s_221), .O(gate492inter4));
  nand2 gate2092(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2093(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2094(.a(G1246), .O(gate492inter7));
  inv1  gate2095(.a(G1247), .O(gate492inter8));
  nand2 gate2096(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2097(.a(s_221), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2098(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2099(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2100(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1849(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1850(.a(gate495inter0), .b(s_186), .O(gate495inter1));
  and2  gate1851(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1852(.a(s_186), .O(gate495inter3));
  inv1  gate1853(.a(s_187), .O(gate495inter4));
  nand2 gate1854(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1855(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1856(.a(G1252), .O(gate495inter7));
  inv1  gate1857(.a(G1253), .O(gate495inter8));
  nand2 gate1858(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1859(.a(s_187), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1860(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1861(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1862(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate1611(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1612(.a(gate496inter0), .b(s_152), .O(gate496inter1));
  and2  gate1613(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1614(.a(s_152), .O(gate496inter3));
  inv1  gate1615(.a(s_153), .O(gate496inter4));
  nand2 gate1616(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1617(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1618(.a(G1254), .O(gate496inter7));
  inv1  gate1619(.a(G1255), .O(gate496inter8));
  nand2 gate1620(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1621(.a(s_153), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1622(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1623(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1624(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate2157(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2158(.a(gate497inter0), .b(s_230), .O(gate497inter1));
  and2  gate2159(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2160(.a(s_230), .O(gate497inter3));
  inv1  gate2161(.a(s_231), .O(gate497inter4));
  nand2 gate2162(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2163(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2164(.a(G1256), .O(gate497inter7));
  inv1  gate2165(.a(G1257), .O(gate497inter8));
  nand2 gate2166(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2167(.a(s_231), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2168(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2169(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2170(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2479(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2480(.a(gate499inter0), .b(s_276), .O(gate499inter1));
  and2  gate2481(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2482(.a(s_276), .O(gate499inter3));
  inv1  gate2483(.a(s_277), .O(gate499inter4));
  nand2 gate2484(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2485(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2486(.a(G1260), .O(gate499inter7));
  inv1  gate2487(.a(G1261), .O(gate499inter8));
  nand2 gate2488(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2489(.a(s_277), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2490(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2491(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2492(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2493(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2494(.a(gate505inter0), .b(s_278), .O(gate505inter1));
  and2  gate2495(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2496(.a(s_278), .O(gate505inter3));
  inv1  gate2497(.a(s_279), .O(gate505inter4));
  nand2 gate2498(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2499(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2500(.a(G1272), .O(gate505inter7));
  inv1  gate2501(.a(G1273), .O(gate505inter8));
  nand2 gate2502(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2503(.a(s_279), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2504(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2505(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2506(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2353(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2354(.a(gate509inter0), .b(s_258), .O(gate509inter1));
  and2  gate2355(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2356(.a(s_258), .O(gate509inter3));
  inv1  gate2357(.a(s_259), .O(gate509inter4));
  nand2 gate2358(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2359(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2360(.a(G1280), .O(gate509inter7));
  inv1  gate2361(.a(G1281), .O(gate509inter8));
  nand2 gate2362(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2363(.a(s_259), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2364(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2365(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2366(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1821(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1822(.a(gate511inter0), .b(s_182), .O(gate511inter1));
  and2  gate1823(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1824(.a(s_182), .O(gate511inter3));
  inv1  gate1825(.a(s_183), .O(gate511inter4));
  nand2 gate1826(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1827(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1828(.a(G1284), .O(gate511inter7));
  inv1  gate1829(.a(G1285), .O(gate511inter8));
  nand2 gate1830(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1831(.a(s_183), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1832(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1833(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1834(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1457(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1458(.a(gate514inter0), .b(s_130), .O(gate514inter1));
  and2  gate1459(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1460(.a(s_130), .O(gate514inter3));
  inv1  gate1461(.a(s_131), .O(gate514inter4));
  nand2 gate1462(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1463(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1464(.a(G1290), .O(gate514inter7));
  inv1  gate1465(.a(G1291), .O(gate514inter8));
  nand2 gate1466(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1467(.a(s_131), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1468(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1469(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1470(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule