module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1933(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1934(.a(gate11inter0), .b(s_198), .O(gate11inter1));
  and2  gate1935(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1936(.a(s_198), .O(gate11inter3));
  inv1  gate1937(.a(s_199), .O(gate11inter4));
  nand2 gate1938(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1939(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1940(.a(G5), .O(gate11inter7));
  inv1  gate1941(.a(G6), .O(gate11inter8));
  nand2 gate1942(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1943(.a(s_199), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1944(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1945(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1946(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1191(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1192(.a(gate18inter0), .b(s_92), .O(gate18inter1));
  and2  gate1193(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1194(.a(s_92), .O(gate18inter3));
  inv1  gate1195(.a(s_93), .O(gate18inter4));
  nand2 gate1196(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1197(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1198(.a(G19), .O(gate18inter7));
  inv1  gate1199(.a(G20), .O(gate18inter8));
  nand2 gate1200(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1201(.a(s_93), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1202(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1203(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1204(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1121(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1122(.a(gate22inter0), .b(s_82), .O(gate22inter1));
  and2  gate1123(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1124(.a(s_82), .O(gate22inter3));
  inv1  gate1125(.a(s_83), .O(gate22inter4));
  nand2 gate1126(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1127(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1128(.a(G27), .O(gate22inter7));
  inv1  gate1129(.a(G28), .O(gate22inter8));
  nand2 gate1130(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1131(.a(s_83), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1132(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1133(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1134(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2199(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2200(.a(gate24inter0), .b(s_236), .O(gate24inter1));
  and2  gate2201(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2202(.a(s_236), .O(gate24inter3));
  inv1  gate2203(.a(s_237), .O(gate24inter4));
  nand2 gate2204(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2205(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2206(.a(G31), .O(gate24inter7));
  inv1  gate2207(.a(G32), .O(gate24inter8));
  nand2 gate2208(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2209(.a(s_237), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2210(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2211(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2212(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1023(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1024(.a(gate27inter0), .b(s_68), .O(gate27inter1));
  and2  gate1025(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1026(.a(s_68), .O(gate27inter3));
  inv1  gate1027(.a(s_69), .O(gate27inter4));
  nand2 gate1028(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1029(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1030(.a(G2), .O(gate27inter7));
  inv1  gate1031(.a(G6), .O(gate27inter8));
  nand2 gate1032(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1033(.a(s_69), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1034(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1035(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1036(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1709(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1710(.a(gate30inter0), .b(s_166), .O(gate30inter1));
  and2  gate1711(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1712(.a(s_166), .O(gate30inter3));
  inv1  gate1713(.a(s_167), .O(gate30inter4));
  nand2 gate1714(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1715(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1716(.a(G11), .O(gate30inter7));
  inv1  gate1717(.a(G15), .O(gate30inter8));
  nand2 gate1718(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1719(.a(s_167), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1720(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1721(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1722(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1737(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1738(.a(gate32inter0), .b(s_170), .O(gate32inter1));
  and2  gate1739(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1740(.a(s_170), .O(gate32inter3));
  inv1  gate1741(.a(s_171), .O(gate32inter4));
  nand2 gate1742(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1743(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1744(.a(G12), .O(gate32inter7));
  inv1  gate1745(.a(G16), .O(gate32inter8));
  nand2 gate1746(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1747(.a(s_171), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1748(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1749(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1750(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate869(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate870(.a(gate33inter0), .b(s_46), .O(gate33inter1));
  and2  gate871(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate872(.a(s_46), .O(gate33inter3));
  inv1  gate873(.a(s_47), .O(gate33inter4));
  nand2 gate874(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate875(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate876(.a(G17), .O(gate33inter7));
  inv1  gate877(.a(G21), .O(gate33inter8));
  nand2 gate878(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate879(.a(s_47), .b(gate33inter3), .O(gate33inter10));
  nor2  gate880(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate881(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate882(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1443(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1444(.a(gate40inter0), .b(s_128), .O(gate40inter1));
  and2  gate1445(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1446(.a(s_128), .O(gate40inter3));
  inv1  gate1447(.a(s_129), .O(gate40inter4));
  nand2 gate1448(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1449(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1450(.a(G28), .O(gate40inter7));
  inv1  gate1451(.a(G32), .O(gate40inter8));
  nand2 gate1452(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1453(.a(s_129), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1454(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1455(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1456(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1135(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1136(.a(gate44inter0), .b(s_84), .O(gate44inter1));
  and2  gate1137(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1138(.a(s_84), .O(gate44inter3));
  inv1  gate1139(.a(s_85), .O(gate44inter4));
  nand2 gate1140(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1141(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1142(.a(G4), .O(gate44inter7));
  inv1  gate1143(.a(G269), .O(gate44inter8));
  nand2 gate1144(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1145(.a(s_85), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1146(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1147(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1148(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1331(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1332(.a(gate47inter0), .b(s_112), .O(gate47inter1));
  and2  gate1333(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1334(.a(s_112), .O(gate47inter3));
  inv1  gate1335(.a(s_113), .O(gate47inter4));
  nand2 gate1336(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1337(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1338(.a(G7), .O(gate47inter7));
  inv1  gate1339(.a(G275), .O(gate47inter8));
  nand2 gate1340(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1341(.a(s_113), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1342(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1343(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1344(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1303(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1304(.a(gate48inter0), .b(s_108), .O(gate48inter1));
  and2  gate1305(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1306(.a(s_108), .O(gate48inter3));
  inv1  gate1307(.a(s_109), .O(gate48inter4));
  nand2 gate1308(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1309(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1310(.a(G8), .O(gate48inter7));
  inv1  gate1311(.a(G275), .O(gate48inter8));
  nand2 gate1312(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1313(.a(s_109), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1314(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1315(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1316(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2423(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2424(.a(gate50inter0), .b(s_268), .O(gate50inter1));
  and2  gate2425(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2426(.a(s_268), .O(gate50inter3));
  inv1  gate2427(.a(s_269), .O(gate50inter4));
  nand2 gate2428(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2429(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2430(.a(G10), .O(gate50inter7));
  inv1  gate2431(.a(G278), .O(gate50inter8));
  nand2 gate2432(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2433(.a(s_269), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2434(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2435(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2436(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate757(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate758(.a(gate52inter0), .b(s_30), .O(gate52inter1));
  and2  gate759(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate760(.a(s_30), .O(gate52inter3));
  inv1  gate761(.a(s_31), .O(gate52inter4));
  nand2 gate762(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate763(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate764(.a(G12), .O(gate52inter7));
  inv1  gate765(.a(G281), .O(gate52inter8));
  nand2 gate766(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate767(.a(s_31), .b(gate52inter3), .O(gate52inter10));
  nor2  gate768(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate769(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate770(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate547(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate548(.a(gate56inter0), .b(s_0), .O(gate56inter1));
  and2  gate549(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate550(.a(s_0), .O(gate56inter3));
  inv1  gate551(.a(s_1), .O(gate56inter4));
  nand2 gate552(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate553(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate554(.a(G16), .O(gate56inter7));
  inv1  gate555(.a(G287), .O(gate56inter8));
  nand2 gate556(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate557(.a(s_1), .b(gate56inter3), .O(gate56inter10));
  nor2  gate558(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate559(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate560(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate2045(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2046(.a(gate63inter0), .b(s_214), .O(gate63inter1));
  and2  gate2047(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2048(.a(s_214), .O(gate63inter3));
  inv1  gate2049(.a(s_215), .O(gate63inter4));
  nand2 gate2050(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2051(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2052(.a(G23), .O(gate63inter7));
  inv1  gate2053(.a(G299), .O(gate63inter8));
  nand2 gate2054(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2055(.a(s_215), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2056(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2057(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2058(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2255(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2256(.a(gate64inter0), .b(s_244), .O(gate64inter1));
  and2  gate2257(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2258(.a(s_244), .O(gate64inter3));
  inv1  gate2259(.a(s_245), .O(gate64inter4));
  nand2 gate2260(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2261(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2262(.a(G24), .O(gate64inter7));
  inv1  gate2263(.a(G299), .O(gate64inter8));
  nand2 gate2264(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2265(.a(s_245), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2266(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2267(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2268(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1499(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1500(.a(gate66inter0), .b(s_136), .O(gate66inter1));
  and2  gate1501(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1502(.a(s_136), .O(gate66inter3));
  inv1  gate1503(.a(s_137), .O(gate66inter4));
  nand2 gate1504(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1505(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1506(.a(G26), .O(gate66inter7));
  inv1  gate1507(.a(G302), .O(gate66inter8));
  nand2 gate1508(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1509(.a(s_137), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1510(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1511(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1512(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1205(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1206(.a(gate70inter0), .b(s_94), .O(gate70inter1));
  and2  gate1207(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1208(.a(s_94), .O(gate70inter3));
  inv1  gate1209(.a(s_95), .O(gate70inter4));
  nand2 gate1210(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1211(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1212(.a(G30), .O(gate70inter7));
  inv1  gate1213(.a(G308), .O(gate70inter8));
  nand2 gate1214(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1215(.a(s_95), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1216(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1217(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1218(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2003(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2004(.a(gate74inter0), .b(s_208), .O(gate74inter1));
  and2  gate2005(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2006(.a(s_208), .O(gate74inter3));
  inv1  gate2007(.a(s_209), .O(gate74inter4));
  nand2 gate2008(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2009(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2010(.a(G5), .O(gate74inter7));
  inv1  gate2011(.a(G314), .O(gate74inter8));
  nand2 gate2012(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2013(.a(s_209), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2014(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2015(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2016(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1177(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1178(.a(gate75inter0), .b(s_90), .O(gate75inter1));
  and2  gate1179(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1180(.a(s_90), .O(gate75inter3));
  inv1  gate1181(.a(s_91), .O(gate75inter4));
  nand2 gate1182(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1183(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1184(.a(G9), .O(gate75inter7));
  inv1  gate1185(.a(G317), .O(gate75inter8));
  nand2 gate1186(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1187(.a(s_91), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1188(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1189(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1190(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1975(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1976(.a(gate81inter0), .b(s_204), .O(gate81inter1));
  and2  gate1977(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1978(.a(s_204), .O(gate81inter3));
  inv1  gate1979(.a(s_205), .O(gate81inter4));
  nand2 gate1980(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1981(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1982(.a(G3), .O(gate81inter7));
  inv1  gate1983(.a(G326), .O(gate81inter8));
  nand2 gate1984(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1985(.a(s_205), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1986(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1987(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1988(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate953(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate954(.a(gate82inter0), .b(s_58), .O(gate82inter1));
  and2  gate955(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate956(.a(s_58), .O(gate82inter3));
  inv1  gate957(.a(s_59), .O(gate82inter4));
  nand2 gate958(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate959(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate960(.a(G7), .O(gate82inter7));
  inv1  gate961(.a(G326), .O(gate82inter8));
  nand2 gate962(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate963(.a(s_59), .b(gate82inter3), .O(gate82inter10));
  nor2  gate964(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate965(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate966(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1541(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1542(.a(gate83inter0), .b(s_142), .O(gate83inter1));
  and2  gate1543(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1544(.a(s_142), .O(gate83inter3));
  inv1  gate1545(.a(s_143), .O(gate83inter4));
  nand2 gate1546(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1547(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1548(.a(G11), .O(gate83inter7));
  inv1  gate1549(.a(G329), .O(gate83inter8));
  nand2 gate1550(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1551(.a(s_143), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1552(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1553(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1554(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1583(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1584(.a(gate92inter0), .b(s_148), .O(gate92inter1));
  and2  gate1585(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1586(.a(s_148), .O(gate92inter3));
  inv1  gate1587(.a(s_149), .O(gate92inter4));
  nand2 gate1588(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1589(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1590(.a(G29), .O(gate92inter7));
  inv1  gate1591(.a(G341), .O(gate92inter8));
  nand2 gate1592(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1593(.a(s_149), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1594(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1595(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1596(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1863(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1864(.a(gate93inter0), .b(s_188), .O(gate93inter1));
  and2  gate1865(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1866(.a(s_188), .O(gate93inter3));
  inv1  gate1867(.a(s_189), .O(gate93inter4));
  nand2 gate1868(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1869(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1870(.a(G18), .O(gate93inter7));
  inv1  gate1871(.a(G344), .O(gate93inter8));
  nand2 gate1872(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1873(.a(s_189), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1874(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1875(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1876(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate715(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate716(.a(gate95inter0), .b(s_24), .O(gate95inter1));
  and2  gate717(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate718(.a(s_24), .O(gate95inter3));
  inv1  gate719(.a(s_25), .O(gate95inter4));
  nand2 gate720(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate721(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate722(.a(G26), .O(gate95inter7));
  inv1  gate723(.a(G347), .O(gate95inter8));
  nand2 gate724(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate725(.a(s_25), .b(gate95inter3), .O(gate95inter10));
  nor2  gate726(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate727(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate728(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate659(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate660(.a(gate96inter0), .b(s_16), .O(gate96inter1));
  and2  gate661(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate662(.a(s_16), .O(gate96inter3));
  inv1  gate663(.a(s_17), .O(gate96inter4));
  nand2 gate664(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate665(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate666(.a(G30), .O(gate96inter7));
  inv1  gate667(.a(G347), .O(gate96inter8));
  nand2 gate668(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate669(.a(s_17), .b(gate96inter3), .O(gate96inter10));
  nor2  gate670(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate671(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate672(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1345(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1346(.a(gate99inter0), .b(s_114), .O(gate99inter1));
  and2  gate1347(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1348(.a(s_114), .O(gate99inter3));
  inv1  gate1349(.a(s_115), .O(gate99inter4));
  nand2 gate1350(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1351(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1352(.a(G27), .O(gate99inter7));
  inv1  gate1353(.a(G353), .O(gate99inter8));
  nand2 gate1354(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1355(.a(s_115), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1356(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1357(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1358(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1625(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1626(.a(gate102inter0), .b(s_154), .O(gate102inter1));
  and2  gate1627(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1628(.a(s_154), .O(gate102inter3));
  inv1  gate1629(.a(s_155), .O(gate102inter4));
  nand2 gate1630(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1631(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1632(.a(G24), .O(gate102inter7));
  inv1  gate1633(.a(G356), .O(gate102inter8));
  nand2 gate1634(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1635(.a(s_155), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1636(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1637(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1638(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1051(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1052(.a(gate103inter0), .b(s_72), .O(gate103inter1));
  and2  gate1053(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1054(.a(s_72), .O(gate103inter3));
  inv1  gate1055(.a(s_73), .O(gate103inter4));
  nand2 gate1056(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1057(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1058(.a(G28), .O(gate103inter7));
  inv1  gate1059(.a(G359), .O(gate103inter8));
  nand2 gate1060(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1061(.a(s_73), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1062(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1063(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1064(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2129(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2130(.a(gate105inter0), .b(s_226), .O(gate105inter1));
  and2  gate2131(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2132(.a(s_226), .O(gate105inter3));
  inv1  gate2133(.a(s_227), .O(gate105inter4));
  nand2 gate2134(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2135(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2136(.a(G362), .O(gate105inter7));
  inv1  gate2137(.a(G363), .O(gate105inter8));
  nand2 gate2138(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2139(.a(s_227), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2140(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2141(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2142(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1793(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1794(.a(gate108inter0), .b(s_178), .O(gate108inter1));
  and2  gate1795(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1796(.a(s_178), .O(gate108inter3));
  inv1  gate1797(.a(s_179), .O(gate108inter4));
  nand2 gate1798(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1799(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1800(.a(G368), .O(gate108inter7));
  inv1  gate1801(.a(G369), .O(gate108inter8));
  nand2 gate1802(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1803(.a(s_179), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1804(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1805(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1806(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate967(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate968(.a(gate109inter0), .b(s_60), .O(gate109inter1));
  and2  gate969(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate970(.a(s_60), .O(gate109inter3));
  inv1  gate971(.a(s_61), .O(gate109inter4));
  nand2 gate972(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate973(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate974(.a(G370), .O(gate109inter7));
  inv1  gate975(.a(G371), .O(gate109inter8));
  nand2 gate976(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate977(.a(s_61), .b(gate109inter3), .O(gate109inter10));
  nor2  gate978(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate979(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate980(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1485(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1486(.a(gate110inter0), .b(s_134), .O(gate110inter1));
  and2  gate1487(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1488(.a(s_134), .O(gate110inter3));
  inv1  gate1489(.a(s_135), .O(gate110inter4));
  nand2 gate1490(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1491(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1492(.a(G372), .O(gate110inter7));
  inv1  gate1493(.a(G373), .O(gate110inter8));
  nand2 gate1494(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1495(.a(s_135), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1496(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1497(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1498(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1149(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1150(.a(gate111inter0), .b(s_86), .O(gate111inter1));
  and2  gate1151(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1152(.a(s_86), .O(gate111inter3));
  inv1  gate1153(.a(s_87), .O(gate111inter4));
  nand2 gate1154(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1155(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1156(.a(G374), .O(gate111inter7));
  inv1  gate1157(.a(G375), .O(gate111inter8));
  nand2 gate1158(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1159(.a(s_87), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1160(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1161(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1162(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate673(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate674(.a(gate112inter0), .b(s_18), .O(gate112inter1));
  and2  gate675(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate676(.a(s_18), .O(gate112inter3));
  inv1  gate677(.a(s_19), .O(gate112inter4));
  nand2 gate678(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate679(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate680(.a(G376), .O(gate112inter7));
  inv1  gate681(.a(G377), .O(gate112inter8));
  nand2 gate682(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate683(.a(s_19), .b(gate112inter3), .O(gate112inter10));
  nor2  gate684(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate685(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate686(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1611(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1612(.a(gate113inter0), .b(s_152), .O(gate113inter1));
  and2  gate1613(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1614(.a(s_152), .O(gate113inter3));
  inv1  gate1615(.a(s_153), .O(gate113inter4));
  nand2 gate1616(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1617(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1618(.a(G378), .O(gate113inter7));
  inv1  gate1619(.a(G379), .O(gate113inter8));
  nand2 gate1620(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1621(.a(s_153), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1622(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1623(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1624(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2409(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2410(.a(gate118inter0), .b(s_266), .O(gate118inter1));
  and2  gate2411(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2412(.a(s_266), .O(gate118inter3));
  inv1  gate2413(.a(s_267), .O(gate118inter4));
  nand2 gate2414(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2415(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2416(.a(G388), .O(gate118inter7));
  inv1  gate2417(.a(G389), .O(gate118inter8));
  nand2 gate2418(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2419(.a(s_267), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2420(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2421(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2422(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2325(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2326(.a(gate126inter0), .b(s_254), .O(gate126inter1));
  and2  gate2327(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2328(.a(s_254), .O(gate126inter3));
  inv1  gate2329(.a(s_255), .O(gate126inter4));
  nand2 gate2330(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2331(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2332(.a(G404), .O(gate126inter7));
  inv1  gate2333(.a(G405), .O(gate126inter8));
  nand2 gate2334(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2335(.a(s_255), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2336(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2337(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2338(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1765(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1766(.a(gate127inter0), .b(s_174), .O(gate127inter1));
  and2  gate1767(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1768(.a(s_174), .O(gate127inter3));
  inv1  gate1769(.a(s_175), .O(gate127inter4));
  nand2 gate1770(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1771(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1772(.a(G406), .O(gate127inter7));
  inv1  gate1773(.a(G407), .O(gate127inter8));
  nand2 gate1774(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1775(.a(s_175), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1776(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1777(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1778(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate603(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate604(.a(gate132inter0), .b(s_8), .O(gate132inter1));
  and2  gate605(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate606(.a(s_8), .O(gate132inter3));
  inv1  gate607(.a(s_9), .O(gate132inter4));
  nand2 gate608(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate609(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate610(.a(G416), .O(gate132inter7));
  inv1  gate611(.a(G417), .O(gate132inter8));
  nand2 gate612(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate613(.a(s_9), .b(gate132inter3), .O(gate132inter10));
  nor2  gate614(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate615(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate616(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate589(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate590(.a(gate135inter0), .b(s_6), .O(gate135inter1));
  and2  gate591(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate592(.a(s_6), .O(gate135inter3));
  inv1  gate593(.a(s_7), .O(gate135inter4));
  nand2 gate594(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate595(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate596(.a(G422), .O(gate135inter7));
  inv1  gate597(.a(G423), .O(gate135inter8));
  nand2 gate598(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate599(.a(s_7), .b(gate135inter3), .O(gate135inter10));
  nor2  gate600(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate601(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate602(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate2437(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2438(.a(gate136inter0), .b(s_270), .O(gate136inter1));
  and2  gate2439(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2440(.a(s_270), .O(gate136inter3));
  inv1  gate2441(.a(s_271), .O(gate136inter4));
  nand2 gate2442(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2443(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2444(.a(G424), .O(gate136inter7));
  inv1  gate2445(.a(G425), .O(gate136inter8));
  nand2 gate2446(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2447(.a(s_271), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2448(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2449(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2450(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1905(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1906(.a(gate142inter0), .b(s_194), .O(gate142inter1));
  and2  gate1907(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1908(.a(s_194), .O(gate142inter3));
  inv1  gate1909(.a(s_195), .O(gate142inter4));
  nand2 gate1910(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1911(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1912(.a(G456), .O(gate142inter7));
  inv1  gate1913(.a(G459), .O(gate142inter8));
  nand2 gate1914(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1915(.a(s_195), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1916(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1917(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1918(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2059(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2060(.a(gate144inter0), .b(s_216), .O(gate144inter1));
  and2  gate2061(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2062(.a(s_216), .O(gate144inter3));
  inv1  gate2063(.a(s_217), .O(gate144inter4));
  nand2 gate2064(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2065(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2066(.a(G468), .O(gate144inter7));
  inv1  gate2067(.a(G471), .O(gate144inter8));
  nand2 gate2068(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2069(.a(s_217), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2070(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2071(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2072(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2395(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2396(.a(gate147inter0), .b(s_264), .O(gate147inter1));
  and2  gate2397(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2398(.a(s_264), .O(gate147inter3));
  inv1  gate2399(.a(s_265), .O(gate147inter4));
  nand2 gate2400(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2401(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2402(.a(G486), .O(gate147inter7));
  inv1  gate2403(.a(G489), .O(gate147inter8));
  nand2 gate2404(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2405(.a(s_265), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2406(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2407(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2408(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate2283(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2284(.a(gate148inter0), .b(s_248), .O(gate148inter1));
  and2  gate2285(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2286(.a(s_248), .O(gate148inter3));
  inv1  gate2287(.a(s_249), .O(gate148inter4));
  nand2 gate2288(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2289(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2290(.a(G492), .O(gate148inter7));
  inv1  gate2291(.a(G495), .O(gate148inter8));
  nand2 gate2292(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2293(.a(s_249), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2294(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2295(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2296(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1653(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1654(.a(gate155inter0), .b(s_158), .O(gate155inter1));
  and2  gate1655(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1656(.a(s_158), .O(gate155inter3));
  inv1  gate1657(.a(s_159), .O(gate155inter4));
  nand2 gate1658(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1659(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1660(.a(G432), .O(gate155inter7));
  inv1  gate1661(.a(G525), .O(gate155inter8));
  nand2 gate1662(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1663(.a(s_159), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1664(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1665(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1666(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1989(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1990(.a(gate158inter0), .b(s_206), .O(gate158inter1));
  and2  gate1991(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1992(.a(s_206), .O(gate158inter3));
  inv1  gate1993(.a(s_207), .O(gate158inter4));
  nand2 gate1994(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1995(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1996(.a(G441), .O(gate158inter7));
  inv1  gate1997(.a(G528), .O(gate158inter8));
  nand2 gate1998(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1999(.a(s_207), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2000(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2001(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2002(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1821(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1822(.a(gate159inter0), .b(s_182), .O(gate159inter1));
  and2  gate1823(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1824(.a(s_182), .O(gate159inter3));
  inv1  gate1825(.a(s_183), .O(gate159inter4));
  nand2 gate1826(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1827(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1828(.a(G444), .O(gate159inter7));
  inv1  gate1829(.a(G531), .O(gate159inter8));
  nand2 gate1830(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1831(.a(s_183), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1832(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1833(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1834(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate883(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate884(.a(gate163inter0), .b(s_48), .O(gate163inter1));
  and2  gate885(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate886(.a(s_48), .O(gate163inter3));
  inv1  gate887(.a(s_49), .O(gate163inter4));
  nand2 gate888(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate889(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate890(.a(G456), .O(gate163inter7));
  inv1  gate891(.a(G537), .O(gate163inter8));
  nand2 gate892(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate893(.a(s_49), .b(gate163inter3), .O(gate163inter10));
  nor2  gate894(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate895(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate896(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2213(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2214(.a(gate168inter0), .b(s_238), .O(gate168inter1));
  and2  gate2215(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2216(.a(s_238), .O(gate168inter3));
  inv1  gate2217(.a(s_239), .O(gate168inter4));
  nand2 gate2218(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2219(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2220(.a(G471), .O(gate168inter7));
  inv1  gate2221(.a(G543), .O(gate168inter8));
  nand2 gate2222(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2223(.a(s_239), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2224(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2225(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2226(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1513(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1514(.a(gate170inter0), .b(s_138), .O(gate170inter1));
  and2  gate1515(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1516(.a(s_138), .O(gate170inter3));
  inv1  gate1517(.a(s_139), .O(gate170inter4));
  nand2 gate1518(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1519(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1520(.a(G477), .O(gate170inter7));
  inv1  gate1521(.a(G546), .O(gate170inter8));
  nand2 gate1522(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1523(.a(s_139), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1524(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1525(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1526(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1429(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1430(.a(gate172inter0), .b(s_126), .O(gate172inter1));
  and2  gate1431(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1432(.a(s_126), .O(gate172inter3));
  inv1  gate1433(.a(s_127), .O(gate172inter4));
  nand2 gate1434(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1435(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1436(.a(G483), .O(gate172inter7));
  inv1  gate1437(.a(G549), .O(gate172inter8));
  nand2 gate1438(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1439(.a(s_127), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1440(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1441(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1442(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1681(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1682(.a(gate176inter0), .b(s_162), .O(gate176inter1));
  and2  gate1683(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1684(.a(s_162), .O(gate176inter3));
  inv1  gate1685(.a(s_163), .O(gate176inter4));
  nand2 gate1686(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1687(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1688(.a(G495), .O(gate176inter7));
  inv1  gate1689(.a(G555), .O(gate176inter8));
  nand2 gate1690(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1691(.a(s_163), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1692(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1693(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1694(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate2311(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2312(.a(gate177inter0), .b(s_252), .O(gate177inter1));
  and2  gate2313(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2314(.a(s_252), .O(gate177inter3));
  inv1  gate2315(.a(s_253), .O(gate177inter4));
  nand2 gate2316(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2317(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2318(.a(G498), .O(gate177inter7));
  inv1  gate2319(.a(G558), .O(gate177inter8));
  nand2 gate2320(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2321(.a(s_253), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2322(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2323(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2324(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1219(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1220(.a(gate180inter0), .b(s_96), .O(gate180inter1));
  and2  gate1221(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1222(.a(s_96), .O(gate180inter3));
  inv1  gate1223(.a(s_97), .O(gate180inter4));
  nand2 gate1224(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1225(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1226(.a(G507), .O(gate180inter7));
  inv1  gate1227(.a(G561), .O(gate180inter8));
  nand2 gate1228(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1229(.a(s_97), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1230(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1231(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1232(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1275(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1276(.a(gate184inter0), .b(s_104), .O(gate184inter1));
  and2  gate1277(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1278(.a(s_104), .O(gate184inter3));
  inv1  gate1279(.a(s_105), .O(gate184inter4));
  nand2 gate1280(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1281(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1282(.a(G519), .O(gate184inter7));
  inv1  gate1283(.a(G567), .O(gate184inter8));
  nand2 gate1284(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1285(.a(s_105), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1286(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1287(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1288(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate925(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate926(.a(gate185inter0), .b(s_54), .O(gate185inter1));
  and2  gate927(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate928(.a(s_54), .O(gate185inter3));
  inv1  gate929(.a(s_55), .O(gate185inter4));
  nand2 gate930(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate931(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate932(.a(G570), .O(gate185inter7));
  inv1  gate933(.a(G571), .O(gate185inter8));
  nand2 gate934(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate935(.a(s_55), .b(gate185inter3), .O(gate185inter10));
  nor2  gate936(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate937(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate938(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1835(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1836(.a(gate189inter0), .b(s_184), .O(gate189inter1));
  and2  gate1837(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1838(.a(s_184), .O(gate189inter3));
  inv1  gate1839(.a(s_185), .O(gate189inter4));
  nand2 gate1840(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1841(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1842(.a(G578), .O(gate189inter7));
  inv1  gate1843(.a(G579), .O(gate189inter8));
  nand2 gate1844(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1845(.a(s_185), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1846(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1847(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1848(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate687(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate688(.a(gate190inter0), .b(s_20), .O(gate190inter1));
  and2  gate689(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate690(.a(s_20), .O(gate190inter3));
  inv1  gate691(.a(s_21), .O(gate190inter4));
  nand2 gate692(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate693(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate694(.a(G580), .O(gate190inter7));
  inv1  gate695(.a(G581), .O(gate190inter8));
  nand2 gate696(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate697(.a(s_21), .b(gate190inter3), .O(gate190inter10));
  nor2  gate698(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate699(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate700(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1261(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1262(.a(gate195inter0), .b(s_102), .O(gate195inter1));
  and2  gate1263(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1264(.a(s_102), .O(gate195inter3));
  inv1  gate1265(.a(s_103), .O(gate195inter4));
  nand2 gate1266(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1267(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1268(.a(G590), .O(gate195inter7));
  inv1  gate1269(.a(G591), .O(gate195inter8));
  nand2 gate1270(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1271(.a(s_103), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1272(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1273(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1274(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2087(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2088(.a(gate196inter0), .b(s_220), .O(gate196inter1));
  and2  gate2089(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2090(.a(s_220), .O(gate196inter3));
  inv1  gate2091(.a(s_221), .O(gate196inter4));
  nand2 gate2092(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2093(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2094(.a(G592), .O(gate196inter7));
  inv1  gate2095(.a(G593), .O(gate196inter8));
  nand2 gate2096(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2097(.a(s_221), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2098(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2099(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2100(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate617(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate618(.a(gate207inter0), .b(s_10), .O(gate207inter1));
  and2  gate619(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate620(.a(s_10), .O(gate207inter3));
  inv1  gate621(.a(s_11), .O(gate207inter4));
  nand2 gate622(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate623(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate624(.a(G622), .O(gate207inter7));
  inv1  gate625(.a(G632), .O(gate207inter8));
  nand2 gate626(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate627(.a(s_11), .b(gate207inter3), .O(gate207inter10));
  nor2  gate628(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate629(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate630(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1667(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1668(.a(gate209inter0), .b(s_160), .O(gate209inter1));
  and2  gate1669(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1670(.a(s_160), .O(gate209inter3));
  inv1  gate1671(.a(s_161), .O(gate209inter4));
  nand2 gate1672(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1673(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1674(.a(G602), .O(gate209inter7));
  inv1  gate1675(.a(G666), .O(gate209inter8));
  nand2 gate1676(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1677(.a(s_161), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1678(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1679(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1680(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2269(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2270(.a(gate210inter0), .b(s_246), .O(gate210inter1));
  and2  gate2271(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2272(.a(s_246), .O(gate210inter3));
  inv1  gate2273(.a(s_247), .O(gate210inter4));
  nand2 gate2274(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2275(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2276(.a(G607), .O(gate210inter7));
  inv1  gate2277(.a(G666), .O(gate210inter8));
  nand2 gate2278(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2279(.a(s_247), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2280(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2281(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2282(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1779(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1780(.a(gate212inter0), .b(s_176), .O(gate212inter1));
  and2  gate1781(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1782(.a(s_176), .O(gate212inter3));
  inv1  gate1783(.a(s_177), .O(gate212inter4));
  nand2 gate1784(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1785(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1786(.a(G617), .O(gate212inter7));
  inv1  gate1787(.a(G669), .O(gate212inter8));
  nand2 gate1788(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1789(.a(s_177), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1790(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1791(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1792(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2017(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2018(.a(gate217inter0), .b(s_210), .O(gate217inter1));
  and2  gate2019(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2020(.a(s_210), .O(gate217inter3));
  inv1  gate2021(.a(s_211), .O(gate217inter4));
  nand2 gate2022(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2023(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2024(.a(G622), .O(gate217inter7));
  inv1  gate2025(.a(G678), .O(gate217inter8));
  nand2 gate2026(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2027(.a(s_211), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2028(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2029(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2030(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1401(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1402(.a(gate226inter0), .b(s_122), .O(gate226inter1));
  and2  gate1403(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1404(.a(s_122), .O(gate226inter3));
  inv1  gate1405(.a(s_123), .O(gate226inter4));
  nand2 gate1406(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1407(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1408(.a(G692), .O(gate226inter7));
  inv1  gate1409(.a(G693), .O(gate226inter8));
  nand2 gate1410(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1411(.a(s_123), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1412(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1413(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1414(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate785(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate786(.a(gate228inter0), .b(s_34), .O(gate228inter1));
  and2  gate787(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate788(.a(s_34), .O(gate228inter3));
  inv1  gate789(.a(s_35), .O(gate228inter4));
  nand2 gate790(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate791(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate792(.a(G696), .O(gate228inter7));
  inv1  gate793(.a(G697), .O(gate228inter8));
  nand2 gate794(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate795(.a(s_35), .b(gate228inter3), .O(gate228inter10));
  nor2  gate796(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate797(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate798(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate813(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate814(.a(gate231inter0), .b(s_38), .O(gate231inter1));
  and2  gate815(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate816(.a(s_38), .O(gate231inter3));
  inv1  gate817(.a(s_39), .O(gate231inter4));
  nand2 gate818(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate819(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate820(.a(G702), .O(gate231inter7));
  inv1  gate821(.a(G703), .O(gate231inter8));
  nand2 gate822(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate823(.a(s_39), .b(gate231inter3), .O(gate231inter10));
  nor2  gate824(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate825(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate826(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate995(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate996(.a(gate234inter0), .b(s_64), .O(gate234inter1));
  and2  gate997(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate998(.a(s_64), .O(gate234inter3));
  inv1  gate999(.a(s_65), .O(gate234inter4));
  nand2 gate1000(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1001(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1002(.a(G245), .O(gate234inter7));
  inv1  gate1003(.a(G721), .O(gate234inter8));
  nand2 gate1004(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1005(.a(s_65), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1006(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1007(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1008(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1359(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1360(.a(gate237inter0), .b(s_116), .O(gate237inter1));
  and2  gate1361(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1362(.a(s_116), .O(gate237inter3));
  inv1  gate1363(.a(s_117), .O(gate237inter4));
  nand2 gate1364(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1365(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1366(.a(G254), .O(gate237inter7));
  inv1  gate1367(.a(G706), .O(gate237inter8));
  nand2 gate1368(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1369(.a(s_117), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1370(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1371(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1372(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1079(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1080(.a(gate238inter0), .b(s_76), .O(gate238inter1));
  and2  gate1081(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1082(.a(s_76), .O(gate238inter3));
  inv1  gate1083(.a(s_77), .O(gate238inter4));
  nand2 gate1084(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1085(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1086(.a(G257), .O(gate238inter7));
  inv1  gate1087(.a(G709), .O(gate238inter8));
  nand2 gate1088(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1089(.a(s_77), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1090(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1091(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1092(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1415(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1416(.a(gate243inter0), .b(s_124), .O(gate243inter1));
  and2  gate1417(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1418(.a(s_124), .O(gate243inter3));
  inv1  gate1419(.a(s_125), .O(gate243inter4));
  nand2 gate1420(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1421(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1422(.a(G245), .O(gate243inter7));
  inv1  gate1423(.a(G733), .O(gate243inter8));
  nand2 gate1424(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1425(.a(s_125), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1426(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1427(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1428(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1877(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1878(.a(gate244inter0), .b(s_190), .O(gate244inter1));
  and2  gate1879(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1880(.a(s_190), .O(gate244inter3));
  inv1  gate1881(.a(s_191), .O(gate244inter4));
  nand2 gate1882(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1883(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1884(.a(G721), .O(gate244inter7));
  inv1  gate1885(.a(G733), .O(gate244inter8));
  nand2 gate1886(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1887(.a(s_191), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1888(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1889(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1890(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate729(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate730(.a(gate247inter0), .b(s_26), .O(gate247inter1));
  and2  gate731(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate732(.a(s_26), .O(gate247inter3));
  inv1  gate733(.a(s_27), .O(gate247inter4));
  nand2 gate734(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate735(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate736(.a(G251), .O(gate247inter7));
  inv1  gate737(.a(G739), .O(gate247inter8));
  nand2 gate738(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate739(.a(s_27), .b(gate247inter3), .O(gate247inter10));
  nor2  gate740(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate741(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate742(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate827(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate828(.a(gate248inter0), .b(s_40), .O(gate248inter1));
  and2  gate829(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate830(.a(s_40), .O(gate248inter3));
  inv1  gate831(.a(s_41), .O(gate248inter4));
  nand2 gate832(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate833(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate834(.a(G727), .O(gate248inter7));
  inv1  gate835(.a(G739), .O(gate248inter8));
  nand2 gate836(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate837(.a(s_41), .b(gate248inter3), .O(gate248inter10));
  nor2  gate838(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate839(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate840(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1849(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1850(.a(gate250inter0), .b(s_186), .O(gate250inter1));
  and2  gate1851(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1852(.a(s_186), .O(gate250inter3));
  inv1  gate1853(.a(s_187), .O(gate250inter4));
  nand2 gate1854(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1855(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1856(.a(G706), .O(gate250inter7));
  inv1  gate1857(.a(G742), .O(gate250inter8));
  nand2 gate1858(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1859(.a(s_187), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1860(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1861(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1862(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1317(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1318(.a(gate253inter0), .b(s_110), .O(gate253inter1));
  and2  gate1319(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1320(.a(s_110), .O(gate253inter3));
  inv1  gate1321(.a(s_111), .O(gate253inter4));
  nand2 gate1322(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1323(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1324(.a(G260), .O(gate253inter7));
  inv1  gate1325(.a(G748), .O(gate253inter8));
  nand2 gate1326(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1327(.a(s_111), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1328(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1329(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1330(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate855(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate856(.a(gate258inter0), .b(s_44), .O(gate258inter1));
  and2  gate857(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate858(.a(s_44), .O(gate258inter3));
  inv1  gate859(.a(s_45), .O(gate258inter4));
  nand2 gate860(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate861(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate862(.a(G756), .O(gate258inter7));
  inv1  gate863(.a(G757), .O(gate258inter8));
  nand2 gate864(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate865(.a(s_45), .b(gate258inter3), .O(gate258inter10));
  nor2  gate866(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate867(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate868(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate2171(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2172(.a(gate259inter0), .b(s_232), .O(gate259inter1));
  and2  gate2173(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2174(.a(s_232), .O(gate259inter3));
  inv1  gate2175(.a(s_233), .O(gate259inter4));
  nand2 gate2176(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2177(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2178(.a(G758), .O(gate259inter7));
  inv1  gate2179(.a(G759), .O(gate259inter8));
  nand2 gate2180(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2181(.a(s_233), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2182(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2183(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2184(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2157(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2158(.a(gate267inter0), .b(s_230), .O(gate267inter1));
  and2  gate2159(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2160(.a(s_230), .O(gate267inter3));
  inv1  gate2161(.a(s_231), .O(gate267inter4));
  nand2 gate2162(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2163(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2164(.a(G648), .O(gate267inter7));
  inv1  gate2165(.a(G776), .O(gate267inter8));
  nand2 gate2166(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2167(.a(s_231), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2168(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2169(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2170(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2367(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2368(.a(gate270inter0), .b(s_260), .O(gate270inter1));
  and2  gate2369(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2370(.a(s_260), .O(gate270inter3));
  inv1  gate2371(.a(s_261), .O(gate270inter4));
  nand2 gate2372(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2373(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2374(.a(G657), .O(gate270inter7));
  inv1  gate2375(.a(G785), .O(gate270inter8));
  nand2 gate2376(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2377(.a(s_261), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2378(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2379(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2380(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate575(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate576(.a(gate275inter0), .b(s_4), .O(gate275inter1));
  and2  gate577(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate578(.a(s_4), .O(gate275inter3));
  inv1  gate579(.a(s_5), .O(gate275inter4));
  nand2 gate580(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate581(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate582(.a(G645), .O(gate275inter7));
  inv1  gate583(.a(G797), .O(gate275inter8));
  nand2 gate584(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate585(.a(s_5), .b(gate275inter3), .O(gate275inter10));
  nor2  gate586(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate587(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate588(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate631(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate632(.a(gate277inter0), .b(s_12), .O(gate277inter1));
  and2  gate633(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate634(.a(s_12), .O(gate277inter3));
  inv1  gate635(.a(s_13), .O(gate277inter4));
  nand2 gate636(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate637(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate638(.a(G648), .O(gate277inter7));
  inv1  gate639(.a(G800), .O(gate277inter8));
  nand2 gate640(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate641(.a(s_13), .b(gate277inter3), .O(gate277inter10));
  nor2  gate642(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate643(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate644(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate701(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate702(.a(gate280inter0), .b(s_22), .O(gate280inter1));
  and2  gate703(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate704(.a(s_22), .O(gate280inter3));
  inv1  gate705(.a(s_23), .O(gate280inter4));
  nand2 gate706(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate707(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate708(.a(G779), .O(gate280inter7));
  inv1  gate709(.a(G803), .O(gate280inter8));
  nand2 gate710(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate711(.a(s_23), .b(gate280inter3), .O(gate280inter10));
  nor2  gate712(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate713(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate714(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1891(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1892(.a(gate281inter0), .b(s_192), .O(gate281inter1));
  and2  gate1893(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1894(.a(s_192), .O(gate281inter3));
  inv1  gate1895(.a(s_193), .O(gate281inter4));
  nand2 gate1896(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1897(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1898(.a(G654), .O(gate281inter7));
  inv1  gate1899(.a(G806), .O(gate281inter8));
  nand2 gate1900(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1901(.a(s_193), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1902(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1903(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1904(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2339(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2340(.a(gate282inter0), .b(s_256), .O(gate282inter1));
  and2  gate2341(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2342(.a(s_256), .O(gate282inter3));
  inv1  gate2343(.a(s_257), .O(gate282inter4));
  nand2 gate2344(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2345(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2346(.a(G782), .O(gate282inter7));
  inv1  gate2347(.a(G806), .O(gate282inter8));
  nand2 gate2348(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2349(.a(s_257), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2350(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2351(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2352(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate2353(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2354(.a(gate284inter0), .b(s_258), .O(gate284inter1));
  and2  gate2355(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2356(.a(s_258), .O(gate284inter3));
  inv1  gate2357(.a(s_259), .O(gate284inter4));
  nand2 gate2358(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2359(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2360(.a(G785), .O(gate284inter7));
  inv1  gate2361(.a(G809), .O(gate284inter8));
  nand2 gate2362(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2363(.a(s_259), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2364(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2365(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2366(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1107(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1108(.a(gate285inter0), .b(s_80), .O(gate285inter1));
  and2  gate1109(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1110(.a(s_80), .O(gate285inter3));
  inv1  gate1111(.a(s_81), .O(gate285inter4));
  nand2 gate1112(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1113(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1114(.a(G660), .O(gate285inter7));
  inv1  gate1115(.a(G812), .O(gate285inter8));
  nand2 gate1116(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1117(.a(s_81), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1118(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1119(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1120(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2381(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2382(.a(gate292inter0), .b(s_262), .O(gate292inter1));
  and2  gate2383(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2384(.a(s_262), .O(gate292inter3));
  inv1  gate2385(.a(s_263), .O(gate292inter4));
  nand2 gate2386(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2387(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2388(.a(G824), .O(gate292inter7));
  inv1  gate2389(.a(G825), .O(gate292inter8));
  nand2 gate2390(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2391(.a(s_263), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2392(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2393(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2394(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2115(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2116(.a(gate294inter0), .b(s_224), .O(gate294inter1));
  and2  gate2117(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2118(.a(s_224), .O(gate294inter3));
  inv1  gate2119(.a(s_225), .O(gate294inter4));
  nand2 gate2120(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2121(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2122(.a(G832), .O(gate294inter7));
  inv1  gate2123(.a(G833), .O(gate294inter8));
  nand2 gate2124(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2125(.a(s_225), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2126(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2127(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2128(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate939(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate940(.a(gate387inter0), .b(s_56), .O(gate387inter1));
  and2  gate941(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate942(.a(s_56), .O(gate387inter3));
  inv1  gate943(.a(s_57), .O(gate387inter4));
  nand2 gate944(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate945(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate946(.a(G1), .O(gate387inter7));
  inv1  gate947(.a(G1036), .O(gate387inter8));
  nand2 gate948(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate949(.a(s_57), .b(gate387inter3), .O(gate387inter10));
  nor2  gate950(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate951(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate952(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2185(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2186(.a(gate389inter0), .b(s_234), .O(gate389inter1));
  and2  gate2187(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2188(.a(s_234), .O(gate389inter3));
  inv1  gate2189(.a(s_235), .O(gate389inter4));
  nand2 gate2190(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2191(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2192(.a(G3), .O(gate389inter7));
  inv1  gate2193(.a(G1042), .O(gate389inter8));
  nand2 gate2194(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2195(.a(s_235), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2196(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2197(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2198(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate911(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate912(.a(gate394inter0), .b(s_52), .O(gate394inter1));
  and2  gate913(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate914(.a(s_52), .O(gate394inter3));
  inv1  gate915(.a(s_53), .O(gate394inter4));
  nand2 gate916(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate917(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate918(.a(G8), .O(gate394inter7));
  inv1  gate919(.a(G1057), .O(gate394inter8));
  nand2 gate920(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate921(.a(s_53), .b(gate394inter3), .O(gate394inter10));
  nor2  gate922(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate923(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate924(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate561(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate562(.a(gate395inter0), .b(s_2), .O(gate395inter1));
  and2  gate563(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate564(.a(s_2), .O(gate395inter3));
  inv1  gate565(.a(s_3), .O(gate395inter4));
  nand2 gate566(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate567(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate568(.a(G9), .O(gate395inter7));
  inv1  gate569(.a(G1060), .O(gate395inter8));
  nand2 gate570(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate571(.a(s_3), .b(gate395inter3), .O(gate395inter10));
  nor2  gate572(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate573(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate574(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2101(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2102(.a(gate397inter0), .b(s_222), .O(gate397inter1));
  and2  gate2103(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2104(.a(s_222), .O(gate397inter3));
  inv1  gate2105(.a(s_223), .O(gate397inter4));
  nand2 gate2106(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2107(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2108(.a(G11), .O(gate397inter7));
  inv1  gate2109(.a(G1066), .O(gate397inter8));
  nand2 gate2110(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2111(.a(s_223), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2112(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2113(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2114(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1919(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1920(.a(gate399inter0), .b(s_196), .O(gate399inter1));
  and2  gate1921(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1922(.a(s_196), .O(gate399inter3));
  inv1  gate1923(.a(s_197), .O(gate399inter4));
  nand2 gate1924(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1925(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1926(.a(G13), .O(gate399inter7));
  inv1  gate1927(.a(G1072), .O(gate399inter8));
  nand2 gate1928(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1929(.a(s_197), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1930(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1931(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1932(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1639(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1640(.a(gate400inter0), .b(s_156), .O(gate400inter1));
  and2  gate1641(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1642(.a(s_156), .O(gate400inter3));
  inv1  gate1643(.a(s_157), .O(gate400inter4));
  nand2 gate1644(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1645(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1646(.a(G14), .O(gate400inter7));
  inv1  gate1647(.a(G1075), .O(gate400inter8));
  nand2 gate1648(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1649(.a(s_157), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1650(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1651(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1652(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1723(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1724(.a(gate401inter0), .b(s_168), .O(gate401inter1));
  and2  gate1725(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1726(.a(s_168), .O(gate401inter3));
  inv1  gate1727(.a(s_169), .O(gate401inter4));
  nand2 gate1728(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1729(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1730(.a(G15), .O(gate401inter7));
  inv1  gate1731(.a(G1078), .O(gate401inter8));
  nand2 gate1732(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1733(.a(s_169), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1734(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1735(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1736(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1233(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1234(.a(gate402inter0), .b(s_98), .O(gate402inter1));
  and2  gate1235(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1236(.a(s_98), .O(gate402inter3));
  inv1  gate1237(.a(s_99), .O(gate402inter4));
  nand2 gate1238(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1239(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1240(.a(G16), .O(gate402inter7));
  inv1  gate1241(.a(G1081), .O(gate402inter8));
  nand2 gate1242(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1243(.a(s_99), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1244(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1245(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1246(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1457(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1458(.a(gate406inter0), .b(s_130), .O(gate406inter1));
  and2  gate1459(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1460(.a(s_130), .O(gate406inter3));
  inv1  gate1461(.a(s_131), .O(gate406inter4));
  nand2 gate1462(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1463(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1464(.a(G20), .O(gate406inter7));
  inv1  gate1465(.a(G1093), .O(gate406inter8));
  nand2 gate1466(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1467(.a(s_131), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1468(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1469(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1470(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate841(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate842(.a(gate407inter0), .b(s_42), .O(gate407inter1));
  and2  gate843(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate844(.a(s_42), .O(gate407inter3));
  inv1  gate845(.a(s_43), .O(gate407inter4));
  nand2 gate846(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate847(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate848(.a(G21), .O(gate407inter7));
  inv1  gate849(.a(G1096), .O(gate407inter8));
  nand2 gate850(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate851(.a(s_43), .b(gate407inter3), .O(gate407inter10));
  nor2  gate852(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate853(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate854(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1947(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1948(.a(gate408inter0), .b(s_200), .O(gate408inter1));
  and2  gate1949(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1950(.a(s_200), .O(gate408inter3));
  inv1  gate1951(.a(s_201), .O(gate408inter4));
  nand2 gate1952(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1953(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1954(.a(G22), .O(gate408inter7));
  inv1  gate1955(.a(G1099), .O(gate408inter8));
  nand2 gate1956(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1957(.a(s_201), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1958(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1959(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1960(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1961(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1962(.a(gate409inter0), .b(s_202), .O(gate409inter1));
  and2  gate1963(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1964(.a(s_202), .O(gate409inter3));
  inv1  gate1965(.a(s_203), .O(gate409inter4));
  nand2 gate1966(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1967(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1968(.a(G23), .O(gate409inter7));
  inv1  gate1969(.a(G1102), .O(gate409inter8));
  nand2 gate1970(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1971(.a(s_203), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1972(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1973(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1974(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1289(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1290(.a(gate410inter0), .b(s_106), .O(gate410inter1));
  and2  gate1291(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1292(.a(s_106), .O(gate410inter3));
  inv1  gate1293(.a(s_107), .O(gate410inter4));
  nand2 gate1294(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1295(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1296(.a(G24), .O(gate410inter7));
  inv1  gate1297(.a(G1105), .O(gate410inter8));
  nand2 gate1298(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1299(.a(s_107), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1300(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1301(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1302(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate799(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate800(.a(gate412inter0), .b(s_36), .O(gate412inter1));
  and2  gate801(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate802(.a(s_36), .O(gate412inter3));
  inv1  gate803(.a(s_37), .O(gate412inter4));
  nand2 gate804(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate805(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate806(.a(G26), .O(gate412inter7));
  inv1  gate807(.a(G1111), .O(gate412inter8));
  nand2 gate808(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate809(.a(s_37), .b(gate412inter3), .O(gate412inter10));
  nor2  gate810(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate811(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate812(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2227(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2228(.a(gate419inter0), .b(s_240), .O(gate419inter1));
  and2  gate2229(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2230(.a(s_240), .O(gate419inter3));
  inv1  gate2231(.a(s_241), .O(gate419inter4));
  nand2 gate2232(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2233(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2234(.a(G1), .O(gate419inter7));
  inv1  gate2235(.a(G1132), .O(gate419inter8));
  nand2 gate2236(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2237(.a(s_241), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2238(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2239(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2240(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1555(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1556(.a(gate421inter0), .b(s_144), .O(gate421inter1));
  and2  gate1557(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1558(.a(s_144), .O(gate421inter3));
  inv1  gate1559(.a(s_145), .O(gate421inter4));
  nand2 gate1560(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1561(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1562(.a(G2), .O(gate421inter7));
  inv1  gate1563(.a(G1135), .O(gate421inter8));
  nand2 gate1564(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1565(.a(s_145), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1566(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1567(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1568(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2297(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2298(.a(gate422inter0), .b(s_250), .O(gate422inter1));
  and2  gate2299(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2300(.a(s_250), .O(gate422inter3));
  inv1  gate2301(.a(s_251), .O(gate422inter4));
  nand2 gate2302(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2303(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2304(.a(G1039), .O(gate422inter7));
  inv1  gate2305(.a(G1135), .O(gate422inter8));
  nand2 gate2306(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2307(.a(s_251), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2308(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2309(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2310(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2073(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2074(.a(gate426inter0), .b(s_218), .O(gate426inter1));
  and2  gate2075(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2076(.a(s_218), .O(gate426inter3));
  inv1  gate2077(.a(s_219), .O(gate426inter4));
  nand2 gate2078(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2079(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2080(.a(G1045), .O(gate426inter7));
  inv1  gate2081(.a(G1141), .O(gate426inter8));
  nand2 gate2082(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2083(.a(s_219), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2084(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2085(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2086(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate981(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate982(.a(gate434inter0), .b(s_62), .O(gate434inter1));
  and2  gate983(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate984(.a(s_62), .O(gate434inter3));
  inv1  gate985(.a(s_63), .O(gate434inter4));
  nand2 gate986(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate987(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate988(.a(G1057), .O(gate434inter7));
  inv1  gate989(.a(G1153), .O(gate434inter8));
  nand2 gate990(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate991(.a(s_63), .b(gate434inter3), .O(gate434inter10));
  nor2  gate992(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate993(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate994(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1065(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1066(.a(gate438inter0), .b(s_74), .O(gate438inter1));
  and2  gate1067(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1068(.a(s_74), .O(gate438inter3));
  inv1  gate1069(.a(s_75), .O(gate438inter4));
  nand2 gate1070(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1071(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1072(.a(G1063), .O(gate438inter7));
  inv1  gate1073(.a(G1159), .O(gate438inter8));
  nand2 gate1074(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1075(.a(s_75), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1076(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1077(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1078(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1569(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1570(.a(gate442inter0), .b(s_146), .O(gate442inter1));
  and2  gate1571(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1572(.a(s_146), .O(gate442inter3));
  inv1  gate1573(.a(s_147), .O(gate442inter4));
  nand2 gate1574(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1575(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1576(.a(G1069), .O(gate442inter7));
  inv1  gate1577(.a(G1165), .O(gate442inter8));
  nand2 gate1578(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1579(.a(s_147), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1580(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1581(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1582(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1751(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1752(.a(gate445inter0), .b(s_172), .O(gate445inter1));
  and2  gate1753(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1754(.a(s_172), .O(gate445inter3));
  inv1  gate1755(.a(s_173), .O(gate445inter4));
  nand2 gate1756(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1757(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1758(.a(G14), .O(gate445inter7));
  inv1  gate1759(.a(G1171), .O(gate445inter8));
  nand2 gate1760(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1761(.a(s_173), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1762(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1763(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1764(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate897(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate898(.a(gate450inter0), .b(s_50), .O(gate450inter1));
  and2  gate899(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate900(.a(s_50), .O(gate450inter3));
  inv1  gate901(.a(s_51), .O(gate450inter4));
  nand2 gate902(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate903(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate904(.a(G1081), .O(gate450inter7));
  inv1  gate905(.a(G1177), .O(gate450inter8));
  nand2 gate906(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate907(.a(s_51), .b(gate450inter3), .O(gate450inter10));
  nor2  gate908(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate909(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate910(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1807(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1808(.a(gate453inter0), .b(s_180), .O(gate453inter1));
  and2  gate1809(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1810(.a(s_180), .O(gate453inter3));
  inv1  gate1811(.a(s_181), .O(gate453inter4));
  nand2 gate1812(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1813(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1814(.a(G18), .O(gate453inter7));
  inv1  gate1815(.a(G1183), .O(gate453inter8));
  nand2 gate1816(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1817(.a(s_181), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1818(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1819(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1820(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate771(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate772(.a(gate454inter0), .b(s_32), .O(gate454inter1));
  and2  gate773(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate774(.a(s_32), .O(gate454inter3));
  inv1  gate775(.a(s_33), .O(gate454inter4));
  nand2 gate776(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate777(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate778(.a(G1087), .O(gate454inter7));
  inv1  gate779(.a(G1183), .O(gate454inter8));
  nand2 gate780(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate781(.a(s_33), .b(gate454inter3), .O(gate454inter10));
  nor2  gate782(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate783(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate784(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1093(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1094(.a(gate456inter0), .b(s_78), .O(gate456inter1));
  and2  gate1095(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1096(.a(s_78), .O(gate456inter3));
  inv1  gate1097(.a(s_79), .O(gate456inter4));
  nand2 gate1098(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1099(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1100(.a(G1090), .O(gate456inter7));
  inv1  gate1101(.a(G1186), .O(gate456inter8));
  nand2 gate1102(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1103(.a(s_79), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1104(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1105(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1106(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate2241(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2242(.a(gate457inter0), .b(s_242), .O(gate457inter1));
  and2  gate2243(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2244(.a(s_242), .O(gate457inter3));
  inv1  gate2245(.a(s_243), .O(gate457inter4));
  nand2 gate2246(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2247(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2248(.a(G20), .O(gate457inter7));
  inv1  gate2249(.a(G1189), .O(gate457inter8));
  nand2 gate2250(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2251(.a(s_243), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2252(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2253(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2254(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1695(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1696(.a(gate461inter0), .b(s_164), .O(gate461inter1));
  and2  gate1697(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1698(.a(s_164), .O(gate461inter3));
  inv1  gate1699(.a(s_165), .O(gate461inter4));
  nand2 gate1700(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1701(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1702(.a(G22), .O(gate461inter7));
  inv1  gate1703(.a(G1195), .O(gate461inter8));
  nand2 gate1704(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1705(.a(s_165), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1706(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1707(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1708(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate1163(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1164(.a(gate462inter0), .b(s_88), .O(gate462inter1));
  and2  gate1165(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1166(.a(s_88), .O(gate462inter3));
  inv1  gate1167(.a(s_89), .O(gate462inter4));
  nand2 gate1168(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1169(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1170(.a(G1099), .O(gate462inter7));
  inv1  gate1171(.a(G1195), .O(gate462inter8));
  nand2 gate1172(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1173(.a(s_89), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1174(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1175(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1176(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1247(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1248(.a(gate463inter0), .b(s_100), .O(gate463inter1));
  and2  gate1249(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1250(.a(s_100), .O(gate463inter3));
  inv1  gate1251(.a(s_101), .O(gate463inter4));
  nand2 gate1252(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1253(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1254(.a(G23), .O(gate463inter7));
  inv1  gate1255(.a(G1198), .O(gate463inter8));
  nand2 gate1256(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1257(.a(s_101), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1258(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1259(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1260(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1471(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1472(.a(gate476inter0), .b(s_132), .O(gate476inter1));
  and2  gate1473(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1474(.a(s_132), .O(gate476inter3));
  inv1  gate1475(.a(s_133), .O(gate476inter4));
  nand2 gate1476(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1477(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1478(.a(G1120), .O(gate476inter7));
  inv1  gate1479(.a(G1216), .O(gate476inter8));
  nand2 gate1480(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1481(.a(s_133), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1482(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1483(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1484(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1527(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1528(.a(gate481inter0), .b(s_140), .O(gate481inter1));
  and2  gate1529(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1530(.a(s_140), .O(gate481inter3));
  inv1  gate1531(.a(s_141), .O(gate481inter4));
  nand2 gate1532(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1533(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1534(.a(G32), .O(gate481inter7));
  inv1  gate1535(.a(G1225), .O(gate481inter8));
  nand2 gate1536(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1537(.a(s_141), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1538(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1539(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1540(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate645(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate646(.a(gate483inter0), .b(s_14), .O(gate483inter1));
  and2  gate647(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate648(.a(s_14), .O(gate483inter3));
  inv1  gate649(.a(s_15), .O(gate483inter4));
  nand2 gate650(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate651(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate652(.a(G1228), .O(gate483inter7));
  inv1  gate653(.a(G1229), .O(gate483inter8));
  nand2 gate654(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate655(.a(s_15), .b(gate483inter3), .O(gate483inter10));
  nor2  gate656(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate657(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate658(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate2031(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2032(.a(gate487inter0), .b(s_212), .O(gate487inter1));
  and2  gate2033(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2034(.a(s_212), .O(gate487inter3));
  inv1  gate2035(.a(s_213), .O(gate487inter4));
  nand2 gate2036(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2037(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2038(.a(G1236), .O(gate487inter7));
  inv1  gate2039(.a(G1237), .O(gate487inter8));
  nand2 gate2040(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2041(.a(s_213), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2042(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2043(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2044(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1009(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1010(.a(gate490inter0), .b(s_66), .O(gate490inter1));
  and2  gate1011(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1012(.a(s_66), .O(gate490inter3));
  inv1  gate1013(.a(s_67), .O(gate490inter4));
  nand2 gate1014(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1015(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1016(.a(G1242), .O(gate490inter7));
  inv1  gate1017(.a(G1243), .O(gate490inter8));
  nand2 gate1018(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1019(.a(s_67), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1020(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1021(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1022(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate2143(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2144(.a(gate491inter0), .b(s_228), .O(gate491inter1));
  and2  gate2145(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2146(.a(s_228), .O(gate491inter3));
  inv1  gate2147(.a(s_229), .O(gate491inter4));
  nand2 gate2148(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2149(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2150(.a(G1244), .O(gate491inter7));
  inv1  gate2151(.a(G1245), .O(gate491inter8));
  nand2 gate2152(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2153(.a(s_229), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2154(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2155(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2156(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1387(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1388(.a(gate492inter0), .b(s_120), .O(gate492inter1));
  and2  gate1389(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1390(.a(s_120), .O(gate492inter3));
  inv1  gate1391(.a(s_121), .O(gate492inter4));
  nand2 gate1392(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1393(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1394(.a(G1246), .O(gate492inter7));
  inv1  gate1395(.a(G1247), .O(gate492inter8));
  nand2 gate1396(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1397(.a(s_121), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1398(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1399(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1400(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1373(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1374(.a(gate497inter0), .b(s_118), .O(gate497inter1));
  and2  gate1375(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1376(.a(s_118), .O(gate497inter3));
  inv1  gate1377(.a(s_119), .O(gate497inter4));
  nand2 gate1378(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1379(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1380(.a(G1256), .O(gate497inter7));
  inv1  gate1381(.a(G1257), .O(gate497inter8));
  nand2 gate1382(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1383(.a(s_119), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1384(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1385(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1386(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1597(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1598(.a(gate505inter0), .b(s_150), .O(gate505inter1));
  and2  gate1599(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1600(.a(s_150), .O(gate505inter3));
  inv1  gate1601(.a(s_151), .O(gate505inter4));
  nand2 gate1602(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1603(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1604(.a(G1272), .O(gate505inter7));
  inv1  gate1605(.a(G1273), .O(gate505inter8));
  nand2 gate1606(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1607(.a(s_151), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1608(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1609(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1610(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate743(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate744(.a(gate508inter0), .b(s_28), .O(gate508inter1));
  and2  gate745(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate746(.a(s_28), .O(gate508inter3));
  inv1  gate747(.a(s_29), .O(gate508inter4));
  nand2 gate748(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate749(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate750(.a(G1278), .O(gate508inter7));
  inv1  gate751(.a(G1279), .O(gate508inter8));
  nand2 gate752(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate753(.a(s_29), .b(gate508inter3), .O(gate508inter10));
  nor2  gate754(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate755(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate756(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1037(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1038(.a(gate513inter0), .b(s_70), .O(gate513inter1));
  and2  gate1039(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1040(.a(s_70), .O(gate513inter3));
  inv1  gate1041(.a(s_71), .O(gate513inter4));
  nand2 gate1042(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1043(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1044(.a(G1288), .O(gate513inter7));
  inv1  gate1045(.a(G1289), .O(gate513inter8));
  nand2 gate1046(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1047(.a(s_71), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1048(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1049(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1050(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule