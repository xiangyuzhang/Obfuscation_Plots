module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1975(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1976(.a(gate9inter0), .b(s_204), .O(gate9inter1));
  and2  gate1977(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1978(.a(s_204), .O(gate9inter3));
  inv1  gate1979(.a(s_205), .O(gate9inter4));
  nand2 gate1980(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1981(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1982(.a(G1), .O(gate9inter7));
  inv1  gate1983(.a(G2), .O(gate9inter8));
  nand2 gate1984(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1985(.a(s_205), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1986(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1987(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1988(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1373(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1374(.a(gate14inter0), .b(s_118), .O(gate14inter1));
  and2  gate1375(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1376(.a(s_118), .O(gate14inter3));
  inv1  gate1377(.a(s_119), .O(gate14inter4));
  nand2 gate1378(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1379(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1380(.a(G11), .O(gate14inter7));
  inv1  gate1381(.a(G12), .O(gate14inter8));
  nand2 gate1382(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1383(.a(s_119), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1384(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1385(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1386(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate2535(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2536(.a(gate15inter0), .b(s_284), .O(gate15inter1));
  and2  gate2537(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2538(.a(s_284), .O(gate15inter3));
  inv1  gate2539(.a(s_285), .O(gate15inter4));
  nand2 gate2540(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2541(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2542(.a(G13), .O(gate15inter7));
  inv1  gate2543(.a(G14), .O(gate15inter8));
  nand2 gate2544(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2545(.a(s_285), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2546(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2547(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2548(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2297(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2298(.a(gate21inter0), .b(s_250), .O(gate21inter1));
  and2  gate2299(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2300(.a(s_250), .O(gate21inter3));
  inv1  gate2301(.a(s_251), .O(gate21inter4));
  nand2 gate2302(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2303(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2304(.a(G25), .O(gate21inter7));
  inv1  gate2305(.a(G26), .O(gate21inter8));
  nand2 gate2306(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2307(.a(s_251), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2308(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2309(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2310(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1429(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1430(.a(gate22inter0), .b(s_126), .O(gate22inter1));
  and2  gate1431(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1432(.a(s_126), .O(gate22inter3));
  inv1  gate1433(.a(s_127), .O(gate22inter4));
  nand2 gate1434(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1435(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1436(.a(G27), .O(gate22inter7));
  inv1  gate1437(.a(G28), .O(gate22inter8));
  nand2 gate1438(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1439(.a(s_127), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1440(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1441(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1442(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1919(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1920(.a(gate23inter0), .b(s_196), .O(gate23inter1));
  and2  gate1921(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1922(.a(s_196), .O(gate23inter3));
  inv1  gate1923(.a(s_197), .O(gate23inter4));
  nand2 gate1924(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1925(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1926(.a(G29), .O(gate23inter7));
  inv1  gate1927(.a(G30), .O(gate23inter8));
  nand2 gate1928(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1929(.a(s_197), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1930(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1931(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1932(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1317(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1318(.a(gate25inter0), .b(s_110), .O(gate25inter1));
  and2  gate1319(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1320(.a(s_110), .O(gate25inter3));
  inv1  gate1321(.a(s_111), .O(gate25inter4));
  nand2 gate1322(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1323(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1324(.a(G1), .O(gate25inter7));
  inv1  gate1325(.a(G5), .O(gate25inter8));
  nand2 gate1326(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1327(.a(s_111), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1328(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1329(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1330(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate855(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate856(.a(gate27inter0), .b(s_44), .O(gate27inter1));
  and2  gate857(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate858(.a(s_44), .O(gate27inter3));
  inv1  gate859(.a(s_45), .O(gate27inter4));
  nand2 gate860(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate861(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate862(.a(G2), .O(gate27inter7));
  inv1  gate863(.a(G6), .O(gate27inter8));
  nand2 gate864(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate865(.a(s_45), .b(gate27inter3), .O(gate27inter10));
  nor2  gate866(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate867(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate868(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2227(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2228(.a(gate29inter0), .b(s_240), .O(gate29inter1));
  and2  gate2229(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2230(.a(s_240), .O(gate29inter3));
  inv1  gate2231(.a(s_241), .O(gate29inter4));
  nand2 gate2232(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2233(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2234(.a(G3), .O(gate29inter7));
  inv1  gate2235(.a(G7), .O(gate29inter8));
  nand2 gate2236(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2237(.a(s_241), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2238(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2239(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2240(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2213(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2214(.a(gate33inter0), .b(s_238), .O(gate33inter1));
  and2  gate2215(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2216(.a(s_238), .O(gate33inter3));
  inv1  gate2217(.a(s_239), .O(gate33inter4));
  nand2 gate2218(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2219(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2220(.a(G17), .O(gate33inter7));
  inv1  gate2221(.a(G21), .O(gate33inter8));
  nand2 gate2222(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2223(.a(s_239), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2224(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2225(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2226(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2367(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2368(.a(gate35inter0), .b(s_260), .O(gate35inter1));
  and2  gate2369(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2370(.a(s_260), .O(gate35inter3));
  inv1  gate2371(.a(s_261), .O(gate35inter4));
  nand2 gate2372(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2373(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2374(.a(G18), .O(gate35inter7));
  inv1  gate2375(.a(G22), .O(gate35inter8));
  nand2 gate2376(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2377(.a(s_261), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2378(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2379(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2380(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1261(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1262(.a(gate38inter0), .b(s_102), .O(gate38inter1));
  and2  gate1263(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1264(.a(s_102), .O(gate38inter3));
  inv1  gate1265(.a(s_103), .O(gate38inter4));
  nand2 gate1266(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1267(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1268(.a(G27), .O(gate38inter7));
  inv1  gate1269(.a(G31), .O(gate38inter8));
  nand2 gate1270(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1271(.a(s_103), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1272(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1273(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1274(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2381(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2382(.a(gate39inter0), .b(s_262), .O(gate39inter1));
  and2  gate2383(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2384(.a(s_262), .O(gate39inter3));
  inv1  gate2385(.a(s_263), .O(gate39inter4));
  nand2 gate2386(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2387(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2388(.a(G20), .O(gate39inter7));
  inv1  gate2389(.a(G24), .O(gate39inter8));
  nand2 gate2390(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2391(.a(s_263), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2392(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2393(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2394(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2185(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2186(.a(gate42inter0), .b(s_234), .O(gate42inter1));
  and2  gate2187(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2188(.a(s_234), .O(gate42inter3));
  inv1  gate2189(.a(s_235), .O(gate42inter4));
  nand2 gate2190(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2191(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2192(.a(G2), .O(gate42inter7));
  inv1  gate2193(.a(G266), .O(gate42inter8));
  nand2 gate2194(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2195(.a(s_235), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2196(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2197(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2198(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1597(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1598(.a(gate45inter0), .b(s_150), .O(gate45inter1));
  and2  gate1599(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1600(.a(s_150), .O(gate45inter3));
  inv1  gate1601(.a(s_151), .O(gate45inter4));
  nand2 gate1602(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1603(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1604(.a(G5), .O(gate45inter7));
  inv1  gate1605(.a(G272), .O(gate45inter8));
  nand2 gate1606(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1607(.a(s_151), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1608(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1609(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1610(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1149(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1150(.a(gate46inter0), .b(s_86), .O(gate46inter1));
  and2  gate1151(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1152(.a(s_86), .O(gate46inter3));
  inv1  gate1153(.a(s_87), .O(gate46inter4));
  nand2 gate1154(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1155(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1156(.a(G6), .O(gate46inter7));
  inv1  gate1157(.a(G272), .O(gate46inter8));
  nand2 gate1158(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1159(.a(s_87), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1160(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1161(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1162(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1877(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1878(.a(gate47inter0), .b(s_190), .O(gate47inter1));
  and2  gate1879(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1880(.a(s_190), .O(gate47inter3));
  inv1  gate1881(.a(s_191), .O(gate47inter4));
  nand2 gate1882(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1883(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1884(.a(G7), .O(gate47inter7));
  inv1  gate1885(.a(G275), .O(gate47inter8));
  nand2 gate1886(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1887(.a(s_191), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1888(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1889(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1890(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1401(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1402(.a(gate50inter0), .b(s_122), .O(gate50inter1));
  and2  gate1403(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1404(.a(s_122), .O(gate50inter3));
  inv1  gate1405(.a(s_123), .O(gate50inter4));
  nand2 gate1406(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1407(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1408(.a(G10), .O(gate50inter7));
  inv1  gate1409(.a(G278), .O(gate50inter8));
  nand2 gate1410(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1411(.a(s_123), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1412(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1413(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1414(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1177(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1178(.a(gate57inter0), .b(s_90), .O(gate57inter1));
  and2  gate1179(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1180(.a(s_90), .O(gate57inter3));
  inv1  gate1181(.a(s_91), .O(gate57inter4));
  nand2 gate1182(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1183(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1184(.a(G17), .O(gate57inter7));
  inv1  gate1185(.a(G290), .O(gate57inter8));
  nand2 gate1186(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1187(.a(s_91), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1188(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1189(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1190(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1135(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1136(.a(gate58inter0), .b(s_84), .O(gate58inter1));
  and2  gate1137(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1138(.a(s_84), .O(gate58inter3));
  inv1  gate1139(.a(s_85), .O(gate58inter4));
  nand2 gate1140(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1141(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1142(.a(G18), .O(gate58inter7));
  inv1  gate1143(.a(G290), .O(gate58inter8));
  nand2 gate1144(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1145(.a(s_85), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1146(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1147(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1148(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1793(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1794(.a(gate59inter0), .b(s_178), .O(gate59inter1));
  and2  gate1795(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1796(.a(s_178), .O(gate59inter3));
  inv1  gate1797(.a(s_179), .O(gate59inter4));
  nand2 gate1798(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1799(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1800(.a(G19), .O(gate59inter7));
  inv1  gate1801(.a(G293), .O(gate59inter8));
  nand2 gate1802(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1803(.a(s_179), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1804(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1805(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1806(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1569(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1570(.a(gate71inter0), .b(s_146), .O(gate71inter1));
  and2  gate1571(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1572(.a(s_146), .O(gate71inter3));
  inv1  gate1573(.a(s_147), .O(gate71inter4));
  nand2 gate1574(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1575(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1576(.a(G31), .O(gate71inter7));
  inv1  gate1577(.a(G311), .O(gate71inter8));
  nand2 gate1578(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1579(.a(s_147), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1580(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1581(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1582(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1219(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1220(.a(gate72inter0), .b(s_96), .O(gate72inter1));
  and2  gate1221(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1222(.a(s_96), .O(gate72inter3));
  inv1  gate1223(.a(s_97), .O(gate72inter4));
  nand2 gate1224(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1225(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1226(.a(G32), .O(gate72inter7));
  inv1  gate1227(.a(G311), .O(gate72inter8));
  nand2 gate1228(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1229(.a(s_97), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1230(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1231(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1232(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate897(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate898(.a(gate75inter0), .b(s_50), .O(gate75inter1));
  and2  gate899(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate900(.a(s_50), .O(gate75inter3));
  inv1  gate901(.a(s_51), .O(gate75inter4));
  nand2 gate902(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate903(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate904(.a(G9), .O(gate75inter7));
  inv1  gate905(.a(G317), .O(gate75inter8));
  nand2 gate906(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate907(.a(s_51), .b(gate75inter3), .O(gate75inter10));
  nor2  gate908(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate909(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate910(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1443(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1444(.a(gate76inter0), .b(s_128), .O(gate76inter1));
  and2  gate1445(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1446(.a(s_128), .O(gate76inter3));
  inv1  gate1447(.a(s_129), .O(gate76inter4));
  nand2 gate1448(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1449(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1450(.a(G13), .O(gate76inter7));
  inv1  gate1451(.a(G317), .O(gate76inter8));
  nand2 gate1452(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1453(.a(s_129), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1454(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1455(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1456(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate981(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate982(.a(gate77inter0), .b(s_62), .O(gate77inter1));
  and2  gate983(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate984(.a(s_62), .O(gate77inter3));
  inv1  gate985(.a(s_63), .O(gate77inter4));
  nand2 gate986(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate987(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate988(.a(G2), .O(gate77inter7));
  inv1  gate989(.a(G320), .O(gate77inter8));
  nand2 gate990(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate991(.a(s_63), .b(gate77inter3), .O(gate77inter10));
  nor2  gate992(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate993(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate994(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate2241(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2242(.a(gate78inter0), .b(s_242), .O(gate78inter1));
  and2  gate2243(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2244(.a(s_242), .O(gate78inter3));
  inv1  gate2245(.a(s_243), .O(gate78inter4));
  nand2 gate2246(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2247(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2248(.a(G6), .O(gate78inter7));
  inv1  gate2249(.a(G320), .O(gate78inter8));
  nand2 gate2250(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2251(.a(s_243), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2252(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2253(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2254(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1681(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1682(.a(gate80inter0), .b(s_162), .O(gate80inter1));
  and2  gate1683(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1684(.a(s_162), .O(gate80inter3));
  inv1  gate1685(.a(s_163), .O(gate80inter4));
  nand2 gate1686(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1687(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1688(.a(G14), .O(gate80inter7));
  inv1  gate1689(.a(G323), .O(gate80inter8));
  nand2 gate1690(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1691(.a(s_163), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1692(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1693(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1694(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2689(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2690(.a(gate81inter0), .b(s_306), .O(gate81inter1));
  and2  gate2691(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2692(.a(s_306), .O(gate81inter3));
  inv1  gate2693(.a(s_307), .O(gate81inter4));
  nand2 gate2694(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2695(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2696(.a(G3), .O(gate81inter7));
  inv1  gate2697(.a(G326), .O(gate81inter8));
  nand2 gate2698(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2699(.a(s_307), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2700(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2701(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2702(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate729(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate730(.a(gate90inter0), .b(s_26), .O(gate90inter1));
  and2  gate731(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate732(.a(s_26), .O(gate90inter3));
  inv1  gate733(.a(s_27), .O(gate90inter4));
  nand2 gate734(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate735(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate736(.a(G21), .O(gate90inter7));
  inv1  gate737(.a(G338), .O(gate90inter8));
  nand2 gate738(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate739(.a(s_27), .b(gate90inter3), .O(gate90inter10));
  nor2  gate740(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate741(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate742(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1247(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1248(.a(gate93inter0), .b(s_100), .O(gate93inter1));
  and2  gate1249(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1250(.a(s_100), .O(gate93inter3));
  inv1  gate1251(.a(s_101), .O(gate93inter4));
  nand2 gate1252(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1253(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1254(.a(G18), .O(gate93inter7));
  inv1  gate1255(.a(G344), .O(gate93inter8));
  nand2 gate1256(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1257(.a(s_101), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1258(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1259(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1260(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2143(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2144(.a(gate95inter0), .b(s_228), .O(gate95inter1));
  and2  gate2145(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2146(.a(s_228), .O(gate95inter3));
  inv1  gate2147(.a(s_229), .O(gate95inter4));
  nand2 gate2148(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2149(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2150(.a(G26), .O(gate95inter7));
  inv1  gate2151(.a(G347), .O(gate95inter8));
  nand2 gate2152(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2153(.a(s_229), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2154(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2155(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2156(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2675(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2676(.a(gate97inter0), .b(s_304), .O(gate97inter1));
  and2  gate2677(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2678(.a(s_304), .O(gate97inter3));
  inv1  gate2679(.a(s_305), .O(gate97inter4));
  nand2 gate2680(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2681(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2682(.a(G19), .O(gate97inter7));
  inv1  gate2683(.a(G350), .O(gate97inter8));
  nand2 gate2684(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2685(.a(s_305), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2686(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2687(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2688(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate799(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate800(.a(gate98inter0), .b(s_36), .O(gate98inter1));
  and2  gate801(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate802(.a(s_36), .O(gate98inter3));
  inv1  gate803(.a(s_37), .O(gate98inter4));
  nand2 gate804(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate805(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate806(.a(G23), .O(gate98inter7));
  inv1  gate807(.a(G350), .O(gate98inter8));
  nand2 gate808(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate809(.a(s_37), .b(gate98inter3), .O(gate98inter10));
  nor2  gate810(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate811(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate812(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1863(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1864(.a(gate100inter0), .b(s_188), .O(gate100inter1));
  and2  gate1865(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1866(.a(s_188), .O(gate100inter3));
  inv1  gate1867(.a(s_189), .O(gate100inter4));
  nand2 gate1868(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1869(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1870(.a(G31), .O(gate100inter7));
  inv1  gate1871(.a(G353), .O(gate100inter8));
  nand2 gate1872(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1873(.a(s_189), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1874(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1875(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1876(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1905(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1906(.a(gate102inter0), .b(s_194), .O(gate102inter1));
  and2  gate1907(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1908(.a(s_194), .O(gate102inter3));
  inv1  gate1909(.a(s_195), .O(gate102inter4));
  nand2 gate1910(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1911(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1912(.a(G24), .O(gate102inter7));
  inv1  gate1913(.a(G356), .O(gate102inter8));
  nand2 gate1914(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1915(.a(s_195), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1916(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1917(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1918(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1947(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1948(.a(gate109inter0), .b(s_200), .O(gate109inter1));
  and2  gate1949(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1950(.a(s_200), .O(gate109inter3));
  inv1  gate1951(.a(s_201), .O(gate109inter4));
  nand2 gate1952(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1953(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1954(.a(G370), .O(gate109inter7));
  inv1  gate1955(.a(G371), .O(gate109inter8));
  nand2 gate1956(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1957(.a(s_201), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1958(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1959(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1960(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2325(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2326(.a(gate115inter0), .b(s_254), .O(gate115inter1));
  and2  gate2327(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2328(.a(s_254), .O(gate115inter3));
  inv1  gate2329(.a(s_255), .O(gate115inter4));
  nand2 gate2330(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2331(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2332(.a(G382), .O(gate115inter7));
  inv1  gate2333(.a(G383), .O(gate115inter8));
  nand2 gate2334(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2335(.a(s_255), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2336(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2337(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2338(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1303(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1304(.a(gate118inter0), .b(s_108), .O(gate118inter1));
  and2  gate1305(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1306(.a(s_108), .O(gate118inter3));
  inv1  gate1307(.a(s_109), .O(gate118inter4));
  nand2 gate1308(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1309(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1310(.a(G388), .O(gate118inter7));
  inv1  gate1311(.a(G389), .O(gate118inter8));
  nand2 gate1312(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1313(.a(s_109), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1314(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1315(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1316(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate547(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate548(.a(gate119inter0), .b(s_0), .O(gate119inter1));
  and2  gate549(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate550(.a(s_0), .O(gate119inter3));
  inv1  gate551(.a(s_1), .O(gate119inter4));
  nand2 gate552(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate553(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate554(.a(G390), .O(gate119inter7));
  inv1  gate555(.a(G391), .O(gate119inter8));
  nand2 gate556(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate557(.a(s_1), .b(gate119inter3), .O(gate119inter10));
  nor2  gate558(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate559(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate560(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1555(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1556(.a(gate121inter0), .b(s_144), .O(gate121inter1));
  and2  gate1557(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1558(.a(s_144), .O(gate121inter3));
  inv1  gate1559(.a(s_145), .O(gate121inter4));
  nand2 gate1560(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1561(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1562(.a(G394), .O(gate121inter7));
  inv1  gate1563(.a(G395), .O(gate121inter8));
  nand2 gate1564(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1565(.a(s_145), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1566(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1567(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1568(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2493(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2494(.a(gate122inter0), .b(s_278), .O(gate122inter1));
  and2  gate2495(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2496(.a(s_278), .O(gate122inter3));
  inv1  gate2497(.a(s_279), .O(gate122inter4));
  nand2 gate2498(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2499(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2500(.a(G396), .O(gate122inter7));
  inv1  gate2501(.a(G397), .O(gate122inter8));
  nand2 gate2502(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2503(.a(s_279), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2504(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2505(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2506(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1345(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1346(.a(gate130inter0), .b(s_114), .O(gate130inter1));
  and2  gate1347(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1348(.a(s_114), .O(gate130inter3));
  inv1  gate1349(.a(s_115), .O(gate130inter4));
  nand2 gate1350(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1351(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1352(.a(G412), .O(gate130inter7));
  inv1  gate1353(.a(G413), .O(gate130inter8));
  nand2 gate1354(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1355(.a(s_115), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1356(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1357(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1358(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1541(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1542(.a(gate131inter0), .b(s_142), .O(gate131inter1));
  and2  gate1543(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1544(.a(s_142), .O(gate131inter3));
  inv1  gate1545(.a(s_143), .O(gate131inter4));
  nand2 gate1546(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1547(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1548(.a(G414), .O(gate131inter7));
  inv1  gate1549(.a(G415), .O(gate131inter8));
  nand2 gate1550(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1551(.a(s_143), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1552(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1553(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1554(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1835(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1836(.a(gate139inter0), .b(s_184), .O(gate139inter1));
  and2  gate1837(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1838(.a(s_184), .O(gate139inter3));
  inv1  gate1839(.a(s_185), .O(gate139inter4));
  nand2 gate1840(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1841(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1842(.a(G438), .O(gate139inter7));
  inv1  gate1843(.a(G441), .O(gate139inter8));
  nand2 gate1844(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1845(.a(s_185), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1846(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1847(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1848(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate687(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate688(.a(gate143inter0), .b(s_20), .O(gate143inter1));
  and2  gate689(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate690(.a(s_20), .O(gate143inter3));
  inv1  gate691(.a(s_21), .O(gate143inter4));
  nand2 gate692(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate693(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate694(.a(G462), .O(gate143inter7));
  inv1  gate695(.a(G465), .O(gate143inter8));
  nand2 gate696(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate697(.a(s_21), .b(gate143inter3), .O(gate143inter10));
  nor2  gate698(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate699(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate700(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1933(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1934(.a(gate144inter0), .b(s_198), .O(gate144inter1));
  and2  gate1935(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1936(.a(s_198), .O(gate144inter3));
  inv1  gate1937(.a(s_199), .O(gate144inter4));
  nand2 gate1938(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1939(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1940(.a(G468), .O(gate144inter7));
  inv1  gate1941(.a(G471), .O(gate144inter8));
  nand2 gate1942(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1943(.a(s_199), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1944(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1945(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1946(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2479(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2480(.a(gate146inter0), .b(s_276), .O(gate146inter1));
  and2  gate2481(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2482(.a(s_276), .O(gate146inter3));
  inv1  gate2483(.a(s_277), .O(gate146inter4));
  nand2 gate2484(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2485(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2486(.a(G480), .O(gate146inter7));
  inv1  gate2487(.a(G483), .O(gate146inter8));
  nand2 gate2488(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2489(.a(s_277), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2490(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2491(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2492(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1709(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1710(.a(gate148inter0), .b(s_166), .O(gate148inter1));
  and2  gate1711(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1712(.a(s_166), .O(gate148inter3));
  inv1  gate1713(.a(s_167), .O(gate148inter4));
  nand2 gate1714(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1715(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1716(.a(G492), .O(gate148inter7));
  inv1  gate1717(.a(G495), .O(gate148inter8));
  nand2 gate1718(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1719(.a(s_167), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1720(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1721(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1722(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2059(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2060(.a(gate156inter0), .b(s_216), .O(gate156inter1));
  and2  gate2061(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2062(.a(s_216), .O(gate156inter3));
  inv1  gate2063(.a(s_217), .O(gate156inter4));
  nand2 gate2064(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2065(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2066(.a(G435), .O(gate156inter7));
  inv1  gate2067(.a(G525), .O(gate156inter8));
  nand2 gate2068(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2069(.a(s_217), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2070(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2071(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2072(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate603(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate604(.a(gate157inter0), .b(s_8), .O(gate157inter1));
  and2  gate605(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate606(.a(s_8), .O(gate157inter3));
  inv1  gate607(.a(s_9), .O(gate157inter4));
  nand2 gate608(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate609(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate610(.a(G438), .O(gate157inter7));
  inv1  gate611(.a(G528), .O(gate157inter8));
  nand2 gate612(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate613(.a(s_9), .b(gate157inter3), .O(gate157inter10));
  nor2  gate614(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate615(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate616(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate645(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate646(.a(gate159inter0), .b(s_14), .O(gate159inter1));
  and2  gate647(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate648(.a(s_14), .O(gate159inter3));
  inv1  gate649(.a(s_15), .O(gate159inter4));
  nand2 gate650(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate651(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate652(.a(G444), .O(gate159inter7));
  inv1  gate653(.a(G531), .O(gate159inter8));
  nand2 gate654(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate655(.a(s_15), .b(gate159inter3), .O(gate159inter10));
  nor2  gate656(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate657(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate658(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2633(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2634(.a(gate162inter0), .b(s_298), .O(gate162inter1));
  and2  gate2635(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2636(.a(s_298), .O(gate162inter3));
  inv1  gate2637(.a(s_299), .O(gate162inter4));
  nand2 gate2638(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2639(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2640(.a(G453), .O(gate162inter7));
  inv1  gate2641(.a(G534), .O(gate162inter8));
  nand2 gate2642(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2643(.a(s_299), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2644(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2645(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2646(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2577(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2578(.a(gate165inter0), .b(s_290), .O(gate165inter1));
  and2  gate2579(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2580(.a(s_290), .O(gate165inter3));
  inv1  gate2581(.a(s_291), .O(gate165inter4));
  nand2 gate2582(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2583(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2584(.a(G462), .O(gate165inter7));
  inv1  gate2585(.a(G540), .O(gate165inter8));
  nand2 gate2586(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2587(.a(s_291), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2588(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2589(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2590(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1457(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1458(.a(gate168inter0), .b(s_130), .O(gate168inter1));
  and2  gate1459(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1460(.a(s_130), .O(gate168inter3));
  inv1  gate1461(.a(s_131), .O(gate168inter4));
  nand2 gate1462(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1463(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1464(.a(G471), .O(gate168inter7));
  inv1  gate1465(.a(G543), .O(gate168inter8));
  nand2 gate1466(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1467(.a(s_131), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1468(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1469(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1470(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2003(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2004(.a(gate171inter0), .b(s_208), .O(gate171inter1));
  and2  gate2005(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2006(.a(s_208), .O(gate171inter3));
  inv1  gate2007(.a(s_209), .O(gate171inter4));
  nand2 gate2008(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2009(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2010(.a(G480), .O(gate171inter7));
  inv1  gate2011(.a(G549), .O(gate171inter8));
  nand2 gate2012(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2013(.a(s_209), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2014(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2015(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2016(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2269(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2270(.a(gate172inter0), .b(s_246), .O(gate172inter1));
  and2  gate2271(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2272(.a(s_246), .O(gate172inter3));
  inv1  gate2273(.a(s_247), .O(gate172inter4));
  nand2 gate2274(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2275(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2276(.a(G483), .O(gate172inter7));
  inv1  gate2277(.a(G549), .O(gate172inter8));
  nand2 gate2278(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2279(.a(s_247), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2280(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2281(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2282(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2031(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2032(.a(gate173inter0), .b(s_212), .O(gate173inter1));
  and2  gate2033(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2034(.a(s_212), .O(gate173inter3));
  inv1  gate2035(.a(s_213), .O(gate173inter4));
  nand2 gate2036(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2037(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2038(.a(G486), .O(gate173inter7));
  inv1  gate2039(.a(G552), .O(gate173inter8));
  nand2 gate2040(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2041(.a(s_213), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2042(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2043(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2044(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2157(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2158(.a(gate174inter0), .b(s_230), .O(gate174inter1));
  and2  gate2159(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2160(.a(s_230), .O(gate174inter3));
  inv1  gate2161(.a(s_231), .O(gate174inter4));
  nand2 gate2162(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2163(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2164(.a(G489), .O(gate174inter7));
  inv1  gate2165(.a(G552), .O(gate174inter8));
  nand2 gate2166(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2167(.a(s_231), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2168(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2169(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2170(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2437(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2438(.a(gate175inter0), .b(s_270), .O(gate175inter1));
  and2  gate2439(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2440(.a(s_270), .O(gate175inter3));
  inv1  gate2441(.a(s_271), .O(gate175inter4));
  nand2 gate2442(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2443(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2444(.a(G492), .O(gate175inter7));
  inv1  gate2445(.a(G555), .O(gate175inter8));
  nand2 gate2446(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2447(.a(s_271), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2448(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2449(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2450(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate575(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate576(.a(gate178inter0), .b(s_4), .O(gate178inter1));
  and2  gate577(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate578(.a(s_4), .O(gate178inter3));
  inv1  gate579(.a(s_5), .O(gate178inter4));
  nand2 gate580(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate581(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate582(.a(G501), .O(gate178inter7));
  inv1  gate583(.a(G558), .O(gate178inter8));
  nand2 gate584(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate585(.a(s_5), .b(gate178inter3), .O(gate178inter10));
  nor2  gate586(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate587(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate588(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1387(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1388(.a(gate180inter0), .b(s_120), .O(gate180inter1));
  and2  gate1389(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1390(.a(s_120), .O(gate180inter3));
  inv1  gate1391(.a(s_121), .O(gate180inter4));
  nand2 gate1392(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1393(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1394(.a(G507), .O(gate180inter7));
  inv1  gate1395(.a(G561), .O(gate180inter8));
  nand2 gate1396(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1397(.a(s_121), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1398(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1399(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1400(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate631(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate632(.a(gate181inter0), .b(s_12), .O(gate181inter1));
  and2  gate633(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate634(.a(s_12), .O(gate181inter3));
  inv1  gate635(.a(s_13), .O(gate181inter4));
  nand2 gate636(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate637(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate638(.a(G510), .O(gate181inter7));
  inv1  gate639(.a(G564), .O(gate181inter8));
  nand2 gate640(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate641(.a(s_13), .b(gate181inter3), .O(gate181inter10));
  nor2  gate642(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate643(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate644(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1527(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1528(.a(gate182inter0), .b(s_140), .O(gate182inter1));
  and2  gate1529(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1530(.a(s_140), .O(gate182inter3));
  inv1  gate1531(.a(s_141), .O(gate182inter4));
  nand2 gate1532(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1533(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1534(.a(G513), .O(gate182inter7));
  inv1  gate1535(.a(G564), .O(gate182inter8));
  nand2 gate1536(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1537(.a(s_141), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1538(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1539(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1540(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2647(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2648(.a(gate184inter0), .b(s_300), .O(gate184inter1));
  and2  gate2649(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2650(.a(s_300), .O(gate184inter3));
  inv1  gate2651(.a(s_301), .O(gate184inter4));
  nand2 gate2652(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2653(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2654(.a(G519), .O(gate184inter7));
  inv1  gate2655(.a(G567), .O(gate184inter8));
  nand2 gate2656(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2657(.a(s_301), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2658(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2659(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2660(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate995(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate996(.a(gate188inter0), .b(s_64), .O(gate188inter1));
  and2  gate997(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate998(.a(s_64), .O(gate188inter3));
  inv1  gate999(.a(s_65), .O(gate188inter4));
  nand2 gate1000(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1001(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1002(.a(G576), .O(gate188inter7));
  inv1  gate1003(.a(G577), .O(gate188inter8));
  nand2 gate1004(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1005(.a(s_65), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1006(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1007(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1008(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2703(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2704(.a(gate191inter0), .b(s_308), .O(gate191inter1));
  and2  gate2705(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2706(.a(s_308), .O(gate191inter3));
  inv1  gate2707(.a(s_309), .O(gate191inter4));
  nand2 gate2708(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2709(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2710(.a(G582), .O(gate191inter7));
  inv1  gate2711(.a(G583), .O(gate191inter8));
  nand2 gate2712(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2713(.a(s_309), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2714(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2715(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2716(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2717(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2718(.a(gate192inter0), .b(s_310), .O(gate192inter1));
  and2  gate2719(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2720(.a(s_310), .O(gate192inter3));
  inv1  gate2721(.a(s_311), .O(gate192inter4));
  nand2 gate2722(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2723(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2724(.a(G584), .O(gate192inter7));
  inv1  gate2725(.a(G585), .O(gate192inter8));
  nand2 gate2726(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2727(.a(s_311), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2728(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2729(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2730(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate617(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate618(.a(gate196inter0), .b(s_10), .O(gate196inter1));
  and2  gate619(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate620(.a(s_10), .O(gate196inter3));
  inv1  gate621(.a(s_11), .O(gate196inter4));
  nand2 gate622(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate623(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate624(.a(G592), .O(gate196inter7));
  inv1  gate625(.a(G593), .O(gate196inter8));
  nand2 gate626(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate627(.a(s_11), .b(gate196inter3), .O(gate196inter10));
  nor2  gate628(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate629(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate630(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2423(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2424(.a(gate198inter0), .b(s_268), .O(gate198inter1));
  and2  gate2425(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2426(.a(s_268), .O(gate198inter3));
  inv1  gate2427(.a(s_269), .O(gate198inter4));
  nand2 gate2428(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2429(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2430(.a(G596), .O(gate198inter7));
  inv1  gate2431(.a(G597), .O(gate198inter8));
  nand2 gate2432(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2433(.a(s_269), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2434(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2435(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2436(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate841(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate842(.a(gate199inter0), .b(s_42), .O(gate199inter1));
  and2  gate843(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate844(.a(s_42), .O(gate199inter3));
  inv1  gate845(.a(s_43), .O(gate199inter4));
  nand2 gate846(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate847(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate848(.a(G598), .O(gate199inter7));
  inv1  gate849(.a(G599), .O(gate199inter8));
  nand2 gate850(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate851(.a(s_43), .b(gate199inter3), .O(gate199inter10));
  nor2  gate852(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate853(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate854(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1331(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1332(.a(gate202inter0), .b(s_112), .O(gate202inter1));
  and2  gate1333(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1334(.a(s_112), .O(gate202inter3));
  inv1  gate1335(.a(s_113), .O(gate202inter4));
  nand2 gate1336(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1337(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1338(.a(G612), .O(gate202inter7));
  inv1  gate1339(.a(G617), .O(gate202inter8));
  nand2 gate1340(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1341(.a(s_113), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1342(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1343(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1344(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1667(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1668(.a(gate211inter0), .b(s_160), .O(gate211inter1));
  and2  gate1669(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1670(.a(s_160), .O(gate211inter3));
  inv1  gate1671(.a(s_161), .O(gate211inter4));
  nand2 gate1672(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1673(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1674(.a(G612), .O(gate211inter7));
  inv1  gate1675(.a(G669), .O(gate211inter8));
  nand2 gate1676(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1677(.a(s_161), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1678(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1679(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1680(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate673(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate674(.a(gate214inter0), .b(s_18), .O(gate214inter1));
  and2  gate675(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate676(.a(s_18), .O(gate214inter3));
  inv1  gate677(.a(s_19), .O(gate214inter4));
  nand2 gate678(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate679(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate680(.a(G612), .O(gate214inter7));
  inv1  gate681(.a(G672), .O(gate214inter8));
  nand2 gate682(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate683(.a(s_19), .b(gate214inter3), .O(gate214inter10));
  nor2  gate684(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate685(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate686(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2199(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2200(.a(gate219inter0), .b(s_236), .O(gate219inter1));
  and2  gate2201(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2202(.a(s_236), .O(gate219inter3));
  inv1  gate2203(.a(s_237), .O(gate219inter4));
  nand2 gate2204(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2205(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2206(.a(G632), .O(gate219inter7));
  inv1  gate2207(.a(G681), .O(gate219inter8));
  nand2 gate2208(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2209(.a(s_237), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2210(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2211(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2212(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2591(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2592(.a(gate223inter0), .b(s_292), .O(gate223inter1));
  and2  gate2593(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2594(.a(s_292), .O(gate223inter3));
  inv1  gate2595(.a(s_293), .O(gate223inter4));
  nand2 gate2596(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2597(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2598(.a(G627), .O(gate223inter7));
  inv1  gate2599(.a(G687), .O(gate223inter8));
  nand2 gate2600(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2601(.a(s_293), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2602(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2603(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2604(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1751(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1752(.a(gate224inter0), .b(s_172), .O(gate224inter1));
  and2  gate1753(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1754(.a(s_172), .O(gate224inter3));
  inv1  gate1755(.a(s_173), .O(gate224inter4));
  nand2 gate1756(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1757(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1758(.a(G637), .O(gate224inter7));
  inv1  gate1759(.a(G687), .O(gate224inter8));
  nand2 gate1760(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1761(.a(s_173), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1762(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1763(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1764(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1163(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1164(.a(gate226inter0), .b(s_88), .O(gate226inter1));
  and2  gate1165(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1166(.a(s_88), .O(gate226inter3));
  inv1  gate1167(.a(s_89), .O(gate226inter4));
  nand2 gate1168(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1169(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1170(.a(G692), .O(gate226inter7));
  inv1  gate1171(.a(G693), .O(gate226inter8));
  nand2 gate1172(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1173(.a(s_89), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1174(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1175(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1176(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate911(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate912(.a(gate228inter0), .b(s_52), .O(gate228inter1));
  and2  gate913(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate914(.a(s_52), .O(gate228inter3));
  inv1  gate915(.a(s_53), .O(gate228inter4));
  nand2 gate916(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate917(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate918(.a(G696), .O(gate228inter7));
  inv1  gate919(.a(G697), .O(gate228inter8));
  nand2 gate920(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate921(.a(s_53), .b(gate228inter3), .O(gate228inter10));
  nor2  gate922(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate923(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate924(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate589(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate590(.a(gate229inter0), .b(s_6), .O(gate229inter1));
  and2  gate591(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate592(.a(s_6), .O(gate229inter3));
  inv1  gate593(.a(s_7), .O(gate229inter4));
  nand2 gate594(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate595(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate596(.a(G698), .O(gate229inter7));
  inv1  gate597(.a(G699), .O(gate229inter8));
  nand2 gate598(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate599(.a(s_7), .b(gate229inter3), .O(gate229inter10));
  nor2  gate600(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate601(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate602(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2283(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2284(.a(gate231inter0), .b(s_248), .O(gate231inter1));
  and2  gate2285(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2286(.a(s_248), .O(gate231inter3));
  inv1  gate2287(.a(s_249), .O(gate231inter4));
  nand2 gate2288(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2289(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2290(.a(G702), .O(gate231inter7));
  inv1  gate2291(.a(G703), .O(gate231inter8));
  nand2 gate2292(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2293(.a(s_249), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2294(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2295(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2296(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2353(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2354(.a(gate232inter0), .b(s_258), .O(gate232inter1));
  and2  gate2355(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2356(.a(s_258), .O(gate232inter3));
  inv1  gate2357(.a(s_259), .O(gate232inter4));
  nand2 gate2358(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2359(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2360(.a(G704), .O(gate232inter7));
  inv1  gate2361(.a(G705), .O(gate232inter8));
  nand2 gate2362(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2363(.a(s_259), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2364(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2365(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2366(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate869(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate870(.a(gate233inter0), .b(s_46), .O(gate233inter1));
  and2  gate871(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate872(.a(s_46), .O(gate233inter3));
  inv1  gate873(.a(s_47), .O(gate233inter4));
  nand2 gate874(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate875(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate876(.a(G242), .O(gate233inter7));
  inv1  gate877(.a(G718), .O(gate233inter8));
  nand2 gate878(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate879(.a(s_47), .b(gate233inter3), .O(gate233inter10));
  nor2  gate880(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate881(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate882(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate925(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate926(.a(gate235inter0), .b(s_54), .O(gate235inter1));
  and2  gate927(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate928(.a(s_54), .O(gate235inter3));
  inv1  gate929(.a(s_55), .O(gate235inter4));
  nand2 gate930(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate931(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate932(.a(G248), .O(gate235inter7));
  inv1  gate933(.a(G724), .O(gate235inter8));
  nand2 gate934(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate935(.a(s_55), .b(gate235inter3), .O(gate235inter10));
  nor2  gate936(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate937(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate938(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2087(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2088(.a(gate242inter0), .b(s_220), .O(gate242inter1));
  and2  gate2089(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2090(.a(s_220), .O(gate242inter3));
  inv1  gate2091(.a(s_221), .O(gate242inter4));
  nand2 gate2092(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2093(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2094(.a(G718), .O(gate242inter7));
  inv1  gate2095(.a(G730), .O(gate242inter8));
  nand2 gate2096(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2097(.a(s_221), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2098(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2099(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2100(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1289(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1290(.a(gate244inter0), .b(s_106), .O(gate244inter1));
  and2  gate1291(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1292(.a(s_106), .O(gate244inter3));
  inv1  gate1293(.a(s_107), .O(gate244inter4));
  nand2 gate1294(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1295(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1296(.a(G721), .O(gate244inter7));
  inv1  gate1297(.a(G733), .O(gate244inter8));
  nand2 gate1298(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1299(.a(s_107), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1300(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1301(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1302(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1359(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1360(.a(gate245inter0), .b(s_116), .O(gate245inter1));
  and2  gate1361(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1362(.a(s_116), .O(gate245inter3));
  inv1  gate1363(.a(s_117), .O(gate245inter4));
  nand2 gate1364(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1365(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1366(.a(G248), .O(gate245inter7));
  inv1  gate1367(.a(G736), .O(gate245inter8));
  nand2 gate1368(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1369(.a(s_117), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1370(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1371(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1372(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1849(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1850(.a(gate247inter0), .b(s_186), .O(gate247inter1));
  and2  gate1851(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1852(.a(s_186), .O(gate247inter3));
  inv1  gate1853(.a(s_187), .O(gate247inter4));
  nand2 gate1854(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1855(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1856(.a(G251), .O(gate247inter7));
  inv1  gate1857(.a(G739), .O(gate247inter8));
  nand2 gate1858(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1859(.a(s_187), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1860(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1861(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1862(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2521(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2522(.a(gate248inter0), .b(s_282), .O(gate248inter1));
  and2  gate2523(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2524(.a(s_282), .O(gate248inter3));
  inv1  gate2525(.a(s_283), .O(gate248inter4));
  nand2 gate2526(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2527(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2528(.a(G727), .O(gate248inter7));
  inv1  gate2529(.a(G739), .O(gate248inter8));
  nand2 gate2530(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2531(.a(s_283), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2532(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2533(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2534(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1891(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1892(.a(gate249inter0), .b(s_192), .O(gate249inter1));
  and2  gate1893(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1894(.a(s_192), .O(gate249inter3));
  inv1  gate1895(.a(s_193), .O(gate249inter4));
  nand2 gate1896(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1897(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1898(.a(G254), .O(gate249inter7));
  inv1  gate1899(.a(G742), .O(gate249inter8));
  nand2 gate1900(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1901(.a(s_193), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1902(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1903(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1904(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2017(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2018(.a(gate250inter0), .b(s_210), .O(gate250inter1));
  and2  gate2019(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2020(.a(s_210), .O(gate250inter3));
  inv1  gate2021(.a(s_211), .O(gate250inter4));
  nand2 gate2022(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2023(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2024(.a(G706), .O(gate250inter7));
  inv1  gate2025(.a(G742), .O(gate250inter8));
  nand2 gate2026(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2027(.a(s_211), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2028(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2029(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2030(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2619(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2620(.a(gate251inter0), .b(s_296), .O(gate251inter1));
  and2  gate2621(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2622(.a(s_296), .O(gate251inter3));
  inv1  gate2623(.a(s_297), .O(gate251inter4));
  nand2 gate2624(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2625(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2626(.a(G257), .O(gate251inter7));
  inv1  gate2627(.a(G745), .O(gate251inter8));
  nand2 gate2628(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2629(.a(s_297), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2630(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2631(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2632(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2073(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2074(.a(gate254inter0), .b(s_218), .O(gate254inter1));
  and2  gate2075(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2076(.a(s_218), .O(gate254inter3));
  inv1  gate2077(.a(s_219), .O(gate254inter4));
  nand2 gate2078(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2079(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2080(.a(G712), .O(gate254inter7));
  inv1  gate2081(.a(G748), .O(gate254inter8));
  nand2 gate2082(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2083(.a(s_219), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2084(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2085(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2086(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate659(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate660(.a(gate256inter0), .b(s_16), .O(gate256inter1));
  and2  gate661(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate662(.a(s_16), .O(gate256inter3));
  inv1  gate663(.a(s_17), .O(gate256inter4));
  nand2 gate664(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate665(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate666(.a(G715), .O(gate256inter7));
  inv1  gate667(.a(G751), .O(gate256inter8));
  nand2 gate668(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate669(.a(s_17), .b(gate256inter3), .O(gate256inter10));
  nor2  gate670(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate671(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate672(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1065(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1066(.a(gate261inter0), .b(s_74), .O(gate261inter1));
  and2  gate1067(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1068(.a(s_74), .O(gate261inter3));
  inv1  gate1069(.a(s_75), .O(gate261inter4));
  nand2 gate1070(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1071(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1072(.a(G762), .O(gate261inter7));
  inv1  gate1073(.a(G763), .O(gate261inter8));
  nand2 gate1074(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1075(.a(s_75), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1076(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1077(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1078(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1415(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1416(.a(gate263inter0), .b(s_124), .O(gate263inter1));
  and2  gate1417(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1418(.a(s_124), .O(gate263inter3));
  inv1  gate1419(.a(s_125), .O(gate263inter4));
  nand2 gate1420(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1421(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1422(.a(G766), .O(gate263inter7));
  inv1  gate1423(.a(G767), .O(gate263inter8));
  nand2 gate1424(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1425(.a(s_125), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1426(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1427(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1428(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate883(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate884(.a(gate264inter0), .b(s_48), .O(gate264inter1));
  and2  gate885(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate886(.a(s_48), .O(gate264inter3));
  inv1  gate887(.a(s_49), .O(gate264inter4));
  nand2 gate888(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate889(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate890(.a(G768), .O(gate264inter7));
  inv1  gate891(.a(G769), .O(gate264inter8));
  nand2 gate892(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate893(.a(s_49), .b(gate264inter3), .O(gate264inter10));
  nor2  gate894(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate895(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate896(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate2451(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2452(.a(gate266inter0), .b(s_272), .O(gate266inter1));
  and2  gate2453(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2454(.a(s_272), .O(gate266inter3));
  inv1  gate2455(.a(s_273), .O(gate266inter4));
  nand2 gate2456(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2457(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2458(.a(G645), .O(gate266inter7));
  inv1  gate2459(.a(G773), .O(gate266inter8));
  nand2 gate2460(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2461(.a(s_273), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2462(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2463(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2464(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1765(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1766(.a(gate268inter0), .b(s_174), .O(gate268inter1));
  and2  gate1767(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1768(.a(s_174), .O(gate268inter3));
  inv1  gate1769(.a(s_175), .O(gate268inter4));
  nand2 gate1770(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1771(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1772(.a(G651), .O(gate268inter7));
  inv1  gate1773(.a(G779), .O(gate268inter8));
  nand2 gate1774(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1775(.a(s_175), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1776(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1777(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1778(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate953(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate954(.a(gate275inter0), .b(s_58), .O(gate275inter1));
  and2  gate955(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate956(.a(s_58), .O(gate275inter3));
  inv1  gate957(.a(s_59), .O(gate275inter4));
  nand2 gate958(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate959(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate960(.a(G645), .O(gate275inter7));
  inv1  gate961(.a(G797), .O(gate275inter8));
  nand2 gate962(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate963(.a(s_59), .b(gate275inter3), .O(gate275inter10));
  nor2  gate964(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate965(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate966(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2465(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2466(.a(gate279inter0), .b(s_274), .O(gate279inter1));
  and2  gate2467(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2468(.a(s_274), .O(gate279inter3));
  inv1  gate2469(.a(s_275), .O(gate279inter4));
  nand2 gate2470(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2471(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2472(.a(G651), .O(gate279inter7));
  inv1  gate2473(.a(G803), .O(gate279inter8));
  nand2 gate2474(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2475(.a(s_275), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2476(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2477(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2478(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1079(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1080(.a(gate281inter0), .b(s_76), .O(gate281inter1));
  and2  gate1081(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1082(.a(s_76), .O(gate281inter3));
  inv1  gate1083(.a(s_77), .O(gate281inter4));
  nand2 gate1084(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1085(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1086(.a(G654), .O(gate281inter7));
  inv1  gate1087(.a(G806), .O(gate281inter8));
  nand2 gate1088(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1089(.a(s_77), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1090(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1091(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1092(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1737(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1738(.a(gate282inter0), .b(s_170), .O(gate282inter1));
  and2  gate1739(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1740(.a(s_170), .O(gate282inter3));
  inv1  gate1741(.a(s_171), .O(gate282inter4));
  nand2 gate1742(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1743(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1744(.a(G782), .O(gate282inter7));
  inv1  gate1745(.a(G806), .O(gate282inter8));
  nand2 gate1746(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1747(.a(s_171), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1748(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1749(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1750(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2563(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2564(.a(gate283inter0), .b(s_288), .O(gate283inter1));
  and2  gate2565(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2566(.a(s_288), .O(gate283inter3));
  inv1  gate2567(.a(s_289), .O(gate283inter4));
  nand2 gate2568(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2569(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2570(.a(G657), .O(gate283inter7));
  inv1  gate2571(.a(G809), .O(gate283inter8));
  nand2 gate2572(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2573(.a(s_289), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2574(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2575(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2576(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1779(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1780(.a(gate284inter0), .b(s_176), .O(gate284inter1));
  and2  gate1781(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1782(.a(s_176), .O(gate284inter3));
  inv1  gate1783(.a(s_177), .O(gate284inter4));
  nand2 gate1784(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1785(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1786(.a(G785), .O(gate284inter7));
  inv1  gate1787(.a(G809), .O(gate284inter8));
  nand2 gate1788(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1789(.a(s_177), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1790(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1791(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1792(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate771(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate772(.a(gate285inter0), .b(s_32), .O(gate285inter1));
  and2  gate773(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate774(.a(s_32), .O(gate285inter3));
  inv1  gate775(.a(s_33), .O(gate285inter4));
  nand2 gate776(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate777(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate778(.a(G660), .O(gate285inter7));
  inv1  gate779(.a(G812), .O(gate285inter8));
  nand2 gate780(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate781(.a(s_33), .b(gate285inter3), .O(gate285inter10));
  nor2  gate782(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate783(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate784(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1051(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1052(.a(gate287inter0), .b(s_72), .O(gate287inter1));
  and2  gate1053(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1054(.a(s_72), .O(gate287inter3));
  inv1  gate1055(.a(s_73), .O(gate287inter4));
  nand2 gate1056(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1057(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1058(.a(G663), .O(gate287inter7));
  inv1  gate1059(.a(G815), .O(gate287inter8));
  nand2 gate1060(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1061(.a(s_73), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1062(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1063(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1064(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1513(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1514(.a(gate288inter0), .b(s_138), .O(gate288inter1));
  and2  gate1515(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1516(.a(s_138), .O(gate288inter3));
  inv1  gate1517(.a(s_139), .O(gate288inter4));
  nand2 gate1518(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1519(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1520(.a(G791), .O(gate288inter7));
  inv1  gate1521(.a(G815), .O(gate288inter8));
  nand2 gate1522(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1523(.a(s_139), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1524(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1525(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1526(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1821(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1822(.a(gate292inter0), .b(s_182), .O(gate292inter1));
  and2  gate1823(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1824(.a(s_182), .O(gate292inter3));
  inv1  gate1825(.a(s_183), .O(gate292inter4));
  nand2 gate1826(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1827(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1828(.a(G824), .O(gate292inter7));
  inv1  gate1829(.a(G825), .O(gate292inter8));
  nand2 gate1830(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1831(.a(s_183), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1832(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1833(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1834(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2395(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2396(.a(gate294inter0), .b(s_264), .O(gate294inter1));
  and2  gate2397(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2398(.a(s_264), .O(gate294inter3));
  inv1  gate2399(.a(s_265), .O(gate294inter4));
  nand2 gate2400(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2401(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2402(.a(G832), .O(gate294inter7));
  inv1  gate2403(.a(G833), .O(gate294inter8));
  nand2 gate2404(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2405(.a(s_265), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2406(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2407(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2408(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2311(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2312(.a(gate295inter0), .b(s_252), .O(gate295inter1));
  and2  gate2313(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2314(.a(s_252), .O(gate295inter3));
  inv1  gate2315(.a(s_253), .O(gate295inter4));
  nand2 gate2316(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2317(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2318(.a(G830), .O(gate295inter7));
  inv1  gate2319(.a(G831), .O(gate295inter8));
  nand2 gate2320(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2321(.a(s_253), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2322(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2323(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2324(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2661(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2662(.a(gate391inter0), .b(s_302), .O(gate391inter1));
  and2  gate2663(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2664(.a(s_302), .O(gate391inter3));
  inv1  gate2665(.a(s_303), .O(gate391inter4));
  nand2 gate2666(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2667(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2668(.a(G5), .O(gate391inter7));
  inv1  gate2669(.a(G1048), .O(gate391inter8));
  nand2 gate2670(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2671(.a(s_303), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2672(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2673(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2674(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate757(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate758(.a(gate394inter0), .b(s_30), .O(gate394inter1));
  and2  gate759(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate760(.a(s_30), .O(gate394inter3));
  inv1  gate761(.a(s_31), .O(gate394inter4));
  nand2 gate762(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate763(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate764(.a(G8), .O(gate394inter7));
  inv1  gate765(.a(G1057), .O(gate394inter8));
  nand2 gate766(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate767(.a(s_31), .b(gate394inter3), .O(gate394inter10));
  nor2  gate768(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate769(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate770(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1611(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1612(.a(gate395inter0), .b(s_152), .O(gate395inter1));
  and2  gate1613(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1614(.a(s_152), .O(gate395inter3));
  inv1  gate1615(.a(s_153), .O(gate395inter4));
  nand2 gate1616(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1617(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1618(.a(G9), .O(gate395inter7));
  inv1  gate1619(.a(G1060), .O(gate395inter8));
  nand2 gate1620(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1621(.a(s_153), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1622(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1623(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1624(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate561(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate562(.a(gate396inter0), .b(s_2), .O(gate396inter1));
  and2  gate563(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate564(.a(s_2), .O(gate396inter3));
  inv1  gate565(.a(s_3), .O(gate396inter4));
  nand2 gate566(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate567(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate568(.a(G10), .O(gate396inter7));
  inv1  gate569(.a(G1063), .O(gate396inter8));
  nand2 gate570(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate571(.a(s_3), .b(gate396inter3), .O(gate396inter10));
  nor2  gate572(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate573(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate574(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate967(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate968(.a(gate401inter0), .b(s_60), .O(gate401inter1));
  and2  gate969(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate970(.a(s_60), .O(gate401inter3));
  inv1  gate971(.a(s_61), .O(gate401inter4));
  nand2 gate972(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate973(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate974(.a(G15), .O(gate401inter7));
  inv1  gate975(.a(G1078), .O(gate401inter8));
  nand2 gate976(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate977(.a(s_61), .b(gate401inter3), .O(gate401inter10));
  nor2  gate978(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate979(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate980(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1723(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1724(.a(gate402inter0), .b(s_168), .O(gate402inter1));
  and2  gate1725(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1726(.a(s_168), .O(gate402inter3));
  inv1  gate1727(.a(s_169), .O(gate402inter4));
  nand2 gate1728(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1729(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1730(.a(G16), .O(gate402inter7));
  inv1  gate1731(.a(G1081), .O(gate402inter8));
  nand2 gate1732(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1733(.a(s_169), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1734(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1735(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1736(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1695(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1696(.a(gate404inter0), .b(s_164), .O(gate404inter1));
  and2  gate1697(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1698(.a(s_164), .O(gate404inter3));
  inv1  gate1699(.a(s_165), .O(gate404inter4));
  nand2 gate1700(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1701(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1702(.a(G18), .O(gate404inter7));
  inv1  gate1703(.a(G1087), .O(gate404inter8));
  nand2 gate1704(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1705(.a(s_165), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1706(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1707(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1708(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1583(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1584(.a(gate410inter0), .b(s_148), .O(gate410inter1));
  and2  gate1585(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1586(.a(s_148), .O(gate410inter3));
  inv1  gate1587(.a(s_149), .O(gate410inter4));
  nand2 gate1588(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1589(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1590(.a(G24), .O(gate410inter7));
  inv1  gate1591(.a(G1105), .O(gate410inter8));
  nand2 gate1592(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1593(.a(s_149), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1594(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1595(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1596(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1275(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1276(.a(gate413inter0), .b(s_104), .O(gate413inter1));
  and2  gate1277(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1278(.a(s_104), .O(gate413inter3));
  inv1  gate1279(.a(s_105), .O(gate413inter4));
  nand2 gate1280(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1281(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1282(.a(G27), .O(gate413inter7));
  inv1  gate1283(.a(G1114), .O(gate413inter8));
  nand2 gate1284(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1285(.a(s_105), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1286(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1287(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1288(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1107(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1108(.a(gate414inter0), .b(s_80), .O(gate414inter1));
  and2  gate1109(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1110(.a(s_80), .O(gate414inter3));
  inv1  gate1111(.a(s_81), .O(gate414inter4));
  nand2 gate1112(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1113(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1114(.a(G28), .O(gate414inter7));
  inv1  gate1115(.a(G1117), .O(gate414inter8));
  nand2 gate1116(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1117(.a(s_81), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1118(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1119(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1120(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1989(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1990(.a(gate416inter0), .b(s_206), .O(gate416inter1));
  and2  gate1991(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1992(.a(s_206), .O(gate416inter3));
  inv1  gate1993(.a(s_207), .O(gate416inter4));
  nand2 gate1994(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1995(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1996(.a(G30), .O(gate416inter7));
  inv1  gate1997(.a(G1123), .O(gate416inter8));
  nand2 gate1998(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1999(.a(s_207), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2000(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2001(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2002(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1639(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1640(.a(gate417inter0), .b(s_156), .O(gate417inter1));
  and2  gate1641(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1642(.a(s_156), .O(gate417inter3));
  inv1  gate1643(.a(s_157), .O(gate417inter4));
  nand2 gate1644(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1645(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1646(.a(G31), .O(gate417inter7));
  inv1  gate1647(.a(G1126), .O(gate417inter8));
  nand2 gate1648(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1649(.a(s_157), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1650(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1651(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1652(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2409(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2410(.a(gate420inter0), .b(s_266), .O(gate420inter1));
  and2  gate2411(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2412(.a(s_266), .O(gate420inter3));
  inv1  gate2413(.a(s_267), .O(gate420inter4));
  nand2 gate2414(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2415(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2416(.a(G1036), .O(gate420inter7));
  inv1  gate2417(.a(G1132), .O(gate420inter8));
  nand2 gate2418(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2419(.a(s_267), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2420(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2421(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2422(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2507(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2508(.a(gate421inter0), .b(s_280), .O(gate421inter1));
  and2  gate2509(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2510(.a(s_280), .O(gate421inter3));
  inv1  gate2511(.a(s_281), .O(gate421inter4));
  nand2 gate2512(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2513(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2514(.a(G2), .O(gate421inter7));
  inv1  gate2515(.a(G1135), .O(gate421inter8));
  nand2 gate2516(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2517(.a(s_281), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2518(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2519(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2520(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate743(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate744(.a(gate423inter0), .b(s_28), .O(gate423inter1));
  and2  gate745(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate746(.a(s_28), .O(gate423inter3));
  inv1  gate747(.a(s_29), .O(gate423inter4));
  nand2 gate748(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate749(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate750(.a(G3), .O(gate423inter7));
  inv1  gate751(.a(G1138), .O(gate423inter8));
  nand2 gate752(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate753(.a(s_29), .b(gate423inter3), .O(gate423inter10));
  nor2  gate754(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate755(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate756(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2129(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2130(.a(gate424inter0), .b(s_226), .O(gate424inter1));
  and2  gate2131(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2132(.a(s_226), .O(gate424inter3));
  inv1  gate2133(.a(s_227), .O(gate424inter4));
  nand2 gate2134(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2135(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2136(.a(G1042), .O(gate424inter7));
  inv1  gate2137(.a(G1138), .O(gate424inter8));
  nand2 gate2138(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2139(.a(s_227), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2140(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2141(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2142(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1233(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1234(.a(gate426inter0), .b(s_98), .O(gate426inter1));
  and2  gate1235(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1236(.a(s_98), .O(gate426inter3));
  inv1  gate1237(.a(s_99), .O(gate426inter4));
  nand2 gate1238(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1239(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1240(.a(G1045), .O(gate426inter7));
  inv1  gate1241(.a(G1141), .O(gate426inter8));
  nand2 gate1242(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1243(.a(s_99), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1244(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1245(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1246(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate827(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate828(.a(gate428inter0), .b(s_40), .O(gate428inter1));
  and2  gate829(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate830(.a(s_40), .O(gate428inter3));
  inv1  gate831(.a(s_41), .O(gate428inter4));
  nand2 gate832(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate833(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate834(.a(G1048), .O(gate428inter7));
  inv1  gate835(.a(G1144), .O(gate428inter8));
  nand2 gate836(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate837(.a(s_41), .b(gate428inter3), .O(gate428inter10));
  nor2  gate838(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate839(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate840(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1499(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1500(.a(gate435inter0), .b(s_136), .O(gate435inter1));
  and2  gate1501(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1502(.a(s_136), .O(gate435inter3));
  inv1  gate1503(.a(s_137), .O(gate435inter4));
  nand2 gate1504(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1505(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1506(.a(G9), .O(gate435inter7));
  inv1  gate1507(.a(G1156), .O(gate435inter8));
  nand2 gate1508(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1509(.a(s_137), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1510(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1511(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1512(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1471(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1472(.a(gate437inter0), .b(s_132), .O(gate437inter1));
  and2  gate1473(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1474(.a(s_132), .O(gate437inter3));
  inv1  gate1475(.a(s_133), .O(gate437inter4));
  nand2 gate1476(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1477(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1478(.a(G10), .O(gate437inter7));
  inv1  gate1479(.a(G1159), .O(gate437inter8));
  nand2 gate1480(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1481(.a(s_133), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1482(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1483(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1484(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2549(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2550(.a(gate439inter0), .b(s_286), .O(gate439inter1));
  and2  gate2551(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2552(.a(s_286), .O(gate439inter3));
  inv1  gate2553(.a(s_287), .O(gate439inter4));
  nand2 gate2554(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2555(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2556(.a(G11), .O(gate439inter7));
  inv1  gate2557(.a(G1162), .O(gate439inter8));
  nand2 gate2558(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2559(.a(s_287), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2560(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2561(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2562(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1807(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1808(.a(gate442inter0), .b(s_180), .O(gate442inter1));
  and2  gate1809(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1810(.a(s_180), .O(gate442inter3));
  inv1  gate1811(.a(s_181), .O(gate442inter4));
  nand2 gate1812(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1813(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1814(.a(G1069), .O(gate442inter7));
  inv1  gate1815(.a(G1165), .O(gate442inter8));
  nand2 gate1816(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1817(.a(s_181), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1818(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1819(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1820(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1009(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1010(.a(gate444inter0), .b(s_66), .O(gate444inter1));
  and2  gate1011(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1012(.a(s_66), .O(gate444inter3));
  inv1  gate1013(.a(s_67), .O(gate444inter4));
  nand2 gate1014(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1015(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1016(.a(G1072), .O(gate444inter7));
  inv1  gate1017(.a(G1168), .O(gate444inter8));
  nand2 gate1018(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1019(.a(s_67), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1020(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1021(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1022(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1205(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1206(.a(gate445inter0), .b(s_94), .O(gate445inter1));
  and2  gate1207(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1208(.a(s_94), .O(gate445inter3));
  inv1  gate1209(.a(s_95), .O(gate445inter4));
  nand2 gate1210(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1211(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1212(.a(G14), .O(gate445inter7));
  inv1  gate1213(.a(G1171), .O(gate445inter8));
  nand2 gate1214(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1215(.a(s_95), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1216(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1217(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1218(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate813(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate814(.a(gate447inter0), .b(s_38), .O(gate447inter1));
  and2  gate815(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate816(.a(s_38), .O(gate447inter3));
  inv1  gate817(.a(s_39), .O(gate447inter4));
  nand2 gate818(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate819(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate820(.a(G15), .O(gate447inter7));
  inv1  gate821(.a(G1174), .O(gate447inter8));
  nand2 gate822(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate823(.a(s_39), .b(gate447inter3), .O(gate447inter10));
  nor2  gate824(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate825(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate826(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate785(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate786(.a(gate450inter0), .b(s_34), .O(gate450inter1));
  and2  gate787(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate788(.a(s_34), .O(gate450inter3));
  inv1  gate789(.a(s_35), .O(gate450inter4));
  nand2 gate790(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate791(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate792(.a(G1081), .O(gate450inter7));
  inv1  gate793(.a(G1177), .O(gate450inter8));
  nand2 gate794(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate795(.a(s_35), .b(gate450inter3), .O(gate450inter10));
  nor2  gate796(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate797(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate798(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2339(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2340(.a(gate451inter0), .b(s_256), .O(gate451inter1));
  and2  gate2341(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2342(.a(s_256), .O(gate451inter3));
  inv1  gate2343(.a(s_257), .O(gate451inter4));
  nand2 gate2344(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2345(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2346(.a(G17), .O(gate451inter7));
  inv1  gate2347(.a(G1180), .O(gate451inter8));
  nand2 gate2348(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2349(.a(s_257), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2350(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2351(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2352(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1961(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1962(.a(gate452inter0), .b(s_202), .O(gate452inter1));
  and2  gate1963(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1964(.a(s_202), .O(gate452inter3));
  inv1  gate1965(.a(s_203), .O(gate452inter4));
  nand2 gate1966(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1967(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1968(.a(G1084), .O(gate452inter7));
  inv1  gate1969(.a(G1180), .O(gate452inter8));
  nand2 gate1970(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1971(.a(s_203), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1972(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1973(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1974(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate1485(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1486(.a(gate453inter0), .b(s_134), .O(gate453inter1));
  and2  gate1487(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1488(.a(s_134), .O(gate453inter3));
  inv1  gate1489(.a(s_135), .O(gate453inter4));
  nand2 gate1490(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1491(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1492(.a(G18), .O(gate453inter7));
  inv1  gate1493(.a(G1183), .O(gate453inter8));
  nand2 gate1494(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1495(.a(s_135), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1496(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1497(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1498(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1625(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1626(.a(gate455inter0), .b(s_154), .O(gate455inter1));
  and2  gate1627(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1628(.a(s_154), .O(gate455inter3));
  inv1  gate1629(.a(s_155), .O(gate455inter4));
  nand2 gate1630(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1631(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1632(.a(G19), .O(gate455inter7));
  inv1  gate1633(.a(G1186), .O(gate455inter8));
  nand2 gate1634(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1635(.a(s_155), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1636(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1637(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1638(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate2171(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2172(.a(gate456inter0), .b(s_232), .O(gate456inter1));
  and2  gate2173(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2174(.a(s_232), .O(gate456inter3));
  inv1  gate2175(.a(s_233), .O(gate456inter4));
  nand2 gate2176(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2177(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2178(.a(G1090), .O(gate456inter7));
  inv1  gate2179(.a(G1186), .O(gate456inter8));
  nand2 gate2180(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2181(.a(s_233), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2182(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2183(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2184(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1093(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1094(.a(gate461inter0), .b(s_78), .O(gate461inter1));
  and2  gate1095(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1096(.a(s_78), .O(gate461inter3));
  inv1  gate1097(.a(s_79), .O(gate461inter4));
  nand2 gate1098(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1099(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1100(.a(G22), .O(gate461inter7));
  inv1  gate1101(.a(G1195), .O(gate461inter8));
  nand2 gate1102(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1103(.a(s_79), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1104(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1105(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1106(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1037(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1038(.a(gate463inter0), .b(s_70), .O(gate463inter1));
  and2  gate1039(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1040(.a(s_70), .O(gate463inter3));
  inv1  gate1041(.a(s_71), .O(gate463inter4));
  nand2 gate1042(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1043(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1044(.a(G23), .O(gate463inter7));
  inv1  gate1045(.a(G1198), .O(gate463inter8));
  nand2 gate1046(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1047(.a(s_71), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1048(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1049(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1050(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate715(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate716(.a(gate472inter0), .b(s_24), .O(gate472inter1));
  and2  gate717(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate718(.a(s_24), .O(gate472inter3));
  inv1  gate719(.a(s_25), .O(gate472inter4));
  nand2 gate720(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate721(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate722(.a(G1114), .O(gate472inter7));
  inv1  gate723(.a(G1210), .O(gate472inter8));
  nand2 gate724(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate725(.a(s_25), .b(gate472inter3), .O(gate472inter10));
  nor2  gate726(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate727(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate728(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate939(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate940(.a(gate473inter0), .b(s_56), .O(gate473inter1));
  and2  gate941(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate942(.a(s_56), .O(gate473inter3));
  inv1  gate943(.a(s_57), .O(gate473inter4));
  nand2 gate944(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate945(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate946(.a(G28), .O(gate473inter7));
  inv1  gate947(.a(G1213), .O(gate473inter8));
  nand2 gate948(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate949(.a(s_57), .b(gate473inter3), .O(gate473inter10));
  nor2  gate950(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate951(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate952(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1023(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1024(.a(gate481inter0), .b(s_68), .O(gate481inter1));
  and2  gate1025(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1026(.a(s_68), .O(gate481inter3));
  inv1  gate1027(.a(s_69), .O(gate481inter4));
  nand2 gate1028(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1029(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1030(.a(G32), .O(gate481inter7));
  inv1  gate1031(.a(G1225), .O(gate481inter8));
  nand2 gate1032(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1033(.a(s_69), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1034(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1035(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1036(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1191(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1192(.a(gate485inter0), .b(s_92), .O(gate485inter1));
  and2  gate1193(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1194(.a(s_92), .O(gate485inter3));
  inv1  gate1195(.a(s_93), .O(gate485inter4));
  nand2 gate1196(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1197(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1198(.a(G1232), .O(gate485inter7));
  inv1  gate1199(.a(G1233), .O(gate485inter8));
  nand2 gate1200(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1201(.a(s_93), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1202(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1203(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1204(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2115(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2116(.a(gate489inter0), .b(s_224), .O(gate489inter1));
  and2  gate2117(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2118(.a(s_224), .O(gate489inter3));
  inv1  gate2119(.a(s_225), .O(gate489inter4));
  nand2 gate2120(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2121(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2122(.a(G1240), .O(gate489inter7));
  inv1  gate2123(.a(G1241), .O(gate489inter8));
  nand2 gate2124(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2125(.a(s_225), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2126(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2127(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2128(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1121(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1122(.a(gate490inter0), .b(s_82), .O(gate490inter1));
  and2  gate1123(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1124(.a(s_82), .O(gate490inter3));
  inv1  gate1125(.a(s_83), .O(gate490inter4));
  nand2 gate1126(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1127(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1128(.a(G1242), .O(gate490inter7));
  inv1  gate1129(.a(G1243), .O(gate490inter8));
  nand2 gate1130(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1131(.a(s_83), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1132(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1133(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1134(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2045(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2046(.a(gate493inter0), .b(s_214), .O(gate493inter1));
  and2  gate2047(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2048(.a(s_214), .O(gate493inter3));
  inv1  gate2049(.a(s_215), .O(gate493inter4));
  nand2 gate2050(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2051(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2052(.a(G1248), .O(gate493inter7));
  inv1  gate2053(.a(G1249), .O(gate493inter8));
  nand2 gate2054(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2055(.a(s_215), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2056(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2057(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2058(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2605(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2606(.a(gate497inter0), .b(s_294), .O(gate497inter1));
  and2  gate2607(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2608(.a(s_294), .O(gate497inter3));
  inv1  gate2609(.a(s_295), .O(gate497inter4));
  nand2 gate2610(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2611(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2612(.a(G1256), .O(gate497inter7));
  inv1  gate2613(.a(G1257), .O(gate497inter8));
  nand2 gate2614(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2615(.a(s_295), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2616(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2617(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2618(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1653(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1654(.a(gate498inter0), .b(s_158), .O(gate498inter1));
  and2  gate1655(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1656(.a(s_158), .O(gate498inter3));
  inv1  gate1657(.a(s_159), .O(gate498inter4));
  nand2 gate1658(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1659(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1660(.a(G1258), .O(gate498inter7));
  inv1  gate1661(.a(G1259), .O(gate498inter8));
  nand2 gate1662(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1663(.a(s_159), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1664(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1665(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1666(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2101(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2102(.a(gate500inter0), .b(s_222), .O(gate500inter1));
  and2  gate2103(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2104(.a(s_222), .O(gate500inter3));
  inv1  gate2105(.a(s_223), .O(gate500inter4));
  nand2 gate2106(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2107(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2108(.a(G1262), .O(gate500inter7));
  inv1  gate2109(.a(G1263), .O(gate500inter8));
  nand2 gate2110(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2111(.a(s_223), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2112(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2113(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2114(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2255(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2256(.a(gate507inter0), .b(s_244), .O(gate507inter1));
  and2  gate2257(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2258(.a(s_244), .O(gate507inter3));
  inv1  gate2259(.a(s_245), .O(gate507inter4));
  nand2 gate2260(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2261(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2262(.a(G1276), .O(gate507inter7));
  inv1  gate2263(.a(G1277), .O(gate507inter8));
  nand2 gate2264(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2265(.a(s_245), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2266(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2267(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2268(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate701(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate702(.a(gate508inter0), .b(s_22), .O(gate508inter1));
  and2  gate703(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate704(.a(s_22), .O(gate508inter3));
  inv1  gate705(.a(s_23), .O(gate508inter4));
  nand2 gate706(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate707(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate708(.a(G1278), .O(gate508inter7));
  inv1  gate709(.a(G1279), .O(gate508inter8));
  nand2 gate710(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate711(.a(s_23), .b(gate508inter3), .O(gate508inter10));
  nor2  gate712(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate713(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate714(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule