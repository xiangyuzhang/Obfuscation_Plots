module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;
wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate303inter0, gate303inter1, gate303inter2, gate303inter3, gate303inter4, gate303inter5, gate303inter6, gate303inter7, gate303inter8, gate303inter9, gate303inter10, gate303inter11, gate303inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate346inter0, gate346inter1, gate346inter2, gate346inter3, gate346inter4, gate346inter5, gate346inter6, gate346inter7, gate346inter8, gate346inter9, gate346inter10, gate346inter11, gate346inter12, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate327inter0, gate327inter1, gate327inter2, gate327inter3, gate327inter4, gate327inter5, gate327inter6, gate327inter7, gate327inter8, gate327inter9, gate327inter10, gate327inter11, gate327inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate307inter0, gate307inter1, gate307inter2, gate307inter3, gate307inter4, gate307inter5, gate307inter6, gate307inter7, gate307inter8, gate307inter9, gate307inter10, gate307inter11, gate307inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate311inter0, gate311inter1, gate311inter2, gate311inter3, gate311inter4, gate311inter5, gate311inter6, gate311inter7, gate311inter8, gate311inter9, gate311inter10, gate311inter11, gate311inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate348inter0, gate348inter1, gate348inter2, gate348inter3, gate348inter4, gate348inter5, gate348inter6, gate348inter7, gate348inter8, gate348inter9, gate348inter10, gate348inter11, gate348inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate310inter0, gate310inter1, gate310inter2, gate310inter3, gate310inter4, gate310inter5, gate310inter6, gate310inter7, gate310inter8, gate310inter9, gate310inter10, gate310inter11, gate310inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate330inter0, gate330inter1, gate330inter2, gate330inter3, gate330inter4, gate330inter5, gate330inter6, gate330inter7, gate330inter8, gate330inter9, gate330inter10, gate330inter11, gate330inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate331inter0, gate331inter1, gate331inter2, gate331inter3, gate331inter4, gate331inter5, gate331inter6, gate331inter7, gate331inter8, gate331inter9, gate331inter10, gate331inter11, gate331inter12;


nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );

  xor2  gate818(.a(N96), .b(N91), .O(gate20inter0));
  nand2 gate819(.a(gate20inter0), .b(s_62), .O(gate20inter1));
  and2  gate820(.a(N96), .b(N91), .O(gate20inter2));
  inv1  gate821(.a(s_62), .O(gate20inter3));
  inv1  gate822(.a(s_63), .O(gate20inter4));
  nand2 gate823(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate824(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate825(.a(N91), .O(gate20inter7));
  inv1  gate826(.a(N96), .O(gate20inter8));
  nand2 gate827(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate828(.a(s_63), .b(gate20inter3), .O(gate20inter10));
  nor2  gate829(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate830(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate831(.a(gate20inter12), .b(gate20inter1), .O(N301));
or2 gate21( .a(N91), .b(N96), .O(N302) );

  xor2  gate972(.a(N106), .b(N101), .O(gate22inter0));
  nand2 gate973(.a(gate22inter0), .b(s_84), .O(gate22inter1));
  and2  gate974(.a(N106), .b(N101), .O(gate22inter2));
  inv1  gate975(.a(s_84), .O(gate22inter3));
  inv1  gate976(.a(s_85), .O(gate22inter4));
  nand2 gate977(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate978(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate979(.a(N101), .O(gate22inter7));
  inv1  gate980(.a(N106), .O(gate22inter8));
  nand2 gate981(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate982(.a(s_85), .b(gate22inter3), .O(gate22inter10));
  nor2  gate983(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate984(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate985(.a(gate22inter12), .b(gate22inter1), .O(N303));
or2 gate23( .a(N101), .b(N106), .O(N304) );

  xor2  gate762(.a(N116), .b(N111), .O(gate24inter0));
  nand2 gate763(.a(gate24inter0), .b(s_54), .O(gate24inter1));
  and2  gate764(.a(N116), .b(N111), .O(gate24inter2));
  inv1  gate765(.a(s_54), .O(gate24inter3));
  inv1  gate766(.a(s_55), .O(gate24inter4));
  nand2 gate767(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate768(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate769(.a(N111), .O(gate24inter7));
  inv1  gate770(.a(N116), .O(gate24inter8));
  nand2 gate771(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate772(.a(s_55), .b(gate24inter3), .O(gate24inter10));
  nor2  gate773(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate774(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate775(.a(gate24inter12), .b(gate24inter1), .O(N305));
or2 gate25( .a(N111), .b(N116), .O(N306) );

  xor2  gate1280(.a(N126), .b(N121), .O(gate26inter0));
  nand2 gate1281(.a(gate26inter0), .b(s_128), .O(gate26inter1));
  and2  gate1282(.a(N126), .b(N121), .O(gate26inter2));
  inv1  gate1283(.a(s_128), .O(gate26inter3));
  inv1  gate1284(.a(s_129), .O(gate26inter4));
  nand2 gate1285(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1286(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1287(.a(N121), .O(gate26inter7));
  inv1  gate1288(.a(N126), .O(gate26inter8));
  nand2 gate1289(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1290(.a(s_129), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1291(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1292(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1293(.a(gate26inter12), .b(gate26inter1), .O(N307));
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );

  xor2  gate398(.a(N156), .b(N59), .O(gate33inter0));
  nand2 gate399(.a(gate33inter0), .b(s_2), .O(gate33inter1));
  and2  gate400(.a(N156), .b(N59), .O(gate33inter2));
  inv1  gate401(.a(s_2), .O(gate33inter3));
  inv1  gate402(.a(s_3), .O(gate33inter4));
  nand2 gate403(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate404(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate405(.a(N59), .O(gate33inter7));
  inv1  gate406(.a(N156), .O(gate33inter8));
  nand2 gate407(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate408(.a(s_3), .b(gate33inter3), .O(gate33inter10));
  nor2  gate409(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate410(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate411(.a(gate33inter12), .b(gate33inter1), .O(N319));
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17), .b(N42), .O(N323) );

  xor2  gate734(.a(N165), .b(N159), .O(gate36inter0));
  nand2 gate735(.a(gate36inter0), .b(s_50), .O(gate36inter1));
  and2  gate736(.a(N165), .b(N159), .O(gate36inter2));
  inv1  gate737(.a(s_50), .O(gate36inter3));
  inv1  gate738(.a(s_51), .O(gate36inter4));
  nand2 gate739(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate740(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate741(.a(N159), .O(gate36inter7));
  inv1  gate742(.a(N165), .O(gate36inter8));
  nand2 gate743(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate744(.a(s_51), .b(gate36inter3), .O(gate36inter10));
  nor2  gate745(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate746(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate747(.a(gate36inter12), .b(gate36inter1), .O(N324));
or2 gate37( .a(N159), .b(N165), .O(N325) );

  xor2  gate552(.a(N177), .b(N171), .O(gate38inter0));
  nand2 gate553(.a(gate38inter0), .b(s_24), .O(gate38inter1));
  and2  gate554(.a(N177), .b(N171), .O(gate38inter2));
  inv1  gate555(.a(s_24), .O(gate38inter3));
  inv1  gate556(.a(s_25), .O(gate38inter4));
  nand2 gate557(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate558(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate559(.a(N171), .O(gate38inter7));
  inv1  gate560(.a(N177), .O(gate38inter8));
  nand2 gate561(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate562(.a(s_25), .b(gate38inter3), .O(gate38inter10));
  nor2  gate563(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate564(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate565(.a(gate38inter12), .b(gate38inter1), .O(N326));
or2 gate39( .a(N171), .b(N177), .O(N327) );

  xor2  gate1266(.a(N189), .b(N183), .O(gate40inter0));
  nand2 gate1267(.a(gate40inter0), .b(s_126), .O(gate40inter1));
  and2  gate1268(.a(N189), .b(N183), .O(gate40inter2));
  inv1  gate1269(.a(s_126), .O(gate40inter3));
  inv1  gate1270(.a(s_127), .O(gate40inter4));
  nand2 gate1271(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1272(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1273(.a(N183), .O(gate40inter7));
  inv1  gate1274(.a(N189), .O(gate40inter8));
  nand2 gate1275(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1276(.a(s_127), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1277(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1278(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1279(.a(gate40inter12), .b(gate40inter1), .O(N328));
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
and2 gate49( .a(N255), .b(N259), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );

  xor2  gate748(.a(N284), .b(N280), .O(gate60inter0));
  nand2 gate749(.a(gate60inter0), .b(s_52), .O(gate60inter1));
  and2  gate750(.a(N284), .b(N280), .O(gate60inter2));
  inv1  gate751(.a(s_52), .O(gate60inter3));
  inv1  gate752(.a(s_53), .O(gate60inter4));
  nand2 gate753(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate754(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate755(.a(N280), .O(gate60inter7));
  inv1  gate756(.a(N284), .O(gate60inter8));
  nand2 gate757(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate758(.a(s_53), .b(gate60inter3), .O(gate60inter10));
  nor2  gate759(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate760(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate761(.a(gate60inter12), .b(gate60inter1), .O(N348));
or2 gate61( .a(N280), .b(N285), .O(N349) );
or2 gate62( .a(N280), .b(N286), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );
nand2 gate67( .a(N89), .b(N298), .O(N355) );
and2 gate68( .a(N90), .b(N298), .O(N356) );

  xor2  gate804(.a(N302), .b(N301), .O(gate69inter0));
  nand2 gate805(.a(gate69inter0), .b(s_60), .O(gate69inter1));
  and2  gate806(.a(N302), .b(N301), .O(gate69inter2));
  inv1  gate807(.a(s_60), .O(gate69inter3));
  inv1  gate808(.a(s_61), .O(gate69inter4));
  nand2 gate809(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate810(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate811(.a(N301), .O(gate69inter7));
  inv1  gate812(.a(N302), .O(gate69inter8));
  nand2 gate813(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate814(.a(s_61), .b(gate69inter3), .O(gate69inter10));
  nor2  gate815(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate816(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate817(.a(gate69inter12), .b(gate69inter1), .O(N357));

  xor2  gate1238(.a(N304), .b(N303), .O(gate70inter0));
  nand2 gate1239(.a(gate70inter0), .b(s_122), .O(gate70inter1));
  and2  gate1240(.a(N304), .b(N303), .O(gate70inter2));
  inv1  gate1241(.a(s_122), .O(gate70inter3));
  inv1  gate1242(.a(s_123), .O(gate70inter4));
  nand2 gate1243(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1244(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1245(.a(N303), .O(gate70inter7));
  inv1  gate1246(.a(N304), .O(gate70inter8));
  nand2 gate1247(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1248(.a(s_123), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1249(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1250(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1251(.a(gate70inter12), .b(gate70inter1), .O(N360));

  xor2  gate1294(.a(N306), .b(N305), .O(gate71inter0));
  nand2 gate1295(.a(gate71inter0), .b(s_130), .O(gate71inter1));
  and2  gate1296(.a(N306), .b(N305), .O(gate71inter2));
  inv1  gate1297(.a(s_130), .O(gate71inter3));
  inv1  gate1298(.a(s_131), .O(gate71inter4));
  nand2 gate1299(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1300(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1301(.a(N305), .O(gate71inter7));
  inv1  gate1302(.a(N306), .O(gate71inter8));
  nand2 gate1303(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1304(.a(s_131), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1305(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1306(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1307(.a(gate71inter12), .b(gate71inter1), .O(N363));

  xor2  gate664(.a(N308), .b(N307), .O(gate72inter0));
  nand2 gate665(.a(gate72inter0), .b(s_40), .O(gate72inter1));
  and2  gate666(.a(N308), .b(N307), .O(gate72inter2));
  inv1  gate667(.a(s_40), .O(gate72inter3));
  inv1  gate668(.a(s_41), .O(gate72inter4));
  nand2 gate669(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate670(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate671(.a(N307), .O(gate72inter7));
  inv1  gate672(.a(N308), .O(gate72inter8));
  nand2 gate673(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate674(.a(s_41), .b(gate72inter3), .O(gate72inter10));
  nor2  gate675(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate676(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate677(.a(gate72inter12), .b(gate72inter1), .O(N366));
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );

  xor2  gate538(.a(N327), .b(N326), .O(gate76inter0));
  nand2 gate539(.a(gate76inter0), .b(s_22), .O(gate76inter1));
  and2  gate540(.a(N327), .b(N326), .O(gate76inter2));
  inv1  gate541(.a(s_22), .O(gate76inter3));
  inv1  gate542(.a(s_23), .O(gate76inter4));
  nand2 gate543(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate544(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate545(.a(N326), .O(gate76inter7));
  inv1  gate546(.a(N327), .O(gate76inter8));
  nand2 gate547(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate548(.a(s_23), .b(gate76inter3), .O(gate76inter10));
  nor2  gate549(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate550(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate551(.a(gate76inter12), .b(gate76inter1), .O(N379));
nand2 gate77( .a(N328), .b(N329), .O(N382) );
nand2 gate78( .a(N330), .b(N331), .O(N385) );
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );

  xor2  gate1154(.a(N352), .b(N347), .O(gate96inter0));
  nand2 gate1155(.a(gate96inter0), .b(s_110), .O(gate96inter1));
  and2  gate1156(.a(N352), .b(N347), .O(gate96inter2));
  inv1  gate1157(.a(s_110), .O(gate96inter3));
  inv1  gate1158(.a(s_111), .O(gate96inter4));
  nand2 gate1159(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1160(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1161(.a(N347), .O(gate96inter7));
  inv1  gate1162(.a(N352), .O(gate96inter8));
  nand2 gate1163(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1164(.a(s_111), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1165(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1166(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1167(.a(gate96inter12), .b(gate96inter1), .O(N410));
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );
nor2 gate126( .a(N406), .b(N425), .O(N460) );

  xor2  gate384(.a(N426), .b(N409), .O(gate127inter0));
  nand2 gate385(.a(gate127inter0), .b(s_0), .O(gate127inter1));
  and2  gate386(.a(N426), .b(N409), .O(gate127inter2));
  inv1  gate387(.a(s_0), .O(gate127inter3));
  inv1  gate388(.a(s_1), .O(gate127inter4));
  nand2 gate389(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate390(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate391(.a(N409), .O(gate127inter7));
  inv1  gate392(.a(N426), .O(gate127inter8));
  nand2 gate393(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate394(.a(s_1), .b(gate127inter3), .O(gate127inter10));
  nor2  gate395(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate396(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate397(.a(gate127inter12), .b(gate127inter1), .O(N463));

  xor2  gate622(.a(N410), .b(N442), .O(gate128inter0));
  nand2 gate623(.a(gate128inter0), .b(s_34), .O(gate128inter1));
  and2  gate624(.a(N410), .b(N442), .O(gate128inter2));
  inv1  gate625(.a(s_34), .O(gate128inter3));
  inv1  gate626(.a(s_35), .O(gate128inter4));
  nand2 gate627(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate628(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate629(.a(N442), .O(gate128inter7));
  inv1  gate630(.a(N410), .O(gate128inter8));
  nand2 gate631(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate632(.a(s_35), .b(gate128inter3), .O(gate128inter10));
  nor2  gate633(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate634(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate635(.a(gate128inter12), .b(gate128inter1), .O(N466));
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );

  xor2  gate944(.a(N1), .b(N443), .O(gate137inter0));
  nand2 gate945(.a(gate137inter0), .b(s_80), .O(gate137inter1));
  and2  gate946(.a(N1), .b(N443), .O(gate137inter2));
  inv1  gate947(.a(s_80), .O(gate137inter3));
  inv1  gate948(.a(s_81), .O(gate137inter4));
  nand2 gate949(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate950(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate951(.a(N443), .O(gate137inter7));
  inv1  gate952(.a(N1), .O(gate137inter8));
  nand2 gate953(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate954(.a(s_81), .b(gate137inter3), .O(gate137inter10));
  nor2  gate955(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate956(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate957(.a(gate137inter12), .b(gate137inter1), .O(N483));
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );

  xor2  gate1308(.a(N444), .b(N413), .O(gate142inter0));
  nand2 gate1309(.a(gate142inter0), .b(s_132), .O(gate142inter1));
  and2  gate1310(.a(N444), .b(N413), .O(gate142inter2));
  inv1  gate1311(.a(s_132), .O(gate142inter3));
  inv1  gate1312(.a(s_133), .O(gate142inter4));
  nand2 gate1313(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1314(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1315(.a(N413), .O(gate142inter7));
  inv1  gate1316(.a(N444), .O(gate142inter8));
  nand2 gate1317(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1318(.a(s_133), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1319(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1320(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1321(.a(gate142inter12), .b(gate142inter1), .O(N492));
nor2 gate143( .a(N416), .b(N445), .O(N495) );

  xor2  gate636(.a(N460), .b(N130), .O(gate144inter0));
  nand2 gate637(.a(gate144inter0), .b(s_36), .O(gate144inter1));
  and2  gate638(.a(N460), .b(N130), .O(gate144inter2));
  inv1  gate639(.a(s_36), .O(gate144inter3));
  inv1  gate640(.a(s_37), .O(gate144inter4));
  nand2 gate641(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate642(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate643(.a(N130), .O(gate144inter7));
  inv1  gate644(.a(N460), .O(gate144inter8));
  nand2 gate645(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate646(.a(s_37), .b(gate144inter3), .O(gate144inter10));
  nor2  gate647(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate648(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate649(.a(gate144inter12), .b(gate144inter1), .O(N498));
or2 gate145( .a(N130), .b(N460), .O(N499) );

  xor2  gate916(.a(N135), .b(N463), .O(gate146inter0));
  nand2 gate917(.a(gate146inter0), .b(s_76), .O(gate146inter1));
  and2  gate918(.a(N135), .b(N463), .O(gate146inter2));
  inv1  gate919(.a(s_76), .O(gate146inter3));
  inv1  gate920(.a(s_77), .O(gate146inter4));
  nand2 gate921(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate922(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate923(.a(N463), .O(gate146inter7));
  inv1  gate924(.a(N135), .O(gate146inter8));
  nand2 gate925(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate926(.a(s_77), .b(gate146inter3), .O(gate146inter10));
  nor2  gate927(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate928(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate929(.a(gate146inter12), .b(gate146inter1), .O(N500));
or2 gate147( .a(N463), .b(N135), .O(N501) );
and2 gate148( .a(N91), .b(N466), .O(N502) );

  xor2  gate930(.a(N476), .b(N475), .O(gate149inter0));
  nand2 gate931(.a(gate149inter0), .b(s_78), .O(gate149inter1));
  and2  gate932(.a(N476), .b(N475), .O(gate149inter2));
  inv1  gate933(.a(s_78), .O(gate149inter3));
  inv1  gate934(.a(s_79), .O(gate149inter4));
  nand2 gate935(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate936(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate937(.a(N475), .O(gate149inter7));
  inv1  gate938(.a(N476), .O(gate149inter8));
  nand2 gate939(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate940(.a(s_79), .b(gate149inter3), .O(gate149inter10));
  nor2  gate941(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate942(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate943(.a(gate149inter12), .b(gate149inter1), .O(N503));
and2 gate150( .a(N96), .b(N466), .O(N504) );
nor2 gate151( .a(N477), .b(N478), .O(N505) );
and2 gate152( .a(N101), .b(N466), .O(N506) );

  xor2  gate1210(.a(N480), .b(N479), .O(gate153inter0));
  nand2 gate1211(.a(gate153inter0), .b(s_118), .O(gate153inter1));
  and2  gate1212(.a(N480), .b(N479), .O(gate153inter2));
  inv1  gate1213(.a(s_118), .O(gate153inter3));
  inv1  gate1214(.a(s_119), .O(gate153inter4));
  nand2 gate1215(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1216(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1217(.a(N479), .O(gate153inter7));
  inv1  gate1218(.a(N480), .O(gate153inter8));
  nand2 gate1219(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1220(.a(s_119), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1221(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1222(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1223(.a(gate153inter12), .b(gate153inter1), .O(N507));
and2 gate154( .a(N106), .b(N466), .O(N508) );

  xor2  gate1378(.a(N482), .b(N481), .O(gate155inter0));
  nand2 gate1379(.a(gate155inter0), .b(s_142), .O(gate155inter1));
  and2  gate1380(.a(N482), .b(N481), .O(gate155inter2));
  inv1  gate1381(.a(s_142), .O(gate155inter3));
  inv1  gate1382(.a(s_143), .O(gate155inter4));
  nand2 gate1383(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1384(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1385(.a(N481), .O(gate155inter7));
  inv1  gate1386(.a(N482), .O(gate155inter8));
  nand2 gate1387(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1388(.a(s_143), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1389(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1390(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1391(.a(gate155inter12), .b(gate155inter1), .O(N509));
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );
nand2 gate164( .a(N130), .b(N492), .O(N518) );
or2 gate165( .a(N130), .b(N492), .O(N519) );
nand2 gate166( .a(N495), .b(N207), .O(N520) );
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
and2 gate170( .a(N451), .b(N171), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );

  xor2  gate790(.a(N189), .b(N451), .O(gate173inter0));
  nand2 gate791(.a(gate173inter0), .b(s_58), .O(gate173inter1));
  and2  gate792(.a(N189), .b(N451), .O(gate173inter2));
  inv1  gate793(.a(s_58), .O(gate173inter3));
  inv1  gate794(.a(s_59), .O(gate173inter4));
  nand2 gate795(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate796(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate797(.a(N451), .O(gate173inter7));
  inv1  gate798(.a(N189), .O(gate173inter8));
  nand2 gate799(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate800(.a(s_59), .b(gate173inter3), .O(gate173inter10));
  nor2  gate801(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate802(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate803(.a(gate173inter12), .b(gate173inter1), .O(N527));

  xor2  gate776(.a(N195), .b(N451), .O(gate174inter0));
  nand2 gate777(.a(gate174inter0), .b(s_56), .O(gate174inter1));
  and2  gate778(.a(N195), .b(N451), .O(gate174inter2));
  inv1  gate779(.a(s_56), .O(gate174inter3));
  inv1  gate780(.a(s_57), .O(gate174inter4));
  nand2 gate781(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate782(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate783(.a(N451), .O(gate174inter7));
  inv1  gate784(.a(N195), .O(gate174inter8));
  nand2 gate785(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate786(.a(s_57), .b(gate174inter3), .O(gate174inter10));
  nor2  gate787(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate788(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate789(.a(gate174inter12), .b(gate174inter1), .O(N528));

  xor2  gate468(.a(N201), .b(N451), .O(gate175inter0));
  nand2 gate469(.a(gate175inter0), .b(s_12), .O(gate175inter1));
  and2  gate470(.a(N201), .b(N451), .O(gate175inter2));
  inv1  gate471(.a(s_12), .O(gate175inter3));
  inv1  gate472(.a(s_13), .O(gate175inter4));
  nand2 gate473(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate474(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate475(.a(N451), .O(gate175inter7));
  inv1  gate476(.a(N201), .O(gate175inter8));
  nand2 gate477(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate478(.a(s_13), .b(gate175inter3), .O(gate175inter10));
  nor2  gate479(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate480(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate481(.a(gate175inter12), .b(gate175inter1), .O(N529));
nand2 gate176( .a(N498), .b(N499), .O(N530) );

  xor2  gate1406(.a(N501), .b(N500), .O(gate177inter0));
  nand2 gate1407(.a(gate177inter0), .b(s_146), .O(gate177inter1));
  and2  gate1408(.a(N501), .b(N500), .O(gate177inter2));
  inv1  gate1409(.a(s_146), .O(gate177inter3));
  inv1  gate1410(.a(s_147), .O(gate177inter4));
  nand2 gate1411(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1412(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1413(.a(N500), .O(gate177inter7));
  inv1  gate1414(.a(N501), .O(gate177inter8));
  nand2 gate1415(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1416(.a(s_147), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1417(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1418(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1419(.a(gate177inter12), .b(gate177inter1), .O(N533));

  xor2  gate454(.a(N502), .b(N309), .O(gate178inter0));
  nand2 gate455(.a(gate178inter0), .b(s_10), .O(gate178inter1));
  and2  gate456(.a(N502), .b(N309), .O(gate178inter2));
  inv1  gate457(.a(s_10), .O(gate178inter3));
  inv1  gate458(.a(s_11), .O(gate178inter4));
  nand2 gate459(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate460(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate461(.a(N309), .O(gate178inter7));
  inv1  gate462(.a(N502), .O(gate178inter8));
  nand2 gate463(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate464(.a(s_11), .b(gate178inter3), .O(gate178inter10));
  nor2  gate465(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate466(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate467(.a(gate178inter12), .b(gate178inter1), .O(N536));
nor2 gate179( .a(N316), .b(N504), .O(N537) );

  xor2  gate678(.a(N506), .b(N317), .O(gate180inter0));
  nand2 gate679(.a(gate180inter0), .b(s_42), .O(gate180inter1));
  and2  gate680(.a(N506), .b(N317), .O(gate180inter2));
  inv1  gate681(.a(s_42), .O(gate180inter3));
  inv1  gate682(.a(s_43), .O(gate180inter4));
  nand2 gate683(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate684(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate685(.a(N317), .O(gate180inter7));
  inv1  gate686(.a(N506), .O(gate180inter8));
  nand2 gate687(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate688(.a(s_43), .b(gate180inter3), .O(gate180inter10));
  nor2  gate689(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate690(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate691(.a(gate180inter12), .b(gate180inter1), .O(N538));
nor2 gate181( .a(N318), .b(N508), .O(N539) );
nor2 gate182( .a(N510), .b(N511), .O(N540) );
nor2 gate183( .a(N512), .b(N513), .O(N541) );

  xor2  gate958(.a(N515), .b(N514), .O(gate184inter0));
  nand2 gate959(.a(gate184inter0), .b(s_82), .O(gate184inter1));
  and2  gate960(.a(N515), .b(N514), .O(gate184inter2));
  inv1  gate961(.a(s_82), .O(gate184inter3));
  inv1  gate962(.a(s_83), .O(gate184inter4));
  nand2 gate963(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate964(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate965(.a(N514), .O(gate184inter7));
  inv1  gate966(.a(N515), .O(gate184inter8));
  nand2 gate967(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate968(.a(s_83), .b(gate184inter3), .O(gate184inter10));
  nor2  gate969(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate970(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate971(.a(gate184inter12), .b(gate184inter1), .O(N542));
nor2 gate185( .a(N516), .b(N517), .O(N543) );
nand2 gate186( .a(N518), .b(N519), .O(N544) );

  xor2  gate1224(.a(N521), .b(N520), .O(gate187inter0));
  nand2 gate1225(.a(gate187inter0), .b(s_120), .O(gate187inter1));
  and2  gate1226(.a(N521), .b(N520), .O(gate187inter2));
  inv1  gate1227(.a(s_120), .O(gate187inter3));
  inv1  gate1228(.a(s_121), .O(gate187inter4));
  nand2 gate1229(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1230(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1231(.a(N520), .O(gate187inter7));
  inv1  gate1232(.a(N521), .O(gate187inter8));
  nand2 gate1233(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1234(.a(s_121), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1235(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1236(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1237(.a(gate187inter12), .b(gate187inter1), .O(N547));
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );

  xor2  gate1420(.a(N503), .b(N536), .O(gate191inter0));
  nand2 gate1421(.a(gate191inter0), .b(s_148), .O(gate191inter1));
  and2  gate1422(.a(N503), .b(N536), .O(gate191inter2));
  inv1  gate1423(.a(s_148), .O(gate191inter3));
  inv1  gate1424(.a(s_149), .O(gate191inter4));
  nand2 gate1425(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1426(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1427(.a(N536), .O(gate191inter7));
  inv1  gate1428(.a(N503), .O(gate191inter8));
  nand2 gate1429(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1430(.a(s_149), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1431(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1432(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1433(.a(gate191inter12), .b(gate191inter1), .O(N553));

  xor2  gate1014(.a(N505), .b(N537), .O(gate192inter0));
  nand2 gate1015(.a(gate192inter0), .b(s_90), .O(gate192inter1));
  and2  gate1016(.a(N505), .b(N537), .O(gate192inter2));
  inv1  gate1017(.a(s_90), .O(gate192inter3));
  inv1  gate1018(.a(s_91), .O(gate192inter4));
  nand2 gate1019(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1020(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1021(.a(N537), .O(gate192inter7));
  inv1  gate1022(.a(N505), .O(gate192inter8));
  nand2 gate1023(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1024(.a(s_91), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1025(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1026(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1027(.a(gate192inter12), .b(gate192inter1), .O(N557));
nand2 gate193( .a(N538), .b(N507), .O(N561) );

  xor2  gate1028(.a(N509), .b(N539), .O(gate194inter0));
  nand2 gate1029(.a(gate194inter0), .b(s_92), .O(gate194inter1));
  and2  gate1030(.a(N509), .b(N539), .O(gate194inter2));
  inv1  gate1031(.a(s_92), .O(gate194inter3));
  inv1  gate1032(.a(s_93), .O(gate194inter4));
  nand2 gate1033(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1034(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1035(.a(N539), .O(gate194inter7));
  inv1  gate1036(.a(N509), .O(gate194inter8));
  nand2 gate1037(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1038(.a(s_93), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1039(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1040(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1041(.a(gate194inter12), .b(gate194inter1), .O(N565));

  xor2  gate524(.a(N540), .b(N488), .O(gate195inter0));
  nand2 gate525(.a(gate195inter0), .b(s_20), .O(gate195inter1));
  and2  gate526(.a(N540), .b(N488), .O(gate195inter2));
  inv1  gate527(.a(s_20), .O(gate195inter3));
  inv1  gate528(.a(s_21), .O(gate195inter4));
  nand2 gate529(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate530(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate531(.a(N488), .O(gate195inter7));
  inv1  gate532(.a(N540), .O(gate195inter8));
  nand2 gate533(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate534(.a(s_21), .b(gate195inter3), .O(gate195inter10));
  nor2  gate535(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate536(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate537(.a(gate195inter12), .b(gate195inter1), .O(N569));

  xor2  gate650(.a(N541), .b(N489), .O(gate196inter0));
  nand2 gate651(.a(gate196inter0), .b(s_38), .O(gate196inter1));
  and2  gate652(.a(N541), .b(N489), .O(gate196inter2));
  inv1  gate653(.a(s_38), .O(gate196inter3));
  inv1  gate654(.a(s_39), .O(gate196inter4));
  nand2 gate655(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate656(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate657(.a(N489), .O(gate196inter7));
  inv1  gate658(.a(N541), .O(gate196inter8));
  nand2 gate659(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate660(.a(s_39), .b(gate196inter3), .O(gate196inter10));
  nor2  gate661(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate662(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate663(.a(gate196inter12), .b(gate196inter1), .O(N573));

  xor2  gate1084(.a(N542), .b(N490), .O(gate197inter0));
  nand2 gate1085(.a(gate197inter0), .b(s_100), .O(gate197inter1));
  and2  gate1086(.a(N542), .b(N490), .O(gate197inter2));
  inv1  gate1087(.a(s_100), .O(gate197inter3));
  inv1  gate1088(.a(s_101), .O(gate197inter4));
  nand2 gate1089(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1090(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1091(.a(N490), .O(gate197inter7));
  inv1  gate1092(.a(N542), .O(gate197inter8));
  nand2 gate1093(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1094(.a(s_101), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1095(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1096(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1097(.a(gate197inter12), .b(gate197inter1), .O(N577));

  xor2  gate1350(.a(N543), .b(N491), .O(gate198inter0));
  nand2 gate1351(.a(gate198inter0), .b(s_138), .O(gate198inter1));
  and2  gate1352(.a(N543), .b(N491), .O(gate198inter2));
  inv1  gate1353(.a(s_138), .O(gate198inter3));
  inv1  gate1354(.a(s_139), .O(gate198inter4));
  nand2 gate1355(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1356(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1357(.a(N491), .O(gate198inter7));
  inv1  gate1358(.a(N543), .O(gate198inter8));
  nand2 gate1359(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1360(.a(s_139), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1361(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1362(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1363(.a(gate198inter12), .b(gate198inter1), .O(N581));
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );

  xor2  gate860(.a(N159), .b(N553), .O(gate204inter0));
  nand2 gate861(.a(gate204inter0), .b(s_68), .O(gate204inter1));
  and2  gate862(.a(N159), .b(N553), .O(gate204inter2));
  inv1  gate863(.a(s_68), .O(gate204inter3));
  inv1  gate864(.a(s_69), .O(gate204inter4));
  nand2 gate865(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate866(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate867(.a(N553), .O(gate204inter7));
  inv1  gate868(.a(N159), .O(gate204inter8));
  nand2 gate869(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate870(.a(s_69), .b(gate204inter3), .O(gate204inter10));
  nor2  gate871(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate872(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate873(.a(gate204inter12), .b(gate204inter1), .O(N590));
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );
nand2 gate207( .a(N557), .b(N165), .O(N597) );
or2 gate208( .a(N557), .b(N165), .O(N600) );
and2 gate209( .a(N246), .b(N557), .O(N605) );

  xor2  gate412(.a(N171), .b(N561), .O(gate210inter0));
  nand2 gate413(.a(gate210inter0), .b(s_4), .O(gate210inter1));
  and2  gate414(.a(N171), .b(N561), .O(gate210inter2));
  inv1  gate415(.a(s_4), .O(gate210inter3));
  inv1  gate416(.a(s_5), .O(gate210inter4));
  nand2 gate417(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate418(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate419(.a(N561), .O(gate210inter7));
  inv1  gate420(.a(N171), .O(gate210inter8));
  nand2 gate421(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate422(.a(s_5), .b(gate210inter3), .O(gate210inter10));
  nor2  gate423(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate424(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate425(.a(gate210inter12), .b(gate210inter1), .O(N606));
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );

  xor2  gate1322(.a(N177), .b(N565), .O(gate213inter0));
  nand2 gate1323(.a(gate213inter0), .b(s_134), .O(gate213inter1));
  and2  gate1324(.a(N177), .b(N565), .O(gate213inter2));
  inv1  gate1325(.a(s_134), .O(gate213inter3));
  inv1  gate1326(.a(s_135), .O(gate213inter4));
  nand2 gate1327(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1328(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1329(.a(N565), .O(gate213inter7));
  inv1  gate1330(.a(N177), .O(gate213inter8));
  nand2 gate1331(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1332(.a(s_135), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1333(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1334(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1335(.a(gate213inter12), .b(gate213inter1), .O(N616));
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );
nand2 gate216( .a(N569), .b(N183), .O(N625) );
or2 gate217( .a(N569), .b(N183), .O(N628) );
and2 gate218( .a(N246), .b(N569), .O(N631) );

  xor2  gate482(.a(N189), .b(N573), .O(gate219inter0));
  nand2 gate483(.a(gate219inter0), .b(s_14), .O(gate219inter1));
  and2  gate484(.a(N189), .b(N573), .O(gate219inter2));
  inv1  gate485(.a(s_14), .O(gate219inter3));
  inv1  gate486(.a(s_15), .O(gate219inter4));
  nand2 gate487(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate488(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate489(.a(N573), .O(gate219inter7));
  inv1  gate490(.a(N189), .O(gate219inter8));
  nand2 gate491(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate492(.a(s_15), .b(gate219inter3), .O(gate219inter10));
  nor2  gate493(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate494(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate495(.a(gate219inter12), .b(gate219inter1), .O(N632));
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );

  xor2  gate608(.a(N195), .b(N577), .O(gate222inter0));
  nand2 gate609(.a(gate222inter0), .b(s_32), .O(gate222inter1));
  and2  gate610(.a(N195), .b(N577), .O(gate222inter2));
  inv1  gate611(.a(s_32), .O(gate222inter3));
  inv1  gate612(.a(s_33), .O(gate222inter4));
  nand2 gate613(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate614(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate615(.a(N577), .O(gate222inter7));
  inv1  gate616(.a(N195), .O(gate222inter8));
  nand2 gate617(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate618(.a(s_33), .b(gate222inter3), .O(gate222inter10));
  nor2  gate619(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate620(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate621(.a(gate222inter12), .b(gate222inter1), .O(N641));
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );

  xor2  gate1392(.a(N201), .b(N581), .O(gate225inter0));
  nand2 gate1393(.a(gate225inter0), .b(s_144), .O(gate225inter1));
  and2  gate1394(.a(N201), .b(N581), .O(gate225inter2));
  inv1  gate1395(.a(s_144), .O(gate225inter3));
  inv1  gate1396(.a(s_145), .O(gate225inter4));
  nand2 gate1397(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1398(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1399(.a(N581), .O(gate225inter7));
  inv1  gate1400(.a(N201), .O(gate225inter8));
  nand2 gate1401(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1402(.a(s_145), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1403(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1404(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1405(.a(gate225inter12), .b(gate225inter1), .O(N651));
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );

  xor2  gate874(.a(N588), .b(N552), .O(gate228inter0));
  nand2 gate875(.a(gate228inter0), .b(s_70), .O(gate228inter1));
  and2  gate876(.a(N588), .b(N552), .O(gate228inter2));
  inv1  gate877(.a(s_70), .O(gate228inter3));
  inv1  gate878(.a(s_71), .O(gate228inter4));
  nand2 gate879(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate880(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate881(.a(N552), .O(gate228inter7));
  inv1  gate882(.a(N588), .O(gate228inter8));
  nand2 gate883(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate884(.a(s_71), .b(gate228inter3), .O(gate228inter10));
  nor2  gate885(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate886(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate887(.a(gate228inter12), .b(gate228inter1), .O(N660));
nor2 gate229( .a(N587), .b(N589), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
and2 gate231( .a(N593), .b(N590), .O(N665) );

  xor2  gate1112(.a(N522), .b(N596), .O(gate232inter0));
  nand2 gate1113(.a(gate232inter0), .b(s_104), .O(gate232inter1));
  and2  gate1114(.a(N522), .b(N596), .O(gate232inter2));
  inv1  gate1115(.a(s_104), .O(gate232inter3));
  inv1  gate1116(.a(s_105), .O(gate232inter4));
  nand2 gate1117(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1118(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1119(.a(N596), .O(gate232inter7));
  inv1  gate1120(.a(N522), .O(gate232inter8));
  nand2 gate1121(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1122(.a(s_105), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1123(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1124(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1125(.a(gate232inter12), .b(gate232inter1), .O(N669));
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );
nor2 gate235( .a(N605), .b(N523), .O(N677) );
inv1 gate236( .a(N606), .O(N678) );
and2 gate237( .a(N609), .b(N606), .O(N682) );

  xor2  gate720(.a(N524), .b(N615), .O(gate238inter0));
  nand2 gate721(.a(gate238inter0), .b(s_48), .O(gate238inter1));
  and2  gate722(.a(N524), .b(N615), .O(gate238inter2));
  inv1  gate723(.a(s_48), .O(gate238inter3));
  inv1  gate724(.a(s_49), .O(gate238inter4));
  nand2 gate725(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate726(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate727(.a(N615), .O(gate238inter7));
  inv1  gate728(.a(N524), .O(gate238inter8));
  nand2 gate729(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate730(.a(s_49), .b(gate238inter3), .O(gate238inter10));
  nor2  gate731(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate732(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate733(.a(gate238inter12), .b(gate238inter1), .O(N686));
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );
nor2 gate241( .a(N624), .b(N525), .O(N696) );
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );

  xor2  gate902(.a(N526), .b(N631), .O(gate244inter0));
  nand2 gate903(.a(gate244inter0), .b(s_74), .O(gate244inter1));
  and2  gate904(.a(N526), .b(N631), .O(gate244inter2));
  inv1  gate905(.a(s_74), .O(gate244inter3));
  inv1  gate906(.a(s_75), .O(gate244inter4));
  nand2 gate907(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate908(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate909(.a(N631), .O(gate244inter7));
  inv1  gate910(.a(N526), .O(gate244inter8));
  nand2 gate911(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate912(.a(s_75), .b(gate244inter3), .O(gate244inter10));
  nor2  gate913(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate914(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate915(.a(gate244inter12), .b(gate244inter1), .O(N704));
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );

  xor2  gate1196(.a(N640), .b(N337), .O(gate247inter0));
  nand2 gate1197(.a(gate247inter0), .b(s_116), .O(gate247inter1));
  and2  gate1198(.a(N640), .b(N337), .O(gate247inter2));
  inv1  gate1199(.a(s_116), .O(gate247inter3));
  inv1  gate1200(.a(s_117), .O(gate247inter4));
  nand2 gate1201(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1202(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1203(.a(N337), .O(gate247inter7));
  inv1  gate1204(.a(N640), .O(gate247inter8));
  nand2 gate1205(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1206(.a(s_117), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1207(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1208(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1209(.a(gate247inter12), .b(gate247inter1), .O(N712));
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );

  xor2  gate1042(.a(N650), .b(N339), .O(gate250inter0));
  nand2 gate1043(.a(gate250inter0), .b(s_94), .O(gate250inter1));
  and2  gate1044(.a(N650), .b(N339), .O(gate250inter2));
  inv1  gate1045(.a(s_94), .O(gate250inter3));
  inv1  gate1046(.a(s_95), .O(gate250inter4));
  nand2 gate1047(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1048(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1049(.a(N339), .O(gate250inter7));
  inv1  gate1050(.a(N650), .O(gate250inter8));
  nand2 gate1051(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1052(.a(s_95), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1053(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1054(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1055(.a(gate250inter12), .b(gate250inter1), .O(N721));
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );
nor2 gate253( .a(N341), .b(N659), .O(N731) );

  xor2  gate496(.a(N261), .b(N654), .O(gate254inter0));
  nand2 gate497(.a(gate254inter0), .b(s_16), .O(gate254inter1));
  and2  gate498(.a(N261), .b(N654), .O(gate254inter2));
  inv1  gate499(.a(s_16), .O(gate254inter3));
  inv1  gate500(.a(s_17), .O(gate254inter4));
  nand2 gate501(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate502(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate503(.a(N654), .O(gate254inter7));
  inv1  gate504(.a(N261), .O(gate254inter8));
  nand2 gate505(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate506(.a(s_17), .b(gate254inter3), .O(gate254inter10));
  nor2  gate507(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate508(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate509(.a(gate254inter12), .b(gate254inter1), .O(N732));
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
and2 gate273( .a(N228), .b(N708), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );
nor2 gate279( .a(N727), .b(N261), .O(N757) );
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );

  xor2  gate706(.a(N722), .b(N644), .O(gate283inter0));
  nand2 gate707(.a(gate283inter0), .b(s_46), .O(gate283inter1));
  and2  gate708(.a(N722), .b(N644), .O(gate283inter2));
  inv1  gate709(.a(s_46), .O(gate283inter3));
  inv1  gate710(.a(s_47), .O(gate283inter4));
  nand2 gate711(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate712(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate713(.a(N644), .O(gate283inter7));
  inv1  gate714(.a(N722), .O(gate283inter8));
  nand2 gate715(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate716(.a(s_47), .b(gate283inter3), .O(gate283inter10));
  nor2  gate717(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate718(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate719(.a(gate283inter12), .b(gate283inter1), .O(N761));

  xor2  gate1000(.a(N713), .b(N635), .O(gate284inter0));
  nand2 gate1001(.a(gate284inter0), .b(s_88), .O(gate284inter1));
  and2  gate1002(.a(N713), .b(N635), .O(gate284inter2));
  inv1  gate1003(.a(s_88), .O(gate284inter3));
  inv1  gate1004(.a(s_89), .O(gate284inter4));
  nand2 gate1005(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1006(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1007(.a(N635), .O(gate284inter7));
  inv1  gate1008(.a(N713), .O(gate284inter8));
  nand2 gate1009(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1010(.a(s_89), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1011(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1012(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1013(.a(gate284inter12), .b(gate284inter1), .O(N762));
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );

  xor2  gate692(.a(N687), .b(N609), .O(gate286inter0));
  nand2 gate693(.a(gate286inter0), .b(s_44), .O(gate286inter1));
  and2  gate694(.a(N687), .b(N609), .O(gate286inter2));
  inv1  gate695(.a(s_44), .O(gate286inter3));
  inv1  gate696(.a(s_45), .O(gate286inter4));
  nand2 gate697(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate698(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate699(.a(N609), .O(gate286inter7));
  inv1  gate700(.a(N687), .O(gate286inter8));
  nand2 gate701(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate702(.a(s_45), .b(gate286inter3), .O(gate286inter10));
  nor2  gate703(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate704(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate705(.a(gate286inter12), .b(gate286inter1), .O(N764));
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );

  xor2  gate1126(.a(N737), .b(N736), .O(gate291inter0));
  nand2 gate1127(.a(gate291inter0), .b(s_106), .O(gate291inter1));
  and2  gate1128(.a(N737), .b(N736), .O(gate291inter2));
  inv1  gate1129(.a(s_106), .O(gate291inter3));
  inv1  gate1130(.a(s_107), .O(gate291inter4));
  nand2 gate1131(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1132(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1133(.a(N736), .O(gate291inter7));
  inv1  gate1134(.a(N737), .O(gate291inter8));
  nand2 gate1135(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1136(.a(s_107), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1137(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1138(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1139(.a(gate291inter12), .b(gate291inter1), .O(N769));
nor2 gate292( .a(N739), .b(N740), .O(N770) );

  xor2  gate594(.a(N743), .b(N742), .O(gate293inter0));
  nand2 gate595(.a(gate293inter0), .b(s_30), .O(gate293inter1));
  and2  gate596(.a(N743), .b(N742), .O(gate293inter2));
  inv1  gate597(.a(s_30), .O(gate293inter3));
  inv1  gate598(.a(s_31), .O(gate293inter4));
  nand2 gate599(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate600(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate601(.a(N742), .O(gate293inter7));
  inv1  gate602(.a(N743), .O(gate293inter8));
  nand2 gate603(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate604(.a(s_31), .b(gate293inter3), .O(gate293inter10));
  nor2  gate605(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate606(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate607(.a(gate293inter12), .b(gate293inter1), .O(N771));

  xor2  gate1098(.a(N746), .b(N745), .O(gate294inter0));
  nand2 gate1099(.a(gate294inter0), .b(s_102), .O(gate294inter1));
  and2  gate1100(.a(N746), .b(N745), .O(gate294inter2));
  inv1  gate1101(.a(s_102), .O(gate294inter3));
  inv1  gate1102(.a(s_103), .O(gate294inter4));
  nand2 gate1103(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1104(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1105(.a(N745), .O(gate294inter7));
  inv1  gate1106(.a(N746), .O(gate294inter8));
  nand2 gate1107(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1108(.a(s_103), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1109(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1110(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1111(.a(gate294inter12), .b(gate294inter1), .O(N772));
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );

  xor2  gate1252(.a(N749), .b(N748), .O(gate296inter0));
  nand2 gate1253(.a(gate296inter0), .b(s_124), .O(gate296inter1));
  and2  gate1254(.a(N749), .b(N748), .O(gate296inter2));
  inv1  gate1255(.a(s_124), .O(gate296inter3));
  inv1  gate1256(.a(s_125), .O(gate296inter4));
  nand2 gate1257(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1258(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1259(.a(N748), .O(gate296inter7));
  inv1  gate1260(.a(N749), .O(gate296inter8));
  nand2 gate1261(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1262(.a(s_125), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1263(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1264(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1265(.a(gate296inter12), .b(gate296inter1), .O(N777));
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );

  xor2  gate580(.a(N752), .b(N751), .O(gate298inter0));
  nand2 gate581(.a(gate298inter0), .b(s_28), .O(gate298inter1));
  and2  gate582(.a(N752), .b(N751), .O(gate298inter2));
  inv1  gate583(.a(s_28), .O(gate298inter3));
  inv1  gate584(.a(s_29), .O(gate298inter4));
  nand2 gate585(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate586(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate587(.a(N751), .O(gate298inter7));
  inv1  gate588(.a(N752), .O(gate298inter8));
  nand2 gate589(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate590(.a(s_29), .b(gate298inter3), .O(gate298inter10));
  nor2  gate591(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate592(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate593(.a(gate298inter12), .b(gate298inter1), .O(N781));
nand2 gate299( .a(N756), .b(N732), .O(N782) );

  xor2  gate1364(.a(N755), .b(N754), .O(gate300inter0));
  nand2 gate1365(.a(gate300inter0), .b(s_140), .O(gate300inter1));
  and2  gate1366(.a(N755), .b(N754), .O(gate300inter2));
  inv1  gate1367(.a(s_140), .O(gate300inter3));
  inv1  gate1368(.a(s_141), .O(gate300inter4));
  nand2 gate1369(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate1370(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate1371(.a(N754), .O(gate300inter7));
  inv1  gate1372(.a(N755), .O(gate300inter8));
  nand2 gate1373(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate1374(.a(s_141), .b(gate300inter3), .O(gate300inter10));
  nor2  gate1375(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate1376(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate1377(.a(gate300inter12), .b(gate300inter1), .O(N785));
nor2 gate301( .a(N757), .b(N758), .O(N786) );
nor2 gate302( .a(N759), .b(N760), .O(N787) );

  xor2  gate440(.a(N773), .b(N700), .O(gate303inter0));
  nand2 gate441(.a(gate303inter0), .b(s_8), .O(gate303inter1));
  and2  gate442(.a(N773), .b(N700), .O(gate303inter2));
  inv1  gate443(.a(s_8), .O(gate303inter3));
  inv1  gate444(.a(s_9), .O(gate303inter4));
  nand2 gate445(.a(gate303inter4), .b(gate303inter3), .O(gate303inter5));
  nor2  gate446(.a(gate303inter5), .b(gate303inter2), .O(gate303inter6));
  inv1  gate447(.a(N700), .O(gate303inter7));
  inv1  gate448(.a(N773), .O(gate303inter8));
  nand2 gate449(.a(gate303inter8), .b(gate303inter7), .O(gate303inter9));
  nand2 gate450(.a(s_9), .b(gate303inter3), .O(gate303inter10));
  nor2  gate451(.a(gate303inter10), .b(gate303inter9), .O(gate303inter11));
  nor2  gate452(.a(gate303inter11), .b(gate303inter6), .O(gate303inter12));
  nand2 gate453(.a(gate303inter12), .b(gate303inter1), .O(N788));
and2 gate304( .a(N700), .b(N773), .O(N789) );
nor2 gate305( .a(N708), .b(N778), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );

  xor2  gate888(.a(N782), .b(N717), .O(gate307inter0));
  nand2 gate889(.a(gate307inter0), .b(s_72), .O(gate307inter1));
  and2  gate890(.a(N782), .b(N717), .O(gate307inter2));
  inv1  gate891(.a(s_72), .O(gate307inter3));
  inv1  gate892(.a(s_73), .O(gate307inter4));
  nand2 gate893(.a(gate307inter4), .b(gate307inter3), .O(gate307inter5));
  nor2  gate894(.a(gate307inter5), .b(gate307inter2), .O(gate307inter6));
  inv1  gate895(.a(N717), .O(gate307inter7));
  inv1  gate896(.a(N782), .O(gate307inter8));
  nand2 gate897(.a(gate307inter8), .b(gate307inter7), .O(gate307inter9));
  nand2 gate898(.a(s_73), .b(gate307inter3), .O(gate307inter10));
  nor2  gate899(.a(gate307inter10), .b(gate307inter9), .O(gate307inter11));
  nor2  gate900(.a(gate307inter11), .b(gate307inter6), .O(gate307inter12));
  nand2 gate901(.a(gate307inter12), .b(gate307inter1), .O(N792));
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );

  xor2  gate1168(.a(N773), .b(N628), .O(gate310inter0));
  nand2 gate1169(.a(gate310inter0), .b(s_112), .O(gate310inter1));
  and2  gate1170(.a(N773), .b(N628), .O(gate310inter2));
  inv1  gate1171(.a(s_112), .O(gate310inter3));
  inv1  gate1172(.a(s_113), .O(gate310inter4));
  nand2 gate1173(.a(gate310inter4), .b(gate310inter3), .O(gate310inter5));
  nor2  gate1174(.a(gate310inter5), .b(gate310inter2), .O(gate310inter6));
  inv1  gate1175(.a(N628), .O(gate310inter7));
  inv1  gate1176(.a(N773), .O(gate310inter8));
  nand2 gate1177(.a(gate310inter8), .b(gate310inter7), .O(gate310inter9));
  nand2 gate1178(.a(s_113), .b(gate310inter3), .O(gate310inter10));
  nor2  gate1179(.a(gate310inter10), .b(gate310inter9), .O(gate310inter11));
  nor2  gate1180(.a(gate310inter11), .b(gate310inter6), .O(gate310inter12));
  nand2 gate1181(.a(gate310inter12), .b(gate310inter1), .O(N795));

  xor2  gate986(.a(N747), .b(N795), .O(gate311inter0));
  nand2 gate987(.a(gate311inter0), .b(s_86), .O(gate311inter1));
  and2  gate988(.a(N747), .b(N795), .O(gate311inter2));
  inv1  gate989(.a(s_86), .O(gate311inter3));
  inv1  gate990(.a(s_87), .O(gate311inter4));
  nand2 gate991(.a(gate311inter4), .b(gate311inter3), .O(gate311inter5));
  nor2  gate992(.a(gate311inter5), .b(gate311inter2), .O(gate311inter6));
  inv1  gate993(.a(N795), .O(gate311inter7));
  inv1  gate994(.a(N747), .O(gate311inter8));
  nand2 gate995(.a(gate311inter8), .b(gate311inter7), .O(gate311inter9));
  nand2 gate996(.a(s_87), .b(gate311inter3), .O(gate311inter10));
  nor2  gate997(.a(gate311inter10), .b(gate311inter9), .O(gate311inter11));
  nor2  gate998(.a(gate311inter11), .b(gate311inter6), .O(gate311inter12));
  nand2 gate999(.a(gate311inter12), .b(gate311inter1), .O(N796));

  xor2  gate426(.a(N789), .b(N788), .O(gate312inter0));
  nand2 gate427(.a(gate312inter0), .b(s_6), .O(gate312inter1));
  and2  gate428(.a(N789), .b(N788), .O(gate312inter2));
  inv1  gate429(.a(s_6), .O(gate312inter3));
  inv1  gate430(.a(s_7), .O(gate312inter4));
  nand2 gate431(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate432(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate433(.a(N788), .O(gate312inter7));
  inv1  gate434(.a(N789), .O(gate312inter8));
  nand2 gate435(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate436(.a(s_7), .b(gate312inter3), .O(gate312inter10));
  nor2  gate437(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate438(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate439(.a(gate312inter12), .b(gate312inter1), .O(N802));
nor2 gate313( .a(N790), .b(N791), .O(N803) );
nor2 gate314( .a(N792), .b(N793), .O(N804) );
nor2 gate315( .a(N340), .b(N794), .O(N805) );
nor2 gate316( .a(N692), .b(N796), .O(N806) );
and2 gate317( .a(N692), .b(N796), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );

  xor2  gate832(.a(N796), .b(N619), .O(gate322inter0));
  nand2 gate833(.a(gate322inter0), .b(s_64), .O(gate322inter1));
  and2  gate834(.a(N796), .b(N619), .O(gate322inter2));
  inv1  gate835(.a(s_64), .O(gate322inter3));
  inv1  gate836(.a(s_65), .O(gate322inter4));
  nand2 gate837(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate838(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate839(.a(N619), .O(gate322inter7));
  inv1  gate840(.a(N796), .O(gate322inter8));
  nand2 gate841(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate842(.a(s_65), .b(gate322inter3), .O(gate322inter10));
  nor2  gate843(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate844(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate845(.a(gate322inter12), .b(gate322inter1), .O(N812));
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );

  xor2  gate846(.a(N812), .b(N744), .O(gate327inter0));
  nand2 gate847(.a(gate327inter0), .b(s_66), .O(gate327inter1));
  and2  gate848(.a(N812), .b(N744), .O(gate327inter2));
  inv1  gate849(.a(s_66), .O(gate327inter3));
  inv1  gate850(.a(s_67), .O(gate327inter4));
  nand2 gate851(.a(gate327inter4), .b(gate327inter3), .O(gate327inter5));
  nor2  gate852(.a(gate327inter5), .b(gate327inter2), .O(gate327inter6));
  inv1  gate853(.a(N744), .O(gate327inter7));
  inv1  gate854(.a(N812), .O(gate327inter8));
  nand2 gate855(.a(gate327inter8), .b(gate327inter7), .O(gate327inter9));
  nand2 gate856(.a(s_67), .b(gate327inter3), .O(gate327inter10));
  nor2  gate857(.a(gate327inter10), .b(gate327inter9), .O(gate327inter11));
  nor2  gate858(.a(gate327inter11), .b(gate327inter6), .O(gate327inter12));
  nand2 gate859(.a(gate327inter12), .b(gate327inter1), .O(N822));
nor2 gate328( .a(N806), .b(N807), .O(N825) );
nor2 gate329( .a(N335), .b(N808), .O(N826) );

  xor2  gate1336(.a(N809), .b(N336), .O(gate330inter0));
  nand2 gate1337(.a(gate330inter0), .b(s_136), .O(gate330inter1));
  and2  gate1338(.a(N809), .b(N336), .O(gate330inter2));
  inv1  gate1339(.a(s_136), .O(gate330inter3));
  inv1  gate1340(.a(s_137), .O(gate330inter4));
  nand2 gate1341(.a(gate330inter4), .b(gate330inter3), .O(gate330inter5));
  nor2  gate1342(.a(gate330inter5), .b(gate330inter2), .O(gate330inter6));
  inv1  gate1343(.a(N336), .O(gate330inter7));
  inv1  gate1344(.a(N809), .O(gate330inter8));
  nand2 gate1345(.a(gate330inter8), .b(gate330inter7), .O(gate330inter9));
  nand2 gate1346(.a(s_137), .b(gate330inter3), .O(gate330inter10));
  nor2  gate1347(.a(gate330inter10), .b(gate330inter9), .O(gate330inter11));
  nor2  gate1348(.a(gate330inter11), .b(gate330inter6), .O(gate330inter12));
  nand2 gate1349(.a(gate330inter12), .b(gate330inter1), .O(N827));

  xor2  gate1434(.a(N810), .b(N338), .O(gate331inter0));
  nand2 gate1435(.a(gate331inter0), .b(s_150), .O(gate331inter1));
  and2  gate1436(.a(N810), .b(N338), .O(gate331inter2));
  inv1  gate1437(.a(s_150), .O(gate331inter3));
  inv1  gate1438(.a(s_151), .O(gate331inter4));
  nand2 gate1439(.a(gate331inter4), .b(gate331inter3), .O(gate331inter5));
  nor2  gate1440(.a(gate331inter5), .b(gate331inter2), .O(gate331inter6));
  inv1  gate1441(.a(N338), .O(gate331inter7));
  inv1  gate1442(.a(N810), .O(gate331inter8));
  nand2 gate1443(.a(gate331inter8), .b(gate331inter7), .O(gate331inter9));
  nand2 gate1444(.a(s_151), .b(gate331inter3), .O(gate331inter10));
  nor2  gate1445(.a(gate331inter10), .b(gate331inter9), .O(gate331inter11));
  nor2  gate1446(.a(gate331inter11), .b(gate331inter6), .O(gate331inter12));
  nand2 gate1447(.a(gate331inter12), .b(gate331inter1), .O(N828));
inv1 gate332( .a(N811), .O(N829) );
nor2 gate333( .a(N665), .b(N815), .O(N830) );
and2 gate334( .a(N665), .b(N815), .O(N831) );

  xor2  gate1056(.a(N819), .b(N673), .O(gate335inter0));
  nand2 gate1057(.a(gate335inter0), .b(s_96), .O(gate335inter1));
  and2  gate1058(.a(N819), .b(N673), .O(gate335inter2));
  inv1  gate1059(.a(s_96), .O(gate335inter3));
  inv1  gate1060(.a(s_97), .O(gate335inter4));
  nand2 gate1061(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate1062(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate1063(.a(N673), .O(gate335inter7));
  inv1  gate1064(.a(N819), .O(gate335inter8));
  nand2 gate1065(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate1066(.a(s_97), .b(gate335inter3), .O(gate335inter10));
  nor2  gate1067(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate1068(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate1069(.a(gate335inter12), .b(gate335inter1), .O(N832));
and2 gate336( .a(N673), .b(N819), .O(N833) );

  xor2  gate510(.a(N822), .b(N682), .O(gate337inter0));
  nand2 gate511(.a(gate337inter0), .b(s_18), .O(gate337inter1));
  and2  gate512(.a(N822), .b(N682), .O(gate337inter2));
  inv1  gate513(.a(s_18), .O(gate337inter3));
  inv1  gate514(.a(s_19), .O(gate337inter4));
  nand2 gate515(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate516(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate517(.a(N682), .O(gate337inter7));
  inv1  gate518(.a(N822), .O(gate337inter8));
  nand2 gate519(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate520(.a(s_19), .b(gate337inter3), .O(gate337inter10));
  nor2  gate521(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate522(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate523(.a(gate337inter12), .b(gate337inter1), .O(N834));
and2 gate338( .a(N682), .b(N822), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
nand2 gate344( .a(N815), .b(N593), .O(N841) );
nor2 gate345( .a(N830), .b(N831), .O(N842) );

  xor2  gate566(.a(N833), .b(N832), .O(gate346inter0));
  nand2 gate567(.a(gate346inter0), .b(s_26), .O(gate346inter1));
  and2  gate568(.a(N833), .b(N832), .O(gate346inter2));
  inv1  gate569(.a(s_26), .O(gate346inter3));
  inv1  gate570(.a(s_27), .O(gate346inter4));
  nand2 gate571(.a(gate346inter4), .b(gate346inter3), .O(gate346inter5));
  nor2  gate572(.a(gate346inter5), .b(gate346inter2), .O(gate346inter6));
  inv1  gate573(.a(N832), .O(gate346inter7));
  inv1  gate574(.a(N833), .O(gate346inter8));
  nand2 gate575(.a(gate346inter8), .b(gate346inter7), .O(gate346inter9));
  nand2 gate576(.a(s_27), .b(gate346inter3), .O(gate346inter10));
  nor2  gate577(.a(gate346inter10), .b(gate346inter9), .O(gate346inter11));
  nor2  gate578(.a(gate346inter11), .b(gate346inter6), .O(gate346inter12));
  nand2 gate579(.a(gate346inter12), .b(gate346inter1), .O(N843));

  xor2  gate1070(.a(N835), .b(N834), .O(gate347inter0));
  nand2 gate1071(.a(gate347inter0), .b(s_98), .O(gate347inter1));
  and2  gate1072(.a(N835), .b(N834), .O(gate347inter2));
  inv1  gate1073(.a(s_98), .O(gate347inter3));
  inv1  gate1074(.a(s_99), .O(gate347inter4));
  nand2 gate1075(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate1076(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate1077(.a(N834), .O(gate347inter7));
  inv1  gate1078(.a(N835), .O(gate347inter8));
  nand2 gate1079(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate1080(.a(s_99), .b(gate347inter3), .O(gate347inter10));
  nor2  gate1081(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate1082(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate1083(.a(gate347inter12), .b(gate347inter1), .O(N844));

  xor2  gate1140(.a(N836), .b(N334), .O(gate348inter0));
  nand2 gate1141(.a(gate348inter0), .b(s_108), .O(gate348inter1));
  and2  gate1142(.a(N836), .b(N334), .O(gate348inter2));
  inv1  gate1143(.a(s_108), .O(gate348inter3));
  inv1  gate1144(.a(s_109), .O(gate348inter4));
  nand2 gate1145(.a(gate348inter4), .b(gate348inter3), .O(gate348inter5));
  nor2  gate1146(.a(gate348inter5), .b(gate348inter2), .O(gate348inter6));
  inv1  gate1147(.a(N334), .O(gate348inter7));
  inv1  gate1148(.a(N836), .O(gate348inter8));
  nand2 gate1149(.a(gate348inter8), .b(gate348inter7), .O(gate348inter9));
  nand2 gate1150(.a(s_109), .b(gate348inter3), .O(gate348inter10));
  nor2  gate1151(.a(gate348inter10), .b(gate348inter9), .O(gate348inter11));
  nor2  gate1152(.a(gate348inter11), .b(gate348inter6), .O(gate348inter12));
  nand2 gate1153(.a(gate348inter12), .b(gate348inter1), .O(N845));
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
and2 gate354( .a(N219), .b(N842), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );

  xor2  gate1182(.a(N851), .b(N417), .O(gate362inter0));
  nand2 gate1183(.a(gate362inter0), .b(s_114), .O(gate362inter1));
  and2  gate1184(.a(N851), .b(N417), .O(gate362inter2));
  inv1  gate1185(.a(s_114), .O(gate362inter3));
  inv1  gate1186(.a(s_115), .O(gate362inter4));
  nand2 gate1187(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate1188(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate1189(.a(N417), .O(gate362inter7));
  inv1  gate1190(.a(N851), .O(gate362inter8));
  nand2 gate1191(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate1192(.a(s_115), .b(gate362inter3), .O(gate362inter10));
  nor2  gate1193(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate1194(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate1195(.a(gate362inter12), .b(gate362inter1), .O(N859));
nor2 gate363( .a(N332), .b(N852), .O(N860) );
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

endmodule