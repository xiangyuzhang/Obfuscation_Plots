module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2647(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2648(.a(gate10inter0), .b(s_300), .O(gate10inter1));
  and2  gate2649(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2650(.a(s_300), .O(gate10inter3));
  inv1  gate2651(.a(s_301), .O(gate10inter4));
  nand2 gate2652(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2653(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2654(.a(G3), .O(gate10inter7));
  inv1  gate2655(.a(G4), .O(gate10inter8));
  nand2 gate2656(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2657(.a(s_301), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2658(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2659(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2660(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate2325(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2326(.a(gate11inter0), .b(s_254), .O(gate11inter1));
  and2  gate2327(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2328(.a(s_254), .O(gate11inter3));
  inv1  gate2329(.a(s_255), .O(gate11inter4));
  nand2 gate2330(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2331(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2332(.a(G5), .O(gate11inter7));
  inv1  gate2333(.a(G6), .O(gate11inter8));
  nand2 gate2334(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2335(.a(s_255), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2336(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2337(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2338(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1863(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1864(.a(gate12inter0), .b(s_188), .O(gate12inter1));
  and2  gate1865(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1866(.a(s_188), .O(gate12inter3));
  inv1  gate1867(.a(s_189), .O(gate12inter4));
  nand2 gate1868(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1869(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1870(.a(G7), .O(gate12inter7));
  inv1  gate1871(.a(G8), .O(gate12inter8));
  nand2 gate1872(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1873(.a(s_189), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1874(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1875(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1876(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2801(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2802(.a(gate13inter0), .b(s_322), .O(gate13inter1));
  and2  gate2803(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2804(.a(s_322), .O(gate13inter3));
  inv1  gate2805(.a(s_323), .O(gate13inter4));
  nand2 gate2806(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2807(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2808(.a(G9), .O(gate13inter7));
  inv1  gate2809(.a(G10), .O(gate13inter8));
  nand2 gate2810(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2811(.a(s_323), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2812(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2813(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2814(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2857(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2858(.a(gate18inter0), .b(s_330), .O(gate18inter1));
  and2  gate2859(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2860(.a(s_330), .O(gate18inter3));
  inv1  gate2861(.a(s_331), .O(gate18inter4));
  nand2 gate2862(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2863(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2864(.a(G19), .O(gate18inter7));
  inv1  gate2865(.a(G20), .O(gate18inter8));
  nand2 gate2866(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2867(.a(s_331), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2868(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2869(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2870(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2507(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2508(.a(gate21inter0), .b(s_280), .O(gate21inter1));
  and2  gate2509(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2510(.a(s_280), .O(gate21inter3));
  inv1  gate2511(.a(s_281), .O(gate21inter4));
  nand2 gate2512(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2513(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2514(.a(G25), .O(gate21inter7));
  inv1  gate2515(.a(G26), .O(gate21inter8));
  nand2 gate2516(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2517(.a(s_281), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2518(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2519(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2520(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2381(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2382(.a(gate25inter0), .b(s_262), .O(gate25inter1));
  and2  gate2383(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2384(.a(s_262), .O(gate25inter3));
  inv1  gate2385(.a(s_263), .O(gate25inter4));
  nand2 gate2386(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2387(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2388(.a(G1), .O(gate25inter7));
  inv1  gate2389(.a(G5), .O(gate25inter8));
  nand2 gate2390(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2391(.a(s_263), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2392(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2393(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2394(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate2297(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2298(.a(gate26inter0), .b(s_250), .O(gate26inter1));
  and2  gate2299(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2300(.a(s_250), .O(gate26inter3));
  inv1  gate2301(.a(s_251), .O(gate26inter4));
  nand2 gate2302(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2303(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2304(.a(G9), .O(gate26inter7));
  inv1  gate2305(.a(G13), .O(gate26inter8));
  nand2 gate2306(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2307(.a(s_251), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2308(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2309(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2310(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1485(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1486(.a(gate29inter0), .b(s_134), .O(gate29inter1));
  and2  gate1487(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1488(.a(s_134), .O(gate29inter3));
  inv1  gate1489(.a(s_135), .O(gate29inter4));
  nand2 gate1490(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1491(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1492(.a(G3), .O(gate29inter7));
  inv1  gate1493(.a(G7), .O(gate29inter8));
  nand2 gate1494(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1495(.a(s_135), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1496(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1497(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1498(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2171(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2172(.a(gate36inter0), .b(s_232), .O(gate36inter1));
  and2  gate2173(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2174(.a(s_232), .O(gate36inter3));
  inv1  gate2175(.a(s_233), .O(gate36inter4));
  nand2 gate2176(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2177(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2178(.a(G26), .O(gate36inter7));
  inv1  gate2179(.a(G30), .O(gate36inter8));
  nand2 gate2180(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2181(.a(s_233), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2182(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2183(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2184(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2227(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2228(.a(gate40inter0), .b(s_240), .O(gate40inter1));
  and2  gate2229(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2230(.a(s_240), .O(gate40inter3));
  inv1  gate2231(.a(s_241), .O(gate40inter4));
  nand2 gate2232(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2233(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2234(.a(G28), .O(gate40inter7));
  inv1  gate2235(.a(G32), .O(gate40inter8));
  nand2 gate2236(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2237(.a(s_241), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2238(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2239(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2240(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2983(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2984(.a(gate41inter0), .b(s_348), .O(gate41inter1));
  and2  gate2985(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2986(.a(s_348), .O(gate41inter3));
  inv1  gate2987(.a(s_349), .O(gate41inter4));
  nand2 gate2988(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2989(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2990(.a(G1), .O(gate41inter7));
  inv1  gate2991(.a(G266), .O(gate41inter8));
  nand2 gate2992(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2993(.a(s_349), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2994(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2995(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2996(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2353(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2354(.a(gate42inter0), .b(s_258), .O(gate42inter1));
  and2  gate2355(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2356(.a(s_258), .O(gate42inter3));
  inv1  gate2357(.a(s_259), .O(gate42inter4));
  nand2 gate2358(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2359(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2360(.a(G2), .O(gate42inter7));
  inv1  gate2361(.a(G266), .O(gate42inter8));
  nand2 gate2362(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2363(.a(s_259), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2364(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2365(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2366(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2577(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2578(.a(gate44inter0), .b(s_290), .O(gate44inter1));
  and2  gate2579(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2580(.a(s_290), .O(gate44inter3));
  inv1  gate2581(.a(s_291), .O(gate44inter4));
  nand2 gate2582(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2583(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2584(.a(G4), .O(gate44inter7));
  inv1  gate2585(.a(G269), .O(gate44inter8));
  nand2 gate2586(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2587(.a(s_291), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2588(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2589(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2590(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1121(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1122(.a(gate47inter0), .b(s_82), .O(gate47inter1));
  and2  gate1123(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1124(.a(s_82), .O(gate47inter3));
  inv1  gate1125(.a(s_83), .O(gate47inter4));
  nand2 gate1126(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1127(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1128(.a(G7), .O(gate47inter7));
  inv1  gate1129(.a(G275), .O(gate47inter8));
  nand2 gate1130(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1131(.a(s_83), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1132(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1133(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1134(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1555(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1556(.a(gate49inter0), .b(s_144), .O(gate49inter1));
  and2  gate1557(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1558(.a(s_144), .O(gate49inter3));
  inv1  gate1559(.a(s_145), .O(gate49inter4));
  nand2 gate1560(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1561(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1562(.a(G9), .O(gate49inter7));
  inv1  gate1563(.a(G278), .O(gate49inter8));
  nand2 gate1564(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1565(.a(s_145), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1566(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1567(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1568(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1751(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1752(.a(gate51inter0), .b(s_172), .O(gate51inter1));
  and2  gate1753(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1754(.a(s_172), .O(gate51inter3));
  inv1  gate1755(.a(s_173), .O(gate51inter4));
  nand2 gate1756(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1757(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1758(.a(G11), .O(gate51inter7));
  inv1  gate1759(.a(G281), .O(gate51inter8));
  nand2 gate1760(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1761(.a(s_173), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1762(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1763(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1764(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2843(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2844(.a(gate53inter0), .b(s_328), .O(gate53inter1));
  and2  gate2845(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2846(.a(s_328), .O(gate53inter3));
  inv1  gate2847(.a(s_329), .O(gate53inter4));
  nand2 gate2848(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2849(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2850(.a(G13), .O(gate53inter7));
  inv1  gate2851(.a(G284), .O(gate53inter8));
  nand2 gate2852(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2853(.a(s_329), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2854(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2855(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2856(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate2409(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2410(.a(gate54inter0), .b(s_266), .O(gate54inter1));
  and2  gate2411(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2412(.a(s_266), .O(gate54inter3));
  inv1  gate2413(.a(s_267), .O(gate54inter4));
  nand2 gate2414(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2415(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2416(.a(G14), .O(gate54inter7));
  inv1  gate2417(.a(G284), .O(gate54inter8));
  nand2 gate2418(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2419(.a(s_267), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2420(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2421(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2422(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1597(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1598(.a(gate55inter0), .b(s_150), .O(gate55inter1));
  and2  gate1599(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1600(.a(s_150), .O(gate55inter3));
  inv1  gate1601(.a(s_151), .O(gate55inter4));
  nand2 gate1602(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1603(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1604(.a(G15), .O(gate55inter7));
  inv1  gate1605(.a(G287), .O(gate55inter8));
  nand2 gate1606(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1607(.a(s_151), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1608(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1609(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1610(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1079(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1080(.a(gate58inter0), .b(s_76), .O(gate58inter1));
  and2  gate1081(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1082(.a(s_76), .O(gate58inter3));
  inv1  gate1083(.a(s_77), .O(gate58inter4));
  nand2 gate1084(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1085(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1086(.a(G18), .O(gate58inter7));
  inv1  gate1087(.a(G290), .O(gate58inter8));
  nand2 gate1088(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1089(.a(s_77), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1090(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1091(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1092(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1681(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1682(.a(gate59inter0), .b(s_162), .O(gate59inter1));
  and2  gate1683(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1684(.a(s_162), .O(gate59inter3));
  inv1  gate1685(.a(s_163), .O(gate59inter4));
  nand2 gate1686(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1687(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1688(.a(G19), .O(gate59inter7));
  inv1  gate1689(.a(G293), .O(gate59inter8));
  nand2 gate1690(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1691(.a(s_163), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1692(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1693(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1694(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate2535(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2536(.a(gate60inter0), .b(s_284), .O(gate60inter1));
  and2  gate2537(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2538(.a(s_284), .O(gate60inter3));
  inv1  gate2539(.a(s_285), .O(gate60inter4));
  nand2 gate2540(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2541(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2542(.a(G20), .O(gate60inter7));
  inv1  gate2543(.a(G293), .O(gate60inter8));
  nand2 gate2544(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2545(.a(s_285), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2546(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2547(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2548(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2941(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2942(.a(gate61inter0), .b(s_342), .O(gate61inter1));
  and2  gate2943(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2944(.a(s_342), .O(gate61inter3));
  inv1  gate2945(.a(s_343), .O(gate61inter4));
  nand2 gate2946(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2947(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2948(.a(G21), .O(gate61inter7));
  inv1  gate2949(.a(G296), .O(gate61inter8));
  nand2 gate2950(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2951(.a(s_343), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2952(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2953(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2954(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2689(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2690(.a(gate62inter0), .b(s_306), .O(gate62inter1));
  and2  gate2691(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2692(.a(s_306), .O(gate62inter3));
  inv1  gate2693(.a(s_307), .O(gate62inter4));
  nand2 gate2694(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2695(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2696(.a(G22), .O(gate62inter7));
  inv1  gate2697(.a(G296), .O(gate62inter8));
  nand2 gate2698(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2699(.a(s_307), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2700(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2701(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2702(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2423(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2424(.a(gate64inter0), .b(s_268), .O(gate64inter1));
  and2  gate2425(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2426(.a(s_268), .O(gate64inter3));
  inv1  gate2427(.a(s_269), .O(gate64inter4));
  nand2 gate2428(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2429(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2430(.a(G24), .O(gate64inter7));
  inv1  gate2431(.a(G299), .O(gate64inter8));
  nand2 gate2432(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2433(.a(s_269), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2434(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2435(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2436(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1443(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1444(.a(gate71inter0), .b(s_128), .O(gate71inter1));
  and2  gate1445(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1446(.a(s_128), .O(gate71inter3));
  inv1  gate1447(.a(s_129), .O(gate71inter4));
  nand2 gate1448(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1449(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1450(.a(G31), .O(gate71inter7));
  inv1  gate1451(.a(G311), .O(gate71inter8));
  nand2 gate1452(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1453(.a(s_129), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1454(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1455(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1456(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate743(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate744(.a(gate72inter0), .b(s_28), .O(gate72inter1));
  and2  gate745(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate746(.a(s_28), .O(gate72inter3));
  inv1  gate747(.a(s_29), .O(gate72inter4));
  nand2 gate748(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate749(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate750(.a(G32), .O(gate72inter7));
  inv1  gate751(.a(G311), .O(gate72inter8));
  nand2 gate752(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate753(.a(s_29), .b(gate72inter3), .O(gate72inter10));
  nor2  gate754(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate755(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate756(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate2549(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2550(.a(gate73inter0), .b(s_286), .O(gate73inter1));
  and2  gate2551(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2552(.a(s_286), .O(gate73inter3));
  inv1  gate2553(.a(s_287), .O(gate73inter4));
  nand2 gate2554(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2555(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2556(.a(G1), .O(gate73inter7));
  inv1  gate2557(.a(G314), .O(gate73inter8));
  nand2 gate2558(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2559(.a(s_287), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2560(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2561(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2562(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1639(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1640(.a(gate79inter0), .b(s_156), .O(gate79inter1));
  and2  gate1641(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1642(.a(s_156), .O(gate79inter3));
  inv1  gate1643(.a(s_157), .O(gate79inter4));
  nand2 gate1644(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1645(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1646(.a(G10), .O(gate79inter7));
  inv1  gate1647(.a(G323), .O(gate79inter8));
  nand2 gate1648(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1649(.a(s_157), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1650(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1651(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1652(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1205(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1206(.a(gate80inter0), .b(s_94), .O(gate80inter1));
  and2  gate1207(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1208(.a(s_94), .O(gate80inter3));
  inv1  gate1209(.a(s_95), .O(gate80inter4));
  nand2 gate1210(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1211(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1212(.a(G14), .O(gate80inter7));
  inv1  gate1213(.a(G323), .O(gate80inter8));
  nand2 gate1214(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1215(.a(s_95), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1216(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1217(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1218(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate953(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate954(.a(gate84inter0), .b(s_58), .O(gate84inter1));
  and2  gate955(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate956(.a(s_58), .O(gate84inter3));
  inv1  gate957(.a(s_59), .O(gate84inter4));
  nand2 gate958(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate959(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate960(.a(G15), .O(gate84inter7));
  inv1  gate961(.a(G329), .O(gate84inter8));
  nand2 gate962(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate963(.a(s_59), .b(gate84inter3), .O(gate84inter10));
  nor2  gate964(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate965(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate966(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2731(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2732(.a(gate90inter0), .b(s_312), .O(gate90inter1));
  and2  gate2733(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2734(.a(s_312), .O(gate90inter3));
  inv1  gate2735(.a(s_313), .O(gate90inter4));
  nand2 gate2736(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2737(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2738(.a(G21), .O(gate90inter7));
  inv1  gate2739(.a(G338), .O(gate90inter8));
  nand2 gate2740(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2741(.a(s_313), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2742(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2743(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2744(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1457(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1458(.a(gate97inter0), .b(s_130), .O(gate97inter1));
  and2  gate1459(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1460(.a(s_130), .O(gate97inter3));
  inv1  gate1461(.a(s_131), .O(gate97inter4));
  nand2 gate1462(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1463(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1464(.a(G19), .O(gate97inter7));
  inv1  gate1465(.a(G350), .O(gate97inter8));
  nand2 gate1466(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1467(.a(s_131), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1468(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1469(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1470(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate3025(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate3026(.a(gate99inter0), .b(s_354), .O(gate99inter1));
  and2  gate3027(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate3028(.a(s_354), .O(gate99inter3));
  inv1  gate3029(.a(s_355), .O(gate99inter4));
  nand2 gate3030(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate3031(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate3032(.a(G27), .O(gate99inter7));
  inv1  gate3033(.a(G353), .O(gate99inter8));
  nand2 gate3034(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate3035(.a(s_355), .b(gate99inter3), .O(gate99inter10));
  nor2  gate3036(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate3037(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate3038(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1947(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1948(.a(gate100inter0), .b(s_200), .O(gate100inter1));
  and2  gate1949(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1950(.a(s_200), .O(gate100inter3));
  inv1  gate1951(.a(s_201), .O(gate100inter4));
  nand2 gate1952(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1953(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1954(.a(G31), .O(gate100inter7));
  inv1  gate1955(.a(G353), .O(gate100inter8));
  nand2 gate1956(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1957(.a(s_201), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1958(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1959(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1960(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate2269(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2270(.a(gate103inter0), .b(s_246), .O(gate103inter1));
  and2  gate2271(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2272(.a(s_246), .O(gate103inter3));
  inv1  gate2273(.a(s_247), .O(gate103inter4));
  nand2 gate2274(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2275(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2276(.a(G28), .O(gate103inter7));
  inv1  gate2277(.a(G359), .O(gate103inter8));
  nand2 gate2278(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2279(.a(s_247), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2280(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2281(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2282(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1247(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1248(.a(gate104inter0), .b(s_100), .O(gate104inter1));
  and2  gate1249(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1250(.a(s_100), .O(gate104inter3));
  inv1  gate1251(.a(s_101), .O(gate104inter4));
  nand2 gate1252(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1253(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1254(.a(G32), .O(gate104inter7));
  inv1  gate1255(.a(G359), .O(gate104inter8));
  nand2 gate1256(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1257(.a(s_101), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1258(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1259(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1260(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate547(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate548(.a(gate107inter0), .b(s_0), .O(gate107inter1));
  and2  gate549(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate550(.a(s_0), .O(gate107inter3));
  inv1  gate551(.a(s_1), .O(gate107inter4));
  nand2 gate552(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate553(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate554(.a(G366), .O(gate107inter7));
  inv1  gate555(.a(G367), .O(gate107inter8));
  nand2 gate556(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate557(.a(s_1), .b(gate107inter3), .O(gate107inter10));
  nor2  gate558(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate559(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate560(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1933(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1934(.a(gate110inter0), .b(s_198), .O(gate110inter1));
  and2  gate1935(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1936(.a(s_198), .O(gate110inter3));
  inv1  gate1937(.a(s_199), .O(gate110inter4));
  nand2 gate1938(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1939(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1940(.a(G372), .O(gate110inter7));
  inv1  gate1941(.a(G373), .O(gate110inter8));
  nand2 gate1942(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1943(.a(s_199), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1944(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1945(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1946(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2367(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2368(.a(gate111inter0), .b(s_260), .O(gate111inter1));
  and2  gate2369(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2370(.a(s_260), .O(gate111inter3));
  inv1  gate2371(.a(s_261), .O(gate111inter4));
  nand2 gate2372(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2373(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2374(.a(G374), .O(gate111inter7));
  inv1  gate2375(.a(G375), .O(gate111inter8));
  nand2 gate2376(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2377(.a(s_261), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2378(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2379(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2380(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2927(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2928(.a(gate115inter0), .b(s_340), .O(gate115inter1));
  and2  gate2929(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2930(.a(s_340), .O(gate115inter3));
  inv1  gate2931(.a(s_341), .O(gate115inter4));
  nand2 gate2932(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2933(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2934(.a(G382), .O(gate115inter7));
  inv1  gate2935(.a(G383), .O(gate115inter8));
  nand2 gate2936(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2937(.a(s_341), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2938(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2939(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2940(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1975(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1976(.a(gate121inter0), .b(s_204), .O(gate121inter1));
  and2  gate1977(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1978(.a(s_204), .O(gate121inter3));
  inv1  gate1979(.a(s_205), .O(gate121inter4));
  nand2 gate1980(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1981(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1982(.a(G394), .O(gate121inter7));
  inv1  gate1983(.a(G395), .O(gate121inter8));
  nand2 gate1984(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1985(.a(s_205), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1986(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1987(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1988(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1709(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1710(.a(gate124inter0), .b(s_166), .O(gate124inter1));
  and2  gate1711(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1712(.a(s_166), .O(gate124inter3));
  inv1  gate1713(.a(s_167), .O(gate124inter4));
  nand2 gate1714(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1715(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1716(.a(G400), .O(gate124inter7));
  inv1  gate1717(.a(G401), .O(gate124inter8));
  nand2 gate1718(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1719(.a(s_167), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1720(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1721(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1722(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1415(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1416(.a(gate131inter0), .b(s_124), .O(gate131inter1));
  and2  gate1417(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1418(.a(s_124), .O(gate131inter3));
  inv1  gate1419(.a(s_125), .O(gate131inter4));
  nand2 gate1420(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1421(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1422(.a(G414), .O(gate131inter7));
  inv1  gate1423(.a(G415), .O(gate131inter8));
  nand2 gate1424(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1425(.a(s_125), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1426(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1427(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1428(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate771(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate772(.a(gate132inter0), .b(s_32), .O(gate132inter1));
  and2  gate773(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate774(.a(s_32), .O(gate132inter3));
  inv1  gate775(.a(s_33), .O(gate132inter4));
  nand2 gate776(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate777(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate778(.a(G416), .O(gate132inter7));
  inv1  gate779(.a(G417), .O(gate132inter8));
  nand2 gate780(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate781(.a(s_33), .b(gate132inter3), .O(gate132inter10));
  nor2  gate782(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate783(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate784(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2591(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2592(.a(gate133inter0), .b(s_292), .O(gate133inter1));
  and2  gate2593(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2594(.a(s_292), .O(gate133inter3));
  inv1  gate2595(.a(s_293), .O(gate133inter4));
  nand2 gate2596(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2597(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2598(.a(G418), .O(gate133inter7));
  inv1  gate2599(.a(G419), .O(gate133inter8));
  nand2 gate2600(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2601(.a(s_293), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2602(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2603(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2604(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1303(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1304(.a(gate136inter0), .b(s_108), .O(gate136inter1));
  and2  gate1305(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1306(.a(s_108), .O(gate136inter3));
  inv1  gate1307(.a(s_109), .O(gate136inter4));
  nand2 gate1308(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1309(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1310(.a(G424), .O(gate136inter7));
  inv1  gate1311(.a(G425), .O(gate136inter8));
  nand2 gate1312(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1313(.a(s_109), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1314(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1315(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1316(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2045(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2046(.a(gate137inter0), .b(s_214), .O(gate137inter1));
  and2  gate2047(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2048(.a(s_214), .O(gate137inter3));
  inv1  gate2049(.a(s_215), .O(gate137inter4));
  nand2 gate2050(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2051(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2052(.a(G426), .O(gate137inter7));
  inv1  gate2053(.a(G429), .O(gate137inter8));
  nand2 gate2054(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2055(.a(s_215), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2056(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2057(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2058(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate631(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate632(.a(gate138inter0), .b(s_12), .O(gate138inter1));
  and2  gate633(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate634(.a(s_12), .O(gate138inter3));
  inv1  gate635(.a(s_13), .O(gate138inter4));
  nand2 gate636(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate637(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate638(.a(G432), .O(gate138inter7));
  inv1  gate639(.a(G435), .O(gate138inter8));
  nand2 gate640(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate641(.a(s_13), .b(gate138inter3), .O(gate138inter10));
  nor2  gate642(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate643(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate644(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2185(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2186(.a(gate144inter0), .b(s_234), .O(gate144inter1));
  and2  gate2187(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2188(.a(s_234), .O(gate144inter3));
  inv1  gate2189(.a(s_235), .O(gate144inter4));
  nand2 gate2190(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2191(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2192(.a(G468), .O(gate144inter7));
  inv1  gate2193(.a(G471), .O(gate144inter8));
  nand2 gate2194(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2195(.a(s_235), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2196(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2197(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2198(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate645(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate646(.a(gate145inter0), .b(s_14), .O(gate145inter1));
  and2  gate647(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate648(.a(s_14), .O(gate145inter3));
  inv1  gate649(.a(s_15), .O(gate145inter4));
  nand2 gate650(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate651(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate652(.a(G474), .O(gate145inter7));
  inv1  gate653(.a(G477), .O(gate145inter8));
  nand2 gate654(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate655(.a(s_15), .b(gate145inter3), .O(gate145inter10));
  nor2  gate656(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate657(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate658(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1065(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1066(.a(gate147inter0), .b(s_74), .O(gate147inter1));
  and2  gate1067(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1068(.a(s_74), .O(gate147inter3));
  inv1  gate1069(.a(s_75), .O(gate147inter4));
  nand2 gate1070(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1071(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1072(.a(G486), .O(gate147inter7));
  inv1  gate1073(.a(G489), .O(gate147inter8));
  nand2 gate1074(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1075(.a(s_75), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1076(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1077(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1078(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2913(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2914(.a(gate149inter0), .b(s_338), .O(gate149inter1));
  and2  gate2915(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2916(.a(s_338), .O(gate149inter3));
  inv1  gate2917(.a(s_339), .O(gate149inter4));
  nand2 gate2918(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2919(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2920(.a(G498), .O(gate149inter7));
  inv1  gate2921(.a(G501), .O(gate149inter8));
  nand2 gate2922(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2923(.a(s_339), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2924(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2925(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2926(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2031(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2032(.a(gate150inter0), .b(s_212), .O(gate150inter1));
  and2  gate2033(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2034(.a(s_212), .O(gate150inter3));
  inv1  gate2035(.a(s_213), .O(gate150inter4));
  nand2 gate2036(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2037(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2038(.a(G504), .O(gate150inter7));
  inv1  gate2039(.a(G507), .O(gate150inter8));
  nand2 gate2040(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2041(.a(s_213), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2042(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2043(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2044(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2493(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2494(.a(gate152inter0), .b(s_278), .O(gate152inter1));
  and2  gate2495(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2496(.a(s_278), .O(gate152inter3));
  inv1  gate2497(.a(s_279), .O(gate152inter4));
  nand2 gate2498(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2499(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2500(.a(G516), .O(gate152inter7));
  inv1  gate2501(.a(G519), .O(gate152inter8));
  nand2 gate2502(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2503(.a(s_279), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2504(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2505(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2506(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate3067(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate3068(.a(gate154inter0), .b(s_360), .O(gate154inter1));
  and2  gate3069(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate3070(.a(s_360), .O(gate154inter3));
  inv1  gate3071(.a(s_361), .O(gate154inter4));
  nand2 gate3072(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate3073(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate3074(.a(G429), .O(gate154inter7));
  inv1  gate3075(.a(G522), .O(gate154inter8));
  nand2 gate3076(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate3077(.a(s_361), .b(gate154inter3), .O(gate154inter10));
  nor2  gate3078(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate3079(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate3080(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1009(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1010(.a(gate155inter0), .b(s_66), .O(gate155inter1));
  and2  gate1011(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1012(.a(s_66), .O(gate155inter3));
  inv1  gate1013(.a(s_67), .O(gate155inter4));
  nand2 gate1014(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1015(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1016(.a(G432), .O(gate155inter7));
  inv1  gate1017(.a(G525), .O(gate155inter8));
  nand2 gate1018(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1019(.a(s_67), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1020(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1021(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1022(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate841(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate842(.a(gate156inter0), .b(s_42), .O(gate156inter1));
  and2  gate843(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate844(.a(s_42), .O(gate156inter3));
  inv1  gate845(.a(s_43), .O(gate156inter4));
  nand2 gate846(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate847(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate848(.a(G435), .O(gate156inter7));
  inv1  gate849(.a(G525), .O(gate156inter8));
  nand2 gate850(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate851(.a(s_43), .b(gate156inter3), .O(gate156inter10));
  nor2  gate852(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate853(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate854(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1149(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1150(.a(gate160inter0), .b(s_86), .O(gate160inter1));
  and2  gate1151(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1152(.a(s_86), .O(gate160inter3));
  inv1  gate1153(.a(s_87), .O(gate160inter4));
  nand2 gate1154(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1155(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1156(.a(G447), .O(gate160inter7));
  inv1  gate1157(.a(G531), .O(gate160inter8));
  nand2 gate1158(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1159(.a(s_87), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1160(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1161(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1162(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2703(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2704(.a(gate162inter0), .b(s_308), .O(gate162inter1));
  and2  gate2705(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2706(.a(s_308), .O(gate162inter3));
  inv1  gate2707(.a(s_309), .O(gate162inter4));
  nand2 gate2708(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2709(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2710(.a(G453), .O(gate162inter7));
  inv1  gate2711(.a(G534), .O(gate162inter8));
  nand2 gate2712(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2713(.a(s_309), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2714(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2715(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2716(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate967(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate968(.a(gate165inter0), .b(s_60), .O(gate165inter1));
  and2  gate969(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate970(.a(s_60), .O(gate165inter3));
  inv1  gate971(.a(s_61), .O(gate165inter4));
  nand2 gate972(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate973(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate974(.a(G462), .O(gate165inter7));
  inv1  gate975(.a(G540), .O(gate165inter8));
  nand2 gate976(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate977(.a(s_61), .b(gate165inter3), .O(gate165inter10));
  nor2  gate978(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate979(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate980(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2465(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2466(.a(gate167inter0), .b(s_274), .O(gate167inter1));
  and2  gate2467(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2468(.a(s_274), .O(gate167inter3));
  inv1  gate2469(.a(s_275), .O(gate167inter4));
  nand2 gate2470(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2471(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2472(.a(G468), .O(gate167inter7));
  inv1  gate2473(.a(G543), .O(gate167inter8));
  nand2 gate2474(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2475(.a(s_275), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2476(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2477(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2478(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2451(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2452(.a(gate169inter0), .b(s_272), .O(gate169inter1));
  and2  gate2453(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2454(.a(s_272), .O(gate169inter3));
  inv1  gate2455(.a(s_273), .O(gate169inter4));
  nand2 gate2456(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2457(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2458(.a(G474), .O(gate169inter7));
  inv1  gate2459(.a(G546), .O(gate169inter8));
  nand2 gate2460(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2461(.a(s_273), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2462(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2463(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2464(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1233(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1234(.a(gate170inter0), .b(s_98), .O(gate170inter1));
  and2  gate1235(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1236(.a(s_98), .O(gate170inter3));
  inv1  gate1237(.a(s_99), .O(gate170inter4));
  nand2 gate1238(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1239(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1240(.a(G477), .O(gate170inter7));
  inv1  gate1241(.a(G546), .O(gate170inter8));
  nand2 gate1242(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1243(.a(s_99), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1244(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1245(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1246(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate939(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate940(.a(gate174inter0), .b(s_56), .O(gate174inter1));
  and2  gate941(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate942(.a(s_56), .O(gate174inter3));
  inv1  gate943(.a(s_57), .O(gate174inter4));
  nand2 gate944(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate945(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate946(.a(G489), .O(gate174inter7));
  inv1  gate947(.a(G552), .O(gate174inter8));
  nand2 gate948(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate949(.a(s_57), .b(gate174inter3), .O(gate174inter10));
  nor2  gate950(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate951(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate952(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate575(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate576(.a(gate180inter0), .b(s_4), .O(gate180inter1));
  and2  gate577(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate578(.a(s_4), .O(gate180inter3));
  inv1  gate579(.a(s_5), .O(gate180inter4));
  nand2 gate580(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate581(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate582(.a(G507), .O(gate180inter7));
  inv1  gate583(.a(G561), .O(gate180inter8));
  nand2 gate584(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate585(.a(s_5), .b(gate180inter3), .O(gate180inter10));
  nor2  gate586(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate587(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate588(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2955(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2956(.a(gate183inter0), .b(s_344), .O(gate183inter1));
  and2  gate2957(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2958(.a(s_344), .O(gate183inter3));
  inv1  gate2959(.a(s_345), .O(gate183inter4));
  nand2 gate2960(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2961(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2962(.a(G516), .O(gate183inter7));
  inv1  gate2963(.a(G567), .O(gate183inter8));
  nand2 gate2964(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2965(.a(s_345), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2966(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2967(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2968(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1261(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1262(.a(gate185inter0), .b(s_102), .O(gate185inter1));
  and2  gate1263(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1264(.a(s_102), .O(gate185inter3));
  inv1  gate1265(.a(s_103), .O(gate185inter4));
  nand2 gate1266(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1267(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1268(.a(G570), .O(gate185inter7));
  inv1  gate1269(.a(G571), .O(gate185inter8));
  nand2 gate1270(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1271(.a(s_103), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1272(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1273(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1274(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1919(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1920(.a(gate186inter0), .b(s_196), .O(gate186inter1));
  and2  gate1921(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1922(.a(s_196), .O(gate186inter3));
  inv1  gate1923(.a(s_197), .O(gate186inter4));
  nand2 gate1924(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1925(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1926(.a(G572), .O(gate186inter7));
  inv1  gate1927(.a(G573), .O(gate186inter8));
  nand2 gate1928(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1929(.a(s_197), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1930(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1931(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1932(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1219(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1220(.a(gate190inter0), .b(s_96), .O(gate190inter1));
  and2  gate1221(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1222(.a(s_96), .O(gate190inter3));
  inv1  gate1223(.a(s_97), .O(gate190inter4));
  nand2 gate1224(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1225(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1226(.a(G580), .O(gate190inter7));
  inv1  gate1227(.a(G581), .O(gate190inter8));
  nand2 gate1228(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1229(.a(s_97), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1230(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1231(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1232(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2815(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2816(.a(gate193inter0), .b(s_324), .O(gate193inter1));
  and2  gate2817(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2818(.a(s_324), .O(gate193inter3));
  inv1  gate2819(.a(s_325), .O(gate193inter4));
  nand2 gate2820(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2821(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2822(.a(G586), .O(gate193inter7));
  inv1  gate2823(.a(G587), .O(gate193inter8));
  nand2 gate2824(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2825(.a(s_325), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2826(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2827(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2828(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1877(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1878(.a(gate195inter0), .b(s_190), .O(gate195inter1));
  and2  gate1879(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1880(.a(s_190), .O(gate195inter3));
  inv1  gate1881(.a(s_191), .O(gate195inter4));
  nand2 gate1882(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1883(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1884(.a(G590), .O(gate195inter7));
  inv1  gate1885(.a(G591), .O(gate195inter8));
  nand2 gate1886(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1887(.a(s_191), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1888(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1889(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1890(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate897(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate898(.a(gate197inter0), .b(s_50), .O(gate197inter1));
  and2  gate899(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate900(.a(s_50), .O(gate197inter3));
  inv1  gate901(.a(s_51), .O(gate197inter4));
  nand2 gate902(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate903(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate904(.a(G594), .O(gate197inter7));
  inv1  gate905(.a(G595), .O(gate197inter8));
  nand2 gate906(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate907(.a(s_51), .b(gate197inter3), .O(gate197inter10));
  nor2  gate908(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate909(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate910(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate855(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate856(.a(gate200inter0), .b(s_44), .O(gate200inter1));
  and2  gate857(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate858(.a(s_44), .O(gate200inter3));
  inv1  gate859(.a(s_45), .O(gate200inter4));
  nand2 gate860(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate861(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate862(.a(G600), .O(gate200inter7));
  inv1  gate863(.a(G601), .O(gate200inter8));
  nand2 gate864(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate865(.a(s_45), .b(gate200inter3), .O(gate200inter10));
  nor2  gate866(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate867(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate868(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate2633(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2634(.a(gate201inter0), .b(s_298), .O(gate201inter1));
  and2  gate2635(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2636(.a(s_298), .O(gate201inter3));
  inv1  gate2637(.a(s_299), .O(gate201inter4));
  nand2 gate2638(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2639(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2640(.a(G602), .O(gate201inter7));
  inv1  gate2641(.a(G607), .O(gate201inter8));
  nand2 gate2642(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2643(.a(s_299), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2644(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2645(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2646(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate2311(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2312(.a(gate202inter0), .b(s_252), .O(gate202inter1));
  and2  gate2313(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2314(.a(s_252), .O(gate202inter3));
  inv1  gate2315(.a(s_253), .O(gate202inter4));
  nand2 gate2316(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2317(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2318(.a(G612), .O(gate202inter7));
  inv1  gate2319(.a(G617), .O(gate202inter8));
  nand2 gate2320(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2321(.a(s_253), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2322(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2323(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2324(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1387(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1388(.a(gate204inter0), .b(s_120), .O(gate204inter1));
  and2  gate1389(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1390(.a(s_120), .O(gate204inter3));
  inv1  gate1391(.a(s_121), .O(gate204inter4));
  nand2 gate1392(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1393(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1394(.a(G607), .O(gate204inter7));
  inv1  gate1395(.a(G617), .O(gate204inter8));
  nand2 gate1396(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1397(.a(s_121), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1398(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1399(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1400(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1373(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1374(.a(gate207inter0), .b(s_118), .O(gate207inter1));
  and2  gate1375(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1376(.a(s_118), .O(gate207inter3));
  inv1  gate1377(.a(s_119), .O(gate207inter4));
  nand2 gate1378(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1379(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1380(.a(G622), .O(gate207inter7));
  inv1  gate1381(.a(G632), .O(gate207inter8));
  nand2 gate1382(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1383(.a(s_119), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1384(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1385(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1386(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2283(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2284(.a(gate208inter0), .b(s_248), .O(gate208inter1));
  and2  gate2285(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2286(.a(s_248), .O(gate208inter3));
  inv1  gate2287(.a(s_249), .O(gate208inter4));
  nand2 gate2288(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2289(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2290(.a(G627), .O(gate208inter7));
  inv1  gate2291(.a(G637), .O(gate208inter8));
  nand2 gate2292(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2293(.a(s_249), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2294(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2295(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2296(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2199(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2200(.a(gate211inter0), .b(s_236), .O(gate211inter1));
  and2  gate2201(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2202(.a(s_236), .O(gate211inter3));
  inv1  gate2203(.a(s_237), .O(gate211inter4));
  nand2 gate2204(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2205(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2206(.a(G612), .O(gate211inter7));
  inv1  gate2207(.a(G669), .O(gate211inter8));
  nand2 gate2208(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2209(.a(s_237), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2210(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2211(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2212(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2717(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2718(.a(gate213inter0), .b(s_310), .O(gate213inter1));
  and2  gate2719(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2720(.a(s_310), .O(gate213inter3));
  inv1  gate2721(.a(s_311), .O(gate213inter4));
  nand2 gate2722(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2723(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2724(.a(G602), .O(gate213inter7));
  inv1  gate2725(.a(G672), .O(gate213inter8));
  nand2 gate2726(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2727(.a(s_311), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2728(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2729(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2730(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2339(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2340(.a(gate214inter0), .b(s_256), .O(gate214inter1));
  and2  gate2341(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2342(.a(s_256), .O(gate214inter3));
  inv1  gate2343(.a(s_257), .O(gate214inter4));
  nand2 gate2344(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2345(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2346(.a(G612), .O(gate214inter7));
  inv1  gate2347(.a(G672), .O(gate214inter8));
  nand2 gate2348(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2349(.a(s_257), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2350(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2351(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2352(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2619(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2620(.a(gate215inter0), .b(s_296), .O(gate215inter1));
  and2  gate2621(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2622(.a(s_296), .O(gate215inter3));
  inv1  gate2623(.a(s_297), .O(gate215inter4));
  nand2 gate2624(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2625(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2626(.a(G607), .O(gate215inter7));
  inv1  gate2627(.a(G675), .O(gate215inter8));
  nand2 gate2628(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2629(.a(s_297), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2630(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2631(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2632(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1569(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1570(.a(gate216inter0), .b(s_146), .O(gate216inter1));
  and2  gate1571(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1572(.a(s_146), .O(gate216inter3));
  inv1  gate1573(.a(s_147), .O(gate216inter4));
  nand2 gate1574(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1575(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1576(.a(G617), .O(gate216inter7));
  inv1  gate1577(.a(G675), .O(gate216inter8));
  nand2 gate1578(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1579(.a(s_147), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1580(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1581(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1582(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1191(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1192(.a(gate218inter0), .b(s_92), .O(gate218inter1));
  and2  gate1193(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1194(.a(s_92), .O(gate218inter3));
  inv1  gate1195(.a(s_93), .O(gate218inter4));
  nand2 gate1196(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1197(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1198(.a(G627), .O(gate218inter7));
  inv1  gate1199(.a(G678), .O(gate218inter8));
  nand2 gate1200(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1201(.a(s_93), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1202(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1203(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1204(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2143(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2144(.a(gate219inter0), .b(s_228), .O(gate219inter1));
  and2  gate2145(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2146(.a(s_228), .O(gate219inter3));
  inv1  gate2147(.a(s_229), .O(gate219inter4));
  nand2 gate2148(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2149(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2150(.a(G632), .O(gate219inter7));
  inv1  gate2151(.a(G681), .O(gate219inter8));
  nand2 gate2152(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2153(.a(s_229), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2154(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2155(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2156(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2745(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2746(.a(gate220inter0), .b(s_314), .O(gate220inter1));
  and2  gate2747(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2748(.a(s_314), .O(gate220inter3));
  inv1  gate2749(.a(s_315), .O(gate220inter4));
  nand2 gate2750(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2751(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2752(.a(G637), .O(gate220inter7));
  inv1  gate2753(.a(G681), .O(gate220inter8));
  nand2 gate2754(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2755(.a(s_315), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2756(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2757(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2758(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1667(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1668(.a(gate221inter0), .b(s_160), .O(gate221inter1));
  and2  gate1669(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1670(.a(s_160), .O(gate221inter3));
  inv1  gate1671(.a(s_161), .O(gate221inter4));
  nand2 gate1672(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1673(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1674(.a(G622), .O(gate221inter7));
  inv1  gate1675(.a(G684), .O(gate221inter8));
  nand2 gate1676(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1677(.a(s_161), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1678(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1679(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1680(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1163(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1164(.a(gate223inter0), .b(s_88), .O(gate223inter1));
  and2  gate1165(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1166(.a(s_88), .O(gate223inter3));
  inv1  gate1167(.a(s_89), .O(gate223inter4));
  nand2 gate1168(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1169(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1170(.a(G627), .O(gate223inter7));
  inv1  gate1171(.a(G687), .O(gate223inter8));
  nand2 gate1172(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1173(.a(s_89), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1174(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1175(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1176(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate3053(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate3054(.a(gate231inter0), .b(s_358), .O(gate231inter1));
  and2  gate3055(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate3056(.a(s_358), .O(gate231inter3));
  inv1  gate3057(.a(s_359), .O(gate231inter4));
  nand2 gate3058(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate3059(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate3060(.a(G702), .O(gate231inter7));
  inv1  gate3061(.a(G703), .O(gate231inter8));
  nand2 gate3062(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate3063(.a(s_359), .b(gate231inter3), .O(gate231inter10));
  nor2  gate3064(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate3065(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate3066(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2969(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2970(.a(gate234inter0), .b(s_346), .O(gate234inter1));
  and2  gate2971(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2972(.a(s_346), .O(gate234inter3));
  inv1  gate2973(.a(s_347), .O(gate234inter4));
  nand2 gate2974(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2975(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2976(.a(G245), .O(gate234inter7));
  inv1  gate2977(.a(G721), .O(gate234inter8));
  nand2 gate2978(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2979(.a(s_347), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2980(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2981(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2982(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate561(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate562(.a(gate237inter0), .b(s_2), .O(gate237inter1));
  and2  gate563(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate564(.a(s_2), .O(gate237inter3));
  inv1  gate565(.a(s_3), .O(gate237inter4));
  nand2 gate566(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate567(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate568(.a(G254), .O(gate237inter7));
  inv1  gate569(.a(G706), .O(gate237inter8));
  nand2 gate570(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate571(.a(s_3), .b(gate237inter3), .O(gate237inter10));
  nor2  gate572(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate573(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate574(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1177(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1178(.a(gate238inter0), .b(s_90), .O(gate238inter1));
  and2  gate1179(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1180(.a(s_90), .O(gate238inter3));
  inv1  gate1181(.a(s_91), .O(gate238inter4));
  nand2 gate1182(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1183(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1184(.a(G257), .O(gate238inter7));
  inv1  gate1185(.a(G709), .O(gate238inter8));
  nand2 gate1186(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1187(.a(s_91), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1188(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1189(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1190(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1961(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1962(.a(gate242inter0), .b(s_202), .O(gate242inter1));
  and2  gate1963(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1964(.a(s_202), .O(gate242inter3));
  inv1  gate1965(.a(s_203), .O(gate242inter4));
  nand2 gate1966(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1967(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1968(.a(G718), .O(gate242inter7));
  inv1  gate1969(.a(G730), .O(gate242inter8));
  nand2 gate1970(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1971(.a(s_203), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1972(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1973(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1974(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1107(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1108(.a(gate244inter0), .b(s_80), .O(gate244inter1));
  and2  gate1109(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1110(.a(s_80), .O(gate244inter3));
  inv1  gate1111(.a(s_81), .O(gate244inter4));
  nand2 gate1112(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1113(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1114(.a(G721), .O(gate244inter7));
  inv1  gate1115(.a(G733), .O(gate244inter8));
  nand2 gate1116(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1117(.a(s_81), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1118(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1119(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1120(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1499(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1500(.a(gate245inter0), .b(s_136), .O(gate245inter1));
  and2  gate1501(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1502(.a(s_136), .O(gate245inter3));
  inv1  gate1503(.a(s_137), .O(gate245inter4));
  nand2 gate1504(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1505(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1506(.a(G248), .O(gate245inter7));
  inv1  gate1507(.a(G736), .O(gate245inter8));
  nand2 gate1508(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1509(.a(s_137), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1510(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1511(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1512(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate673(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate674(.a(gate247inter0), .b(s_18), .O(gate247inter1));
  and2  gate675(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate676(.a(s_18), .O(gate247inter3));
  inv1  gate677(.a(s_19), .O(gate247inter4));
  nand2 gate678(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate679(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate680(.a(G251), .O(gate247inter7));
  inv1  gate681(.a(G739), .O(gate247inter8));
  nand2 gate682(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate683(.a(s_19), .b(gate247inter3), .O(gate247inter10));
  nor2  gate684(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate685(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate686(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2087(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2088(.a(gate248inter0), .b(s_220), .O(gate248inter1));
  and2  gate2089(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2090(.a(s_220), .O(gate248inter3));
  inv1  gate2091(.a(s_221), .O(gate248inter4));
  nand2 gate2092(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2093(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2094(.a(G727), .O(gate248inter7));
  inv1  gate2095(.a(G739), .O(gate248inter8));
  nand2 gate2096(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2097(.a(s_221), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2098(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2099(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2100(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2017(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2018(.a(gate249inter0), .b(s_210), .O(gate249inter1));
  and2  gate2019(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2020(.a(s_210), .O(gate249inter3));
  inv1  gate2021(.a(s_211), .O(gate249inter4));
  nand2 gate2022(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2023(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2024(.a(G254), .O(gate249inter7));
  inv1  gate2025(.a(G742), .O(gate249inter8));
  nand2 gate2026(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2027(.a(s_211), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2028(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2029(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2030(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1779(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1780(.a(gate252inter0), .b(s_176), .O(gate252inter1));
  and2  gate1781(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1782(.a(s_176), .O(gate252inter3));
  inv1  gate1783(.a(s_177), .O(gate252inter4));
  nand2 gate1784(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1785(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1786(.a(G709), .O(gate252inter7));
  inv1  gate1787(.a(G745), .O(gate252inter8));
  nand2 gate1788(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1789(.a(s_177), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1790(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1791(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1792(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2787(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2788(.a(gate256inter0), .b(s_320), .O(gate256inter1));
  and2  gate2789(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2790(.a(s_320), .O(gate256inter3));
  inv1  gate2791(.a(s_321), .O(gate256inter4));
  nand2 gate2792(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2793(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2794(.a(G715), .O(gate256inter7));
  inv1  gate2795(.a(G751), .O(gate256inter8));
  nand2 gate2796(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2797(.a(s_321), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2798(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2799(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2800(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2661(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2662(.a(gate258inter0), .b(s_302), .O(gate258inter1));
  and2  gate2663(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2664(.a(s_302), .O(gate258inter3));
  inv1  gate2665(.a(s_303), .O(gate258inter4));
  nand2 gate2666(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2667(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2668(.a(G756), .O(gate258inter7));
  inv1  gate2669(.a(G757), .O(gate258inter8));
  nand2 gate2670(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2671(.a(s_303), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2672(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2673(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2674(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1471(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1472(.a(gate260inter0), .b(s_132), .O(gate260inter1));
  and2  gate1473(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1474(.a(s_132), .O(gate260inter3));
  inv1  gate1475(.a(s_133), .O(gate260inter4));
  nand2 gate1476(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1477(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1478(.a(G760), .O(gate260inter7));
  inv1  gate1479(.a(G761), .O(gate260inter8));
  nand2 gate1480(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1481(.a(s_133), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1482(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1483(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1484(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2059(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2060(.a(gate263inter0), .b(s_216), .O(gate263inter1));
  and2  gate2061(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2062(.a(s_216), .O(gate263inter3));
  inv1  gate2063(.a(s_217), .O(gate263inter4));
  nand2 gate2064(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2065(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2066(.a(G766), .O(gate263inter7));
  inv1  gate2067(.a(G767), .O(gate263inter8));
  nand2 gate2068(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2069(.a(s_217), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2070(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2071(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2072(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1317(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1318(.a(gate264inter0), .b(s_110), .O(gate264inter1));
  and2  gate1319(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1320(.a(s_110), .O(gate264inter3));
  inv1  gate1321(.a(s_111), .O(gate264inter4));
  nand2 gate1322(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1323(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1324(.a(G768), .O(gate264inter7));
  inv1  gate1325(.a(G769), .O(gate264inter8));
  nand2 gate1326(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1327(.a(s_111), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1328(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1329(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1330(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate2157(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2158(.a(gate265inter0), .b(s_230), .O(gate265inter1));
  and2  gate2159(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2160(.a(s_230), .O(gate265inter3));
  inv1  gate2161(.a(s_231), .O(gate265inter4));
  nand2 gate2162(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2163(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2164(.a(G642), .O(gate265inter7));
  inv1  gate2165(.a(G770), .O(gate265inter8));
  nand2 gate2166(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2167(.a(s_231), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2168(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2169(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2170(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate2255(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2256(.a(gate266inter0), .b(s_244), .O(gate266inter1));
  and2  gate2257(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2258(.a(s_244), .O(gate266inter3));
  inv1  gate2259(.a(s_245), .O(gate266inter4));
  nand2 gate2260(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2261(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2262(.a(G645), .O(gate266inter7));
  inv1  gate2263(.a(G773), .O(gate266inter8));
  nand2 gate2264(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2265(.a(s_245), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2266(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2267(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2268(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1891(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1892(.a(gate267inter0), .b(s_192), .O(gate267inter1));
  and2  gate1893(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1894(.a(s_192), .O(gate267inter3));
  inv1  gate1895(.a(s_193), .O(gate267inter4));
  nand2 gate1896(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1897(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1898(.a(G648), .O(gate267inter7));
  inv1  gate1899(.a(G776), .O(gate267inter8));
  nand2 gate1900(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1901(.a(s_193), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1902(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1903(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1904(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1625(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1626(.a(gate268inter0), .b(s_154), .O(gate268inter1));
  and2  gate1627(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1628(.a(s_154), .O(gate268inter3));
  inv1  gate1629(.a(s_155), .O(gate268inter4));
  nand2 gate1630(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1631(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1632(.a(G651), .O(gate268inter7));
  inv1  gate1633(.a(G779), .O(gate268inter8));
  nand2 gate1634(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1635(.a(s_155), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1636(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1637(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1638(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate701(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate702(.a(gate272inter0), .b(s_22), .O(gate272inter1));
  and2  gate703(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate704(.a(s_22), .O(gate272inter3));
  inv1  gate705(.a(s_23), .O(gate272inter4));
  nand2 gate706(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate707(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate708(.a(G663), .O(gate272inter7));
  inv1  gate709(.a(G791), .O(gate272inter8));
  nand2 gate710(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate711(.a(s_23), .b(gate272inter3), .O(gate272inter10));
  nor2  gate712(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate713(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate714(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate3011(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate3012(.a(gate273inter0), .b(s_352), .O(gate273inter1));
  and2  gate3013(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate3014(.a(s_352), .O(gate273inter3));
  inv1  gate3015(.a(s_353), .O(gate273inter4));
  nand2 gate3016(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate3017(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate3018(.a(G642), .O(gate273inter7));
  inv1  gate3019(.a(G794), .O(gate273inter8));
  nand2 gate3020(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate3021(.a(s_353), .b(gate273inter3), .O(gate273inter10));
  nor2  gate3022(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate3023(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate3024(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2003(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2004(.a(gate274inter0), .b(s_208), .O(gate274inter1));
  and2  gate2005(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2006(.a(s_208), .O(gate274inter3));
  inv1  gate2007(.a(s_209), .O(gate274inter4));
  nand2 gate2008(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2009(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2010(.a(G770), .O(gate274inter7));
  inv1  gate2011(.a(G794), .O(gate274inter8));
  nand2 gate2012(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2013(.a(s_209), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2014(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2015(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2016(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1737(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1738(.a(gate275inter0), .b(s_170), .O(gate275inter1));
  and2  gate1739(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1740(.a(s_170), .O(gate275inter3));
  inv1  gate1741(.a(s_171), .O(gate275inter4));
  nand2 gate1742(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1743(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1744(.a(G645), .O(gate275inter7));
  inv1  gate1745(.a(G797), .O(gate275inter8));
  nand2 gate1746(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1747(.a(s_171), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1748(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1749(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1750(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2101(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2102(.a(gate277inter0), .b(s_222), .O(gate277inter1));
  and2  gate2103(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2104(.a(s_222), .O(gate277inter3));
  inv1  gate2105(.a(s_223), .O(gate277inter4));
  nand2 gate2106(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2107(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2108(.a(G648), .O(gate277inter7));
  inv1  gate2109(.a(G800), .O(gate277inter8));
  nand2 gate2110(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2111(.a(s_223), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2112(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2113(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2114(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate687(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate688(.a(gate278inter0), .b(s_20), .O(gate278inter1));
  and2  gate689(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate690(.a(s_20), .O(gate278inter3));
  inv1  gate691(.a(s_21), .O(gate278inter4));
  nand2 gate692(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate693(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate694(.a(G776), .O(gate278inter7));
  inv1  gate695(.a(G800), .O(gate278inter8));
  nand2 gate696(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate697(.a(s_21), .b(gate278inter3), .O(gate278inter10));
  nor2  gate698(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate699(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate700(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1849(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1850(.a(gate279inter0), .b(s_186), .O(gate279inter1));
  and2  gate1851(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1852(.a(s_186), .O(gate279inter3));
  inv1  gate1853(.a(s_187), .O(gate279inter4));
  nand2 gate1854(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1855(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1856(.a(G651), .O(gate279inter7));
  inv1  gate1857(.a(G803), .O(gate279inter8));
  nand2 gate1858(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1859(.a(s_187), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1860(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1861(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1862(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate995(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate996(.a(gate280inter0), .b(s_64), .O(gate280inter1));
  and2  gate997(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate998(.a(s_64), .O(gate280inter3));
  inv1  gate999(.a(s_65), .O(gate280inter4));
  nand2 gate1000(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1001(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1002(.a(G779), .O(gate280inter7));
  inv1  gate1003(.a(G803), .O(gate280inter8));
  nand2 gate1004(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1005(.a(s_65), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1006(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1007(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1008(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1723(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1724(.a(gate282inter0), .b(s_168), .O(gate282inter1));
  and2  gate1725(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1726(.a(s_168), .O(gate282inter3));
  inv1  gate1727(.a(s_169), .O(gate282inter4));
  nand2 gate1728(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1729(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1730(.a(G782), .O(gate282inter7));
  inv1  gate1731(.a(G806), .O(gate282inter8));
  nand2 gate1732(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1733(.a(s_169), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1734(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1735(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1736(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2213(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2214(.a(gate283inter0), .b(s_238), .O(gate283inter1));
  and2  gate2215(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2216(.a(s_238), .O(gate283inter3));
  inv1  gate2217(.a(s_239), .O(gate283inter4));
  nand2 gate2218(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2219(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2220(.a(G657), .O(gate283inter7));
  inv1  gate2221(.a(G809), .O(gate283inter8));
  nand2 gate2222(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2223(.a(s_239), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2224(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2225(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2226(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2885(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2886(.a(gate285inter0), .b(s_334), .O(gate285inter1));
  and2  gate2887(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2888(.a(s_334), .O(gate285inter3));
  inv1  gate2889(.a(s_335), .O(gate285inter4));
  nand2 gate2890(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2891(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2892(.a(G660), .O(gate285inter7));
  inv1  gate2893(.a(G812), .O(gate285inter8));
  nand2 gate2894(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2895(.a(s_335), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2896(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2897(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2898(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1611(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1612(.a(gate288inter0), .b(s_152), .O(gate288inter1));
  and2  gate1613(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1614(.a(s_152), .O(gate288inter3));
  inv1  gate1615(.a(s_153), .O(gate288inter4));
  nand2 gate1616(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1617(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1618(.a(G791), .O(gate288inter7));
  inv1  gate1619(.a(G815), .O(gate288inter8));
  nand2 gate1620(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1621(.a(s_153), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1622(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1623(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1624(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1541(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1542(.a(gate289inter0), .b(s_142), .O(gate289inter1));
  and2  gate1543(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1544(.a(s_142), .O(gate289inter3));
  inv1  gate1545(.a(s_143), .O(gate289inter4));
  nand2 gate1546(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1547(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1548(.a(G818), .O(gate289inter7));
  inv1  gate1549(.a(G819), .O(gate289inter8));
  nand2 gate1550(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1551(.a(s_143), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1552(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1553(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1554(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate869(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate870(.a(gate291inter0), .b(s_46), .O(gate291inter1));
  and2  gate871(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate872(.a(s_46), .O(gate291inter3));
  inv1  gate873(.a(s_47), .O(gate291inter4));
  nand2 gate874(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate875(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate876(.a(G822), .O(gate291inter7));
  inv1  gate877(.a(G823), .O(gate291inter8));
  nand2 gate878(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate879(.a(s_47), .b(gate291inter3), .O(gate291inter10));
  nor2  gate880(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate881(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate882(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1653(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1654(.a(gate294inter0), .b(s_158), .O(gate294inter1));
  and2  gate1655(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1656(.a(s_158), .O(gate294inter3));
  inv1  gate1657(.a(s_159), .O(gate294inter4));
  nand2 gate1658(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1659(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1660(.a(G832), .O(gate294inter7));
  inv1  gate1661(.a(G833), .O(gate294inter8));
  nand2 gate1662(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1663(.a(s_159), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1664(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1665(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1666(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1793(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1794(.a(gate388inter0), .b(s_178), .O(gate388inter1));
  and2  gate1795(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1796(.a(s_178), .O(gate388inter3));
  inv1  gate1797(.a(s_179), .O(gate388inter4));
  nand2 gate1798(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1799(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1800(.a(G2), .O(gate388inter7));
  inv1  gate1801(.a(G1039), .O(gate388inter8));
  nand2 gate1802(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1803(.a(s_179), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1804(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1805(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1806(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1359(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1360(.a(gate395inter0), .b(s_116), .O(gate395inter1));
  and2  gate1361(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1362(.a(s_116), .O(gate395inter3));
  inv1  gate1363(.a(s_117), .O(gate395inter4));
  nand2 gate1364(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1365(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1366(.a(G9), .O(gate395inter7));
  inv1  gate1367(.a(G1060), .O(gate395inter8));
  nand2 gate1368(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1369(.a(s_117), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1370(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1371(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1372(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1695(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1696(.a(gate397inter0), .b(s_164), .O(gate397inter1));
  and2  gate1697(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1698(.a(s_164), .O(gate397inter3));
  inv1  gate1699(.a(s_165), .O(gate397inter4));
  nand2 gate1700(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1701(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1702(.a(G11), .O(gate397inter7));
  inv1  gate1703(.a(G1066), .O(gate397inter8));
  nand2 gate1704(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1705(.a(s_165), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1706(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1707(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1708(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1289(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1290(.a(gate398inter0), .b(s_106), .O(gate398inter1));
  and2  gate1291(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1292(.a(s_106), .O(gate398inter3));
  inv1  gate1293(.a(s_107), .O(gate398inter4));
  nand2 gate1294(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1295(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1296(.a(G12), .O(gate398inter7));
  inv1  gate1297(.a(G1069), .O(gate398inter8));
  nand2 gate1298(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1299(.a(s_107), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1300(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1301(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1302(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1135(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1136(.a(gate401inter0), .b(s_84), .O(gate401inter1));
  and2  gate1137(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1138(.a(s_84), .O(gate401inter3));
  inv1  gate1139(.a(s_85), .O(gate401inter4));
  nand2 gate1140(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1141(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1142(.a(G15), .O(gate401inter7));
  inv1  gate1143(.a(G1078), .O(gate401inter8));
  nand2 gate1144(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1145(.a(s_85), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1146(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1147(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1148(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2773(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2774(.a(gate404inter0), .b(s_318), .O(gate404inter1));
  and2  gate2775(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2776(.a(s_318), .O(gate404inter3));
  inv1  gate2777(.a(s_319), .O(gate404inter4));
  nand2 gate2778(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2779(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2780(.a(G18), .O(gate404inter7));
  inv1  gate2781(.a(G1087), .O(gate404inter8));
  nand2 gate2782(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2783(.a(s_319), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2784(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2785(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2786(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate813(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate814(.a(gate406inter0), .b(s_38), .O(gate406inter1));
  and2  gate815(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate816(.a(s_38), .O(gate406inter3));
  inv1  gate817(.a(s_39), .O(gate406inter4));
  nand2 gate818(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate819(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate820(.a(G20), .O(gate406inter7));
  inv1  gate821(.a(G1093), .O(gate406inter8));
  nand2 gate822(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate823(.a(s_39), .b(gate406inter3), .O(gate406inter10));
  nor2  gate824(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate825(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate826(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1275(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1276(.a(gate407inter0), .b(s_104), .O(gate407inter1));
  and2  gate1277(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1278(.a(s_104), .O(gate407inter3));
  inv1  gate1279(.a(s_105), .O(gate407inter4));
  nand2 gate1280(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1281(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1282(.a(G21), .O(gate407inter7));
  inv1  gate1283(.a(G1096), .O(gate407inter8));
  nand2 gate1284(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1285(.a(s_105), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1286(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1287(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1288(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2997(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2998(.a(gate417inter0), .b(s_350), .O(gate417inter1));
  and2  gate2999(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate3000(.a(s_350), .O(gate417inter3));
  inv1  gate3001(.a(s_351), .O(gate417inter4));
  nand2 gate3002(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate3003(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate3004(.a(G31), .O(gate417inter7));
  inv1  gate3005(.a(G1126), .O(gate417inter8));
  nand2 gate3006(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate3007(.a(s_351), .b(gate417inter3), .O(gate417inter10));
  nor2  gate3008(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate3009(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate3010(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1429(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1430(.a(gate420inter0), .b(s_126), .O(gate420inter1));
  and2  gate1431(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1432(.a(s_126), .O(gate420inter3));
  inv1  gate1433(.a(s_127), .O(gate420inter4));
  nand2 gate1434(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1435(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1436(.a(G1036), .O(gate420inter7));
  inv1  gate1437(.a(G1132), .O(gate420inter8));
  nand2 gate1438(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1439(.a(s_127), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1440(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1441(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1442(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate729(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate730(.a(gate422inter0), .b(s_26), .O(gate422inter1));
  and2  gate731(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate732(.a(s_26), .O(gate422inter3));
  inv1  gate733(.a(s_27), .O(gate422inter4));
  nand2 gate734(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate735(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate736(.a(G1039), .O(gate422inter7));
  inv1  gate737(.a(G1135), .O(gate422inter8));
  nand2 gate738(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate739(.a(s_27), .b(gate422inter3), .O(gate422inter10));
  nor2  gate740(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate741(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate742(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1023(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1024(.a(gate423inter0), .b(s_68), .O(gate423inter1));
  and2  gate1025(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1026(.a(s_68), .O(gate423inter3));
  inv1  gate1027(.a(s_69), .O(gate423inter4));
  nand2 gate1028(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1029(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1030(.a(G3), .O(gate423inter7));
  inv1  gate1031(.a(G1138), .O(gate423inter8));
  nand2 gate1032(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1033(.a(s_69), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1034(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1035(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1036(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2129(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2130(.a(gate424inter0), .b(s_226), .O(gate424inter1));
  and2  gate2131(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2132(.a(s_226), .O(gate424inter3));
  inv1  gate2133(.a(s_227), .O(gate424inter4));
  nand2 gate2134(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2135(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2136(.a(G1042), .O(gate424inter7));
  inv1  gate2137(.a(G1138), .O(gate424inter8));
  nand2 gate2138(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2139(.a(s_227), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2140(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2141(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2142(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1835(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1836(.a(gate425inter0), .b(s_184), .O(gate425inter1));
  and2  gate1837(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1838(.a(s_184), .O(gate425inter3));
  inv1  gate1839(.a(s_185), .O(gate425inter4));
  nand2 gate1840(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1841(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1842(.a(G4), .O(gate425inter7));
  inv1  gate1843(.a(G1141), .O(gate425inter8));
  nand2 gate1844(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1845(.a(s_185), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1846(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1847(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1848(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate659(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate660(.a(gate429inter0), .b(s_16), .O(gate429inter1));
  and2  gate661(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate662(.a(s_16), .O(gate429inter3));
  inv1  gate663(.a(s_17), .O(gate429inter4));
  nand2 gate664(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate665(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate666(.a(G6), .O(gate429inter7));
  inv1  gate667(.a(G1147), .O(gate429inter8));
  nand2 gate668(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate669(.a(s_17), .b(gate429inter3), .O(gate429inter10));
  nor2  gate670(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate671(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate672(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate2241(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2242(.a(gate430inter0), .b(s_242), .O(gate430inter1));
  and2  gate2243(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2244(.a(s_242), .O(gate430inter3));
  inv1  gate2245(.a(s_243), .O(gate430inter4));
  nand2 gate2246(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2247(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2248(.a(G1051), .O(gate430inter7));
  inv1  gate2249(.a(G1147), .O(gate430inter8));
  nand2 gate2250(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2251(.a(s_243), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2252(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2253(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2254(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1527(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1528(.a(gate431inter0), .b(s_140), .O(gate431inter1));
  and2  gate1529(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1530(.a(s_140), .O(gate431inter3));
  inv1  gate1531(.a(s_141), .O(gate431inter4));
  nand2 gate1532(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1533(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1534(.a(G7), .O(gate431inter7));
  inv1  gate1535(.a(G1150), .O(gate431inter8));
  nand2 gate1536(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1537(.a(s_141), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1538(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1539(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1540(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1345(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1346(.a(gate433inter0), .b(s_114), .O(gate433inter1));
  and2  gate1347(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1348(.a(s_114), .O(gate433inter3));
  inv1  gate1349(.a(s_115), .O(gate433inter4));
  nand2 gate1350(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1351(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1352(.a(G8), .O(gate433inter7));
  inv1  gate1353(.a(G1153), .O(gate433inter8));
  nand2 gate1354(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1355(.a(s_115), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1356(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1357(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1358(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2563(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2564(.a(gate435inter0), .b(s_288), .O(gate435inter1));
  and2  gate2565(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2566(.a(s_288), .O(gate435inter3));
  inv1  gate2567(.a(s_289), .O(gate435inter4));
  nand2 gate2568(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2569(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2570(.a(G9), .O(gate435inter7));
  inv1  gate2571(.a(G1156), .O(gate435inter8));
  nand2 gate2572(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2573(.a(s_289), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2574(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2575(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2576(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate2759(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2760(.a(gate436inter0), .b(s_316), .O(gate436inter1));
  and2  gate2761(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2762(.a(s_316), .O(gate436inter3));
  inv1  gate2763(.a(s_317), .O(gate436inter4));
  nand2 gate2764(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2765(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2766(.a(G1060), .O(gate436inter7));
  inv1  gate2767(.a(G1156), .O(gate436inter8));
  nand2 gate2768(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2769(.a(s_317), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2770(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2771(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2772(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1037(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1038(.a(gate437inter0), .b(s_70), .O(gate437inter1));
  and2  gate1039(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1040(.a(s_70), .O(gate437inter3));
  inv1  gate1041(.a(s_71), .O(gate437inter4));
  nand2 gate1042(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1043(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1044(.a(G10), .O(gate437inter7));
  inv1  gate1045(.a(G1159), .O(gate437inter8));
  nand2 gate1046(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1047(.a(s_71), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1048(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1049(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1050(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2395(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2396(.a(gate438inter0), .b(s_264), .O(gate438inter1));
  and2  gate2397(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2398(.a(s_264), .O(gate438inter3));
  inv1  gate2399(.a(s_265), .O(gate438inter4));
  nand2 gate2400(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2401(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2402(.a(G1063), .O(gate438inter7));
  inv1  gate2403(.a(G1159), .O(gate438inter8));
  nand2 gate2404(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2405(.a(s_265), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2406(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2407(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2408(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1583(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1584(.a(gate439inter0), .b(s_148), .O(gate439inter1));
  and2  gate1585(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1586(.a(s_148), .O(gate439inter3));
  inv1  gate1587(.a(s_149), .O(gate439inter4));
  nand2 gate1588(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1589(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1590(.a(G11), .O(gate439inter7));
  inv1  gate1591(.a(G1162), .O(gate439inter8));
  nand2 gate1592(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1593(.a(s_149), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1594(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1595(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1596(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate2437(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2438(.a(gate440inter0), .b(s_270), .O(gate440inter1));
  and2  gate2439(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2440(.a(s_270), .O(gate440inter3));
  inv1  gate2441(.a(s_271), .O(gate440inter4));
  nand2 gate2442(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2443(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2444(.a(G1066), .O(gate440inter7));
  inv1  gate2445(.a(G1162), .O(gate440inter8));
  nand2 gate2446(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2447(.a(s_271), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2448(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2449(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2450(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate981(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate982(.a(gate441inter0), .b(s_62), .O(gate441inter1));
  and2  gate983(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate984(.a(s_62), .O(gate441inter3));
  inv1  gate985(.a(s_63), .O(gate441inter4));
  nand2 gate986(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate987(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate988(.a(G12), .O(gate441inter7));
  inv1  gate989(.a(G1165), .O(gate441inter8));
  nand2 gate990(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate991(.a(s_63), .b(gate441inter3), .O(gate441inter10));
  nor2  gate992(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate993(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate994(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate589(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate590(.a(gate442inter0), .b(s_6), .O(gate442inter1));
  and2  gate591(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate592(.a(s_6), .O(gate442inter3));
  inv1  gate593(.a(s_7), .O(gate442inter4));
  nand2 gate594(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate595(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate596(.a(G1069), .O(gate442inter7));
  inv1  gate597(.a(G1165), .O(gate442inter8));
  nand2 gate598(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate599(.a(s_7), .b(gate442inter3), .O(gate442inter10));
  nor2  gate600(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate601(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate602(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate925(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate926(.a(gate444inter0), .b(s_54), .O(gate444inter1));
  and2  gate927(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate928(.a(s_54), .O(gate444inter3));
  inv1  gate929(.a(s_55), .O(gate444inter4));
  nand2 gate930(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate931(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate932(.a(G1072), .O(gate444inter7));
  inv1  gate933(.a(G1168), .O(gate444inter8));
  nand2 gate934(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate935(.a(s_55), .b(gate444inter3), .O(gate444inter10));
  nor2  gate936(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate937(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate938(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate911(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate912(.a(gate445inter0), .b(s_52), .O(gate445inter1));
  and2  gate913(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate914(.a(s_52), .O(gate445inter3));
  inv1  gate915(.a(s_53), .O(gate445inter4));
  nand2 gate916(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate917(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate918(.a(G14), .O(gate445inter7));
  inv1  gate919(.a(G1171), .O(gate445inter8));
  nand2 gate920(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate921(.a(s_53), .b(gate445inter3), .O(gate445inter10));
  nor2  gate922(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate923(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate924(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate715(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate716(.a(gate446inter0), .b(s_24), .O(gate446inter1));
  and2  gate717(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate718(.a(s_24), .O(gate446inter3));
  inv1  gate719(.a(s_25), .O(gate446inter4));
  nand2 gate720(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate721(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate722(.a(G1075), .O(gate446inter7));
  inv1  gate723(.a(G1171), .O(gate446inter8));
  nand2 gate724(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate725(.a(s_25), .b(gate446inter3), .O(gate446inter10));
  nor2  gate726(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate727(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate728(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2605(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2606(.a(gate447inter0), .b(s_294), .O(gate447inter1));
  and2  gate2607(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2608(.a(s_294), .O(gate447inter3));
  inv1  gate2609(.a(s_295), .O(gate447inter4));
  nand2 gate2610(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2611(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2612(.a(G15), .O(gate447inter7));
  inv1  gate2613(.a(G1174), .O(gate447inter8));
  nand2 gate2614(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2615(.a(s_295), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2616(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2617(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2618(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2675(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2676(.a(gate448inter0), .b(s_304), .O(gate448inter1));
  and2  gate2677(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2678(.a(s_304), .O(gate448inter3));
  inv1  gate2679(.a(s_305), .O(gate448inter4));
  nand2 gate2680(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2681(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2682(.a(G1078), .O(gate448inter7));
  inv1  gate2683(.a(G1174), .O(gate448inter8));
  nand2 gate2684(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2685(.a(s_305), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2686(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2687(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2688(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1331(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1332(.a(gate449inter0), .b(s_112), .O(gate449inter1));
  and2  gate1333(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1334(.a(s_112), .O(gate449inter3));
  inv1  gate1335(.a(s_113), .O(gate449inter4));
  nand2 gate1336(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1337(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1338(.a(G16), .O(gate449inter7));
  inv1  gate1339(.a(G1177), .O(gate449inter8));
  nand2 gate1340(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1341(.a(s_113), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1342(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1343(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1344(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1513(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1514(.a(gate450inter0), .b(s_138), .O(gate450inter1));
  and2  gate1515(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1516(.a(s_138), .O(gate450inter3));
  inv1  gate1517(.a(s_139), .O(gate450inter4));
  nand2 gate1518(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1519(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1520(.a(G1081), .O(gate450inter7));
  inv1  gate1521(.a(G1177), .O(gate450inter8));
  nand2 gate1522(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1523(.a(s_139), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1524(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1525(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1526(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate757(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate758(.a(gate453inter0), .b(s_30), .O(gate453inter1));
  and2  gate759(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate760(.a(s_30), .O(gate453inter3));
  inv1  gate761(.a(s_31), .O(gate453inter4));
  nand2 gate762(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate763(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate764(.a(G18), .O(gate453inter7));
  inv1  gate765(.a(G1183), .O(gate453inter8));
  nand2 gate766(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate767(.a(s_31), .b(gate453inter3), .O(gate453inter10));
  nor2  gate768(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate769(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate770(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate603(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate604(.a(gate454inter0), .b(s_8), .O(gate454inter1));
  and2  gate605(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate606(.a(s_8), .O(gate454inter3));
  inv1  gate607(.a(s_9), .O(gate454inter4));
  nand2 gate608(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate609(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate610(.a(G1087), .O(gate454inter7));
  inv1  gate611(.a(G1183), .O(gate454inter8));
  nand2 gate612(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate613(.a(s_9), .b(gate454inter3), .O(gate454inter10));
  nor2  gate614(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate615(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate616(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1807(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1808(.a(gate456inter0), .b(s_180), .O(gate456inter1));
  and2  gate1809(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1810(.a(s_180), .O(gate456inter3));
  inv1  gate1811(.a(s_181), .O(gate456inter4));
  nand2 gate1812(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1813(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1814(.a(G1090), .O(gate456inter7));
  inv1  gate1815(.a(G1186), .O(gate456inter8));
  nand2 gate1816(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1817(.a(s_181), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1818(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1819(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1820(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate883(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate884(.a(gate463inter0), .b(s_48), .O(gate463inter1));
  and2  gate885(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate886(.a(s_48), .O(gate463inter3));
  inv1  gate887(.a(s_49), .O(gate463inter4));
  nand2 gate888(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate889(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate890(.a(G23), .O(gate463inter7));
  inv1  gate891(.a(G1198), .O(gate463inter8));
  nand2 gate892(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate893(.a(s_49), .b(gate463inter3), .O(gate463inter10));
  nor2  gate894(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate895(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate896(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate799(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate800(.a(gate464inter0), .b(s_36), .O(gate464inter1));
  and2  gate801(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate802(.a(s_36), .O(gate464inter3));
  inv1  gate803(.a(s_37), .O(gate464inter4));
  nand2 gate804(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate805(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate806(.a(G1102), .O(gate464inter7));
  inv1  gate807(.a(G1198), .O(gate464inter8));
  nand2 gate808(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate809(.a(s_37), .b(gate464inter3), .O(gate464inter10));
  nor2  gate810(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate811(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate812(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate3039(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate3040(.a(gate466inter0), .b(s_356), .O(gate466inter1));
  and2  gate3041(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate3042(.a(s_356), .O(gate466inter3));
  inv1  gate3043(.a(s_357), .O(gate466inter4));
  nand2 gate3044(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate3045(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate3046(.a(G1105), .O(gate466inter7));
  inv1  gate3047(.a(G1201), .O(gate466inter8));
  nand2 gate3048(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate3049(.a(s_357), .b(gate466inter3), .O(gate466inter10));
  nor2  gate3050(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate3051(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate3052(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1765(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1766(.a(gate471inter0), .b(s_174), .O(gate471inter1));
  and2  gate1767(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1768(.a(s_174), .O(gate471inter3));
  inv1  gate1769(.a(s_175), .O(gate471inter4));
  nand2 gate1770(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1771(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1772(.a(G27), .O(gate471inter7));
  inv1  gate1773(.a(G1210), .O(gate471inter8));
  nand2 gate1774(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1775(.a(s_175), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1776(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1777(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1778(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2073(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2074(.a(gate474inter0), .b(s_218), .O(gate474inter1));
  and2  gate2075(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2076(.a(s_218), .O(gate474inter3));
  inv1  gate2077(.a(s_219), .O(gate474inter4));
  nand2 gate2078(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2079(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2080(.a(G1117), .O(gate474inter7));
  inv1  gate2081(.a(G1213), .O(gate474inter8));
  nand2 gate2082(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2083(.a(s_219), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2084(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2085(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2086(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate785(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate786(.a(gate476inter0), .b(s_34), .O(gate476inter1));
  and2  gate787(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate788(.a(s_34), .O(gate476inter3));
  inv1  gate789(.a(s_35), .O(gate476inter4));
  nand2 gate790(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate791(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate792(.a(G1120), .O(gate476inter7));
  inv1  gate793(.a(G1216), .O(gate476inter8));
  nand2 gate794(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate795(.a(s_35), .b(gate476inter3), .O(gate476inter10));
  nor2  gate796(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate797(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate798(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1905(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1906(.a(gate477inter0), .b(s_194), .O(gate477inter1));
  and2  gate1907(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1908(.a(s_194), .O(gate477inter3));
  inv1  gate1909(.a(s_195), .O(gate477inter4));
  nand2 gate1910(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1911(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1912(.a(G30), .O(gate477inter7));
  inv1  gate1913(.a(G1219), .O(gate477inter8));
  nand2 gate1914(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1915(.a(s_195), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1916(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1917(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1918(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2115(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2116(.a(gate479inter0), .b(s_224), .O(gate479inter1));
  and2  gate2117(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2118(.a(s_224), .O(gate479inter3));
  inv1  gate2119(.a(s_225), .O(gate479inter4));
  nand2 gate2120(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2121(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2122(.a(G31), .O(gate479inter7));
  inv1  gate2123(.a(G1222), .O(gate479inter8));
  nand2 gate2124(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2125(.a(s_225), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2126(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2127(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2128(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1401(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1402(.a(gate482inter0), .b(s_122), .O(gate482inter1));
  and2  gate1403(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1404(.a(s_122), .O(gate482inter3));
  inv1  gate1405(.a(s_123), .O(gate482inter4));
  nand2 gate1406(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1407(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1408(.a(G1129), .O(gate482inter7));
  inv1  gate1409(.a(G1225), .O(gate482inter8));
  nand2 gate1410(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1411(.a(s_123), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1412(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1413(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1414(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate2479(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2480(.a(gate484inter0), .b(s_276), .O(gate484inter1));
  and2  gate2481(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2482(.a(s_276), .O(gate484inter3));
  inv1  gate2483(.a(s_277), .O(gate484inter4));
  nand2 gate2484(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2485(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2486(.a(G1230), .O(gate484inter7));
  inv1  gate2487(.a(G1231), .O(gate484inter8));
  nand2 gate2488(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2489(.a(s_277), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2490(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2491(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2492(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1051(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1052(.a(gate488inter0), .b(s_72), .O(gate488inter1));
  and2  gate1053(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1054(.a(s_72), .O(gate488inter3));
  inv1  gate1055(.a(s_73), .O(gate488inter4));
  nand2 gate1056(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1057(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1058(.a(G1238), .O(gate488inter7));
  inv1  gate1059(.a(G1239), .O(gate488inter8));
  nand2 gate1060(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1061(.a(s_73), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1062(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1063(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1064(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1989(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1990(.a(gate489inter0), .b(s_206), .O(gate489inter1));
  and2  gate1991(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1992(.a(s_206), .O(gate489inter3));
  inv1  gate1993(.a(s_207), .O(gate489inter4));
  nand2 gate1994(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1995(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1996(.a(G1240), .O(gate489inter7));
  inv1  gate1997(.a(G1241), .O(gate489inter8));
  nand2 gate1998(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1999(.a(s_207), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2000(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2001(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2002(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1821(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1822(.a(gate490inter0), .b(s_182), .O(gate490inter1));
  and2  gate1823(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1824(.a(s_182), .O(gate490inter3));
  inv1  gate1825(.a(s_183), .O(gate490inter4));
  nand2 gate1826(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1827(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1828(.a(G1242), .O(gate490inter7));
  inv1  gate1829(.a(G1243), .O(gate490inter8));
  nand2 gate1830(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1831(.a(s_183), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1832(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1833(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1834(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate2871(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2872(.a(gate491inter0), .b(s_332), .O(gate491inter1));
  and2  gate2873(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2874(.a(s_332), .O(gate491inter3));
  inv1  gate2875(.a(s_333), .O(gate491inter4));
  nand2 gate2876(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2877(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2878(.a(G1244), .O(gate491inter7));
  inv1  gate2879(.a(G1245), .O(gate491inter8));
  nand2 gate2880(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2881(.a(s_333), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2882(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2883(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2884(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2899(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2900(.a(gate496inter0), .b(s_336), .O(gate496inter1));
  and2  gate2901(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2902(.a(s_336), .O(gate496inter3));
  inv1  gate2903(.a(s_337), .O(gate496inter4));
  nand2 gate2904(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2905(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2906(.a(G1254), .O(gate496inter7));
  inv1  gate2907(.a(G1255), .O(gate496inter8));
  nand2 gate2908(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2909(.a(s_337), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2910(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2911(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2912(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2521(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2522(.a(gate499inter0), .b(s_282), .O(gate499inter1));
  and2  gate2523(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2524(.a(s_282), .O(gate499inter3));
  inv1  gate2525(.a(s_283), .O(gate499inter4));
  nand2 gate2526(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2527(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2528(.a(G1260), .O(gate499inter7));
  inv1  gate2529(.a(G1261), .O(gate499inter8));
  nand2 gate2530(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2531(.a(s_283), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2532(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2533(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2534(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2829(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2830(.a(gate502inter0), .b(s_326), .O(gate502inter1));
  and2  gate2831(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2832(.a(s_326), .O(gate502inter3));
  inv1  gate2833(.a(s_327), .O(gate502inter4));
  nand2 gate2834(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2835(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2836(.a(G1266), .O(gate502inter7));
  inv1  gate2837(.a(G1267), .O(gate502inter8));
  nand2 gate2838(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2839(.a(s_327), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2840(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2841(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2842(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate827(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate828(.a(gate503inter0), .b(s_40), .O(gate503inter1));
  and2  gate829(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate830(.a(s_40), .O(gate503inter3));
  inv1  gate831(.a(s_41), .O(gate503inter4));
  nand2 gate832(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate833(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate834(.a(G1268), .O(gate503inter7));
  inv1  gate835(.a(G1269), .O(gate503inter8));
  nand2 gate836(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate837(.a(s_41), .b(gate503inter3), .O(gate503inter10));
  nor2  gate838(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate839(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate840(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate617(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate618(.a(gate506inter0), .b(s_10), .O(gate506inter1));
  and2  gate619(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate620(.a(s_10), .O(gate506inter3));
  inv1  gate621(.a(s_11), .O(gate506inter4));
  nand2 gate622(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate623(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate624(.a(G1274), .O(gate506inter7));
  inv1  gate625(.a(G1275), .O(gate506inter8));
  nand2 gate626(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate627(.a(s_11), .b(gate506inter3), .O(gate506inter10));
  nor2  gate628(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate629(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate630(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1093(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1094(.a(gate514inter0), .b(s_78), .O(gate514inter1));
  and2  gate1095(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1096(.a(s_78), .O(gate514inter3));
  inv1  gate1097(.a(s_79), .O(gate514inter4));
  nand2 gate1098(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1099(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1100(.a(G1290), .O(gate514inter7));
  inv1  gate1101(.a(G1291), .O(gate514inter8));
  nand2 gate1102(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1103(.a(s_79), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1104(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1105(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1106(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule