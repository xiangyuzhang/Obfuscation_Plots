module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12;

  xor2  gate483(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate484(.a(gate1inter0), .b(s_40), .O(gate1inter1));
  and2  gate485(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate486(.a(s_40), .O(gate1inter3));
  inv1  gate487(.a(s_41), .O(gate1inter4));
  nand2 gate488(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate489(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate490(.a(N1), .O(gate1inter7));
  inv1  gate491(.a(N5), .O(gate1inter8));
  nand2 gate492(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate493(.a(s_41), .b(gate1inter3), .O(gate1inter10));
  nor2  gate494(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate495(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate496(.a(gate1inter12), .b(gate1inter1), .O(N250));
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate525(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate526(.a(gate6inter0), .b(s_46), .O(gate6inter1));
  and2  gate527(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate528(.a(s_46), .O(gate6inter3));
  inv1  gate529(.a(s_47), .O(gate6inter4));
  nand2 gate530(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate531(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate532(.a(N41), .O(gate6inter7));
  inv1  gate533(.a(N45), .O(gate6inter8));
  nand2 gate534(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate535(.a(s_47), .b(gate6inter3), .O(gate6inter10));
  nor2  gate536(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate537(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate538(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate693(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate694(.a(gate8inter0), .b(s_70), .O(gate8inter1));
  and2  gate695(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate696(.a(s_70), .O(gate8inter3));
  inv1  gate697(.a(s_71), .O(gate8inter4));
  nand2 gate698(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate699(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate700(.a(N57), .O(gate8inter7));
  inv1  gate701(.a(N61), .O(gate8inter8));
  nand2 gate702(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate703(.a(s_71), .b(gate8inter3), .O(gate8inter10));
  nor2  gate704(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate705(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate706(.a(gate8inter12), .b(gate8inter1), .O(N257));
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );

  xor2  gate385(.a(N93), .b(N89), .O(gate12inter0));
  nand2 gate386(.a(gate12inter0), .b(s_26), .O(gate12inter1));
  and2  gate387(.a(N93), .b(N89), .O(gate12inter2));
  inv1  gate388(.a(s_26), .O(gate12inter3));
  inv1  gate389(.a(s_27), .O(gate12inter4));
  nand2 gate390(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate391(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate392(.a(N89), .O(gate12inter7));
  inv1  gate393(.a(N93), .O(gate12inter8));
  nand2 gate394(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate395(.a(s_27), .b(gate12inter3), .O(gate12inter10));
  nor2  gate396(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate397(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate398(.a(gate12inter12), .b(gate12inter1), .O(N261));
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );

  xor2  gate665(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate666(.a(gate15inter0), .b(s_66), .O(gate15inter1));
  and2  gate667(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate668(.a(s_66), .O(gate15inter3));
  inv1  gate669(.a(s_67), .O(gate15inter4));
  nand2 gate670(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate671(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate672(.a(N113), .O(gate15inter7));
  inv1  gate673(.a(N117), .O(gate15inter8));
  nand2 gate674(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate675(.a(s_67), .b(gate15inter3), .O(gate15inter10));
  nor2  gate676(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate677(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate678(.a(gate15inter12), .b(gate15inter1), .O(N264));
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate287(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate288(.a(gate25inter0), .b(s_12), .O(gate25inter1));
  and2  gate289(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate290(.a(s_12), .O(gate25inter3));
  inv1  gate291(.a(s_13), .O(gate25inter4));
  nand2 gate292(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate293(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate294(.a(N1), .O(gate25inter7));
  inv1  gate295(.a(N17), .O(gate25inter8));
  nand2 gate296(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate297(.a(s_13), .b(gate25inter3), .O(gate25inter10));
  nor2  gate298(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate299(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate300(.a(gate25inter12), .b(gate25inter1), .O(N274));

  xor2  gate273(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate274(.a(gate26inter0), .b(s_10), .O(gate26inter1));
  and2  gate275(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate276(.a(s_10), .O(gate26inter3));
  inv1  gate277(.a(s_11), .O(gate26inter4));
  nand2 gate278(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate279(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate280(.a(N33), .O(gate26inter7));
  inv1  gate281(.a(N49), .O(gate26inter8));
  nand2 gate282(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate283(.a(s_11), .b(gate26inter3), .O(gate26inter10));
  nor2  gate284(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate285(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate286(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );

  xor2  gate553(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate554(.a(gate31inter0), .b(s_50), .O(gate31inter1));
  and2  gate555(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate556(.a(s_50), .O(gate31inter3));
  inv1  gate557(.a(s_51), .O(gate31inter4));
  nand2 gate558(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate559(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate560(.a(N13), .O(gate31inter7));
  inv1  gate561(.a(N29), .O(gate31inter8));
  nand2 gate562(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate563(.a(s_51), .b(gate31inter3), .O(gate31inter10));
  nor2  gate564(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate565(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate566(.a(gate31inter12), .b(gate31inter1), .O(N280));
xor2 gate32( .a(N45), .b(N61), .O(N281) );

  xor2  gate245(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate246(.a(gate33inter0), .b(s_6), .O(gate33inter1));
  and2  gate247(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate248(.a(s_6), .O(gate33inter3));
  inv1  gate249(.a(s_7), .O(gate33inter4));
  nand2 gate250(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate251(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate252(.a(N65), .O(gate33inter7));
  inv1  gate253(.a(N81), .O(gate33inter8));
  nand2 gate254(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate255(.a(s_7), .b(gate33inter3), .O(gate33inter10));
  nor2  gate256(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate257(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate258(.a(gate33inter12), .b(gate33inter1), .O(N282));

  xor2  gate637(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate638(.a(gate34inter0), .b(s_62), .O(gate34inter1));
  and2  gate639(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate640(.a(s_62), .O(gate34inter3));
  inv1  gate641(.a(s_63), .O(gate34inter4));
  nand2 gate642(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate643(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate644(.a(N97), .O(gate34inter7));
  inv1  gate645(.a(N113), .O(gate34inter8));
  nand2 gate646(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate647(.a(s_63), .b(gate34inter3), .O(gate34inter10));
  nor2  gate648(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate649(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate650(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );

  xor2  gate301(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate302(.a(gate36inter0), .b(s_14), .O(gate36inter1));
  and2  gate303(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate304(.a(s_14), .O(gate36inter3));
  inv1  gate305(.a(s_15), .O(gate36inter4));
  nand2 gate306(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate307(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate308(.a(N101), .O(gate36inter7));
  inv1  gate309(.a(N117), .O(gate36inter8));
  nand2 gate310(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate311(.a(s_15), .b(gate36inter3), .O(gate36inter10));
  nor2  gate312(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate313(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate314(.a(gate36inter12), .b(gate36inter1), .O(N285));
xor2 gate37( .a(N73), .b(N89), .O(N286) );

  xor2  gate581(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate582(.a(gate38inter0), .b(s_54), .O(gate38inter1));
  and2  gate583(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate584(.a(s_54), .O(gate38inter3));
  inv1  gate585(.a(s_55), .O(gate38inter4));
  nand2 gate586(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate587(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate588(.a(N105), .O(gate38inter7));
  inv1  gate589(.a(N121), .O(gate38inter8));
  nand2 gate590(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate591(.a(s_55), .b(gate38inter3), .O(gate38inter10));
  nor2  gate592(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate593(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate594(.a(gate38inter12), .b(gate38inter1), .O(N287));

  xor2  gate567(.a(N93), .b(N77), .O(gate39inter0));
  nand2 gate568(.a(gate39inter0), .b(s_52), .O(gate39inter1));
  and2  gate569(.a(N93), .b(N77), .O(gate39inter2));
  inv1  gate570(.a(s_52), .O(gate39inter3));
  inv1  gate571(.a(s_53), .O(gate39inter4));
  nand2 gate572(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate573(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate574(.a(N77), .O(gate39inter7));
  inv1  gate575(.a(N93), .O(gate39inter8));
  nand2 gate576(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate577(.a(s_53), .b(gate39inter3), .O(gate39inter10));
  nor2  gate578(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate579(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate580(.a(gate39inter12), .b(gate39inter1), .O(N288));
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );

  xor2  gate623(.a(N257), .b(N256), .O(gate44inter0));
  nand2 gate624(.a(gate44inter0), .b(s_60), .O(gate44inter1));
  and2  gate625(.a(N257), .b(N256), .O(gate44inter2));
  inv1  gate626(.a(s_60), .O(gate44inter3));
  inv1  gate627(.a(s_61), .O(gate44inter4));
  nand2 gate628(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate629(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate630(.a(N256), .O(gate44inter7));
  inv1  gate631(.a(N257), .O(gate44inter8));
  nand2 gate632(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate633(.a(s_61), .b(gate44inter3), .O(gate44inter10));
  nor2  gate634(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate635(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate636(.a(gate44inter12), .b(gate44inter1), .O(N299));

  xor2  gate217(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate218(.a(gate45inter0), .b(s_2), .O(gate45inter1));
  and2  gate219(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate220(.a(s_2), .O(gate45inter3));
  inv1  gate221(.a(s_3), .O(gate45inter4));
  nand2 gate222(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate223(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate224(.a(N258), .O(gate45inter7));
  inv1  gate225(.a(N259), .O(gate45inter8));
  nand2 gate226(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate227(.a(s_3), .b(gate45inter3), .O(gate45inter10));
  nor2  gate228(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate229(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate230(.a(gate45inter12), .b(gate45inter1), .O(N302));
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate427(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate428(.a(gate47inter0), .b(s_32), .O(gate47inter1));
  and2  gate429(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate430(.a(s_32), .O(gate47inter3));
  inv1  gate431(.a(s_33), .O(gate47inter4));
  nand2 gate432(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate433(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate434(.a(N262), .O(gate47inter7));
  inv1  gate435(.a(N263), .O(gate47inter8));
  nand2 gate436(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate437(.a(s_33), .b(gate47inter3), .O(gate47inter10));
  nor2  gate438(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate439(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate440(.a(gate47inter12), .b(gate47inter1), .O(N308));
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );

  xor2  gate231(.a(N289), .b(N288), .O(gate56inter0));
  nand2 gate232(.a(gate56inter0), .b(s_4), .O(gate56inter1));
  and2  gate233(.a(N289), .b(N288), .O(gate56inter2));
  inv1  gate234(.a(s_4), .O(gate56inter3));
  inv1  gate235(.a(s_5), .O(gate56inter4));
  nand2 gate236(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate237(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate238(.a(N288), .O(gate56inter7));
  inv1  gate239(.a(N289), .O(gate56inter8));
  nand2 gate240(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate241(.a(s_5), .b(gate56inter3), .O(gate56inter10));
  nor2  gate242(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate243(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate244(.a(gate56inter12), .b(gate56inter1), .O(N321));

  xor2  gate399(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate400(.a(gate57inter0), .b(s_28), .O(gate57inter1));
  and2  gate401(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate402(.a(s_28), .O(gate57inter3));
  inv1  gate403(.a(s_29), .O(gate57inter4));
  nand2 gate404(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate405(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate406(.a(N290), .O(gate57inter7));
  inv1  gate407(.a(N293), .O(gate57inter8));
  nand2 gate408(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate409(.a(s_29), .b(gate57inter3), .O(gate57inter10));
  nor2  gate410(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate411(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate412(.a(gate57inter12), .b(gate57inter1), .O(N338));
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );

  xor2  gate329(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate330(.a(gate60inter0), .b(s_18), .O(gate60inter1));
  and2  gate331(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate332(.a(s_18), .O(gate60inter3));
  inv1  gate333(.a(s_19), .O(gate60inter4));
  nand2 gate334(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate335(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate336(.a(N293), .O(gate60inter7));
  inv1  gate337(.a(N299), .O(gate60inter8));
  nand2 gate338(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate339(.a(s_19), .b(gate60inter3), .O(gate60inter10));
  nor2  gate340(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate341(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate342(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate679(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate680(.a(gate62inter0), .b(s_68), .O(gate62inter1));
  and2  gate681(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate682(.a(s_68), .O(gate62inter3));
  inv1  gate683(.a(s_69), .O(gate62inter4));
  nand2 gate684(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate685(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate686(.a(N308), .O(gate62inter7));
  inv1  gate687(.a(N311), .O(gate62inter8));
  nand2 gate688(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate689(.a(s_69), .b(gate62inter3), .O(gate62inter10));
  nor2  gate690(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate691(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate692(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate203(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate204(.a(gate65inter0), .b(s_0), .O(gate65inter1));
  and2  gate205(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate206(.a(s_0), .O(gate65inter3));
  inv1  gate207(.a(s_1), .O(gate65inter4));
  nand2 gate208(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate209(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate210(.a(N266), .O(gate65inter7));
  inv1  gate211(.a(N342), .O(gate65inter8));
  nand2 gate212(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate213(.a(s_1), .b(gate65inter3), .O(gate65inter10));
  nor2  gate214(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate215(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate216(.a(gate65inter12), .b(gate65inter1), .O(N346));
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );

  xor2  gate413(.a(N338), .b(N270), .O(gate69inter0));
  nand2 gate414(.a(gate69inter0), .b(s_30), .O(gate69inter1));
  and2  gate415(.a(N338), .b(N270), .O(gate69inter2));
  inv1  gate416(.a(s_30), .O(gate69inter3));
  inv1  gate417(.a(s_31), .O(gate69inter4));
  nand2 gate418(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate419(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate420(.a(N270), .O(gate69inter7));
  inv1  gate421(.a(N338), .O(gate69inter8));
  nand2 gate422(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate423(.a(s_31), .b(gate69inter3), .O(gate69inter10));
  nor2  gate424(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate425(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate426(.a(gate69inter12), .b(gate69inter1), .O(N350));
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );

  xor2  gate441(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate442(.a(gate74inter0), .b(s_34), .O(gate74inter1));
  and2  gate443(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate444(.a(s_34), .O(gate74inter3));
  inv1  gate445(.a(s_35), .O(gate74inter4));
  nand2 gate446(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate447(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate448(.a(N315), .O(gate74inter7));
  inv1  gate449(.a(N347), .O(gate74inter8));
  nand2 gate450(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate451(.a(s_35), .b(gate74inter3), .O(gate74inter10));
  nor2  gate452(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate453(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate454(.a(gate74inter12), .b(gate74inter1), .O(N367));
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );

  xor2  gate609(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate610(.a(gate77inter0), .b(s_58), .O(gate77inter1));
  and2  gate611(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate612(.a(s_58), .O(gate77inter3));
  inv1  gate613(.a(s_59), .O(gate77inter4));
  nand2 gate614(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate615(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate616(.a(N318), .O(gate77inter7));
  inv1  gate617(.a(N350), .O(gate77inter8));
  nand2 gate618(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate619(.a(s_59), .b(gate77inter3), .O(gate77inter10));
  nor2  gate620(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate621(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate622(.a(gate77inter12), .b(gate77inter1), .O(N406));
xor2 gate78( .a(N319), .b(N351), .O(N419) );

  xor2  gate357(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate358(.a(gate79inter0), .b(s_22), .O(gate79inter1));
  and2  gate359(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate360(.a(s_22), .O(gate79inter3));
  inv1  gate361(.a(s_23), .O(gate79inter4));
  nand2 gate362(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate363(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate364(.a(N320), .O(gate79inter7));
  inv1  gate365(.a(N352), .O(gate79inter8));
  nand2 gate366(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate367(.a(s_23), .b(gate79inter3), .O(gate79inter10));
  nor2  gate368(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate369(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate370(.a(gate79inter12), .b(gate79inter1), .O(N432));
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate651(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate652(.a(gate172inter0), .b(s_64), .O(gate172inter1));
  and2  gate653(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate654(.a(s_64), .O(gate172inter3));
  inv1  gate655(.a(s_65), .O(gate172inter4));
  nand2 gate656(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate657(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate658(.a(N5), .O(gate172inter7));
  inv1  gate659(.a(N693), .O(gate172inter8));
  nand2 gate660(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate661(.a(s_65), .b(gate172inter3), .O(gate172inter10));
  nor2  gate662(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate663(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate664(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );

  xor2  gate595(.a(N695), .b(N13), .O(gate174inter0));
  nand2 gate596(.a(gate174inter0), .b(s_56), .O(gate174inter1));
  and2  gate597(.a(N695), .b(N13), .O(gate174inter2));
  inv1  gate598(.a(s_56), .O(gate174inter3));
  inv1  gate599(.a(s_57), .O(gate174inter4));
  nand2 gate600(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate601(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate602(.a(N13), .O(gate174inter7));
  inv1  gate603(.a(N695), .O(gate174inter8));
  nand2 gate604(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate605(.a(s_57), .b(gate174inter3), .O(gate174inter10));
  nor2  gate606(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate607(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate608(.a(gate174inter12), .b(gate174inter1), .O(N727));
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );

  xor2  gate469(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate470(.a(gate179inter0), .b(s_38), .O(gate179inter1));
  and2  gate471(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate472(.a(s_38), .O(gate179inter3));
  inv1  gate473(.a(s_39), .O(gate179inter4));
  nand2 gate474(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate475(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate476(.a(N33), .O(gate179inter7));
  inv1  gate477(.a(N700), .O(gate179inter8));
  nand2 gate478(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate479(.a(s_39), .b(gate179inter3), .O(gate179inter10));
  nor2  gate480(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate481(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate482(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );

  xor2  gate511(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate512(.a(gate183inter0), .b(s_44), .O(gate183inter1));
  and2  gate513(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate514(.a(s_44), .O(gate183inter3));
  inv1  gate515(.a(s_45), .O(gate183inter4));
  nand2 gate516(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate517(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate518(.a(N49), .O(gate183inter7));
  inv1  gate519(.a(N704), .O(gate183inter8));
  nand2 gate520(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate521(.a(s_45), .b(gate183inter3), .O(gate183inter10));
  nor2  gate522(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate523(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate524(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );

  xor2  gate315(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate316(.a(gate185inter0), .b(s_16), .O(gate185inter1));
  and2  gate317(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate318(.a(s_16), .O(gate185inter3));
  inv1  gate319(.a(s_17), .O(gate185inter4));
  nand2 gate320(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate321(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate322(.a(N57), .O(gate185inter7));
  inv1  gate323(.a(N706), .O(gate185inter8));
  nand2 gate324(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate325(.a(s_17), .b(gate185inter3), .O(gate185inter10));
  nor2  gate326(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate327(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate328(.a(gate185inter12), .b(gate185inter1), .O(N738));

  xor2  gate371(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate372(.a(gate186inter0), .b(s_24), .O(gate186inter1));
  and2  gate373(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate374(.a(s_24), .O(gate186inter3));
  inv1  gate375(.a(s_25), .O(gate186inter4));
  nand2 gate376(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate377(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate378(.a(N61), .O(gate186inter7));
  inv1  gate379(.a(N707), .O(gate186inter8));
  nand2 gate380(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate381(.a(s_25), .b(gate186inter3), .O(gate186inter10));
  nor2  gate382(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate383(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate384(.a(gate186inter12), .b(gate186inter1), .O(N739));

  xor2  gate455(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate456(.a(gate187inter0), .b(s_36), .O(gate187inter1));
  and2  gate457(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate458(.a(s_36), .O(gate187inter3));
  inv1  gate459(.a(s_37), .O(gate187inter4));
  nand2 gate460(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate461(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate462(.a(N65), .O(gate187inter7));
  inv1  gate463(.a(N708), .O(gate187inter8));
  nand2 gate464(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate465(.a(s_37), .b(gate187inter3), .O(gate187inter10));
  nor2  gate466(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate467(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate468(.a(gate187inter12), .b(gate187inter1), .O(N740));

  xor2  gate343(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate344(.a(gate188inter0), .b(s_20), .O(gate188inter1));
  and2  gate345(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate346(.a(s_20), .O(gate188inter3));
  inv1  gate347(.a(s_21), .O(gate188inter4));
  nand2 gate348(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate349(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate350(.a(N69), .O(gate188inter7));
  inv1  gate351(.a(N709), .O(gate188inter8));
  nand2 gate352(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate353(.a(s_21), .b(gate188inter3), .O(gate188inter10));
  nor2  gate354(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate355(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate356(.a(gate188inter12), .b(gate188inter1), .O(N741));
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );

  xor2  gate497(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate498(.a(gate194inter0), .b(s_42), .O(gate194inter1));
  and2  gate499(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate500(.a(s_42), .O(gate194inter3));
  inv1  gate501(.a(s_43), .O(gate194inter4));
  nand2 gate502(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate503(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate504(.a(N93), .O(gate194inter7));
  inv1  gate505(.a(N715), .O(gate194inter8));
  nand2 gate506(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate507(.a(s_43), .b(gate194inter3), .O(gate194inter10));
  nor2  gate508(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate509(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate510(.a(gate194inter12), .b(gate194inter1), .O(N747));
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );

  xor2  gate539(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate540(.a(gate197inter0), .b(s_48), .O(gate197inter1));
  and2  gate541(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate542(.a(s_48), .O(gate197inter3));
  inv1  gate543(.a(s_49), .O(gate197inter4));
  nand2 gate544(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate545(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate546(.a(N105), .O(gate197inter7));
  inv1  gate547(.a(N718), .O(gate197inter8));
  nand2 gate548(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate549(.a(s_49), .b(gate197inter3), .O(gate197inter10));
  nor2  gate550(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate551(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate552(.a(gate197inter12), .b(gate197inter1), .O(N750));

  xor2  gate259(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate260(.a(gate198inter0), .b(s_8), .O(gate198inter1));
  and2  gate261(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate262(.a(s_8), .O(gate198inter3));
  inv1  gate263(.a(s_9), .O(gate198inter4));
  nand2 gate264(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate265(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate266(.a(N109), .O(gate198inter7));
  inv1  gate267(.a(N719), .O(gate198inter8));
  nand2 gate268(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate269(.a(s_9), .b(gate198inter3), .O(gate198inter10));
  nor2  gate270(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate271(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate272(.a(gate198inter12), .b(gate198inter1), .O(N751));
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule