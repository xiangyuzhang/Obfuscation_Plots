module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1275(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1276(.a(gate9inter0), .b(s_104), .O(gate9inter1));
  and2  gate1277(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1278(.a(s_104), .O(gate9inter3));
  inv1  gate1279(.a(s_105), .O(gate9inter4));
  nand2 gate1280(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1281(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1282(.a(G1), .O(gate9inter7));
  inv1  gate1283(.a(G2), .O(gate9inter8));
  nand2 gate1284(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1285(.a(s_105), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1286(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1287(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1288(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2059(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2060(.a(gate17inter0), .b(s_216), .O(gate17inter1));
  and2  gate2061(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2062(.a(s_216), .O(gate17inter3));
  inv1  gate2063(.a(s_217), .O(gate17inter4));
  nand2 gate2064(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2065(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2066(.a(G17), .O(gate17inter7));
  inv1  gate2067(.a(G18), .O(gate17inter8));
  nand2 gate2068(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2069(.a(s_217), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2070(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2071(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2072(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate701(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate702(.a(gate19inter0), .b(s_22), .O(gate19inter1));
  and2  gate703(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate704(.a(s_22), .O(gate19inter3));
  inv1  gate705(.a(s_23), .O(gate19inter4));
  nand2 gate706(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate707(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate708(.a(G21), .O(gate19inter7));
  inv1  gate709(.a(G22), .O(gate19inter8));
  nand2 gate710(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate711(.a(s_23), .b(gate19inter3), .O(gate19inter10));
  nor2  gate712(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate713(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate714(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1513(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1514(.a(gate21inter0), .b(s_138), .O(gate21inter1));
  and2  gate1515(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1516(.a(s_138), .O(gate21inter3));
  inv1  gate1517(.a(s_139), .O(gate21inter4));
  nand2 gate1518(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1519(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1520(.a(G25), .O(gate21inter7));
  inv1  gate1521(.a(G26), .O(gate21inter8));
  nand2 gate1522(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1523(.a(s_139), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1524(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1525(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1526(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1779(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1780(.a(gate24inter0), .b(s_176), .O(gate24inter1));
  and2  gate1781(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1782(.a(s_176), .O(gate24inter3));
  inv1  gate1783(.a(s_177), .O(gate24inter4));
  nand2 gate1784(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1785(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1786(.a(G31), .O(gate24inter7));
  inv1  gate1787(.a(G32), .O(gate24inter8));
  nand2 gate1788(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1789(.a(s_177), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1790(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1791(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1792(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1751(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1752(.a(gate25inter0), .b(s_172), .O(gate25inter1));
  and2  gate1753(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1754(.a(s_172), .O(gate25inter3));
  inv1  gate1755(.a(s_173), .O(gate25inter4));
  nand2 gate1756(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1757(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1758(.a(G1), .O(gate25inter7));
  inv1  gate1759(.a(G5), .O(gate25inter8));
  nand2 gate1760(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1761(.a(s_173), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1762(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1763(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1764(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1793(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1794(.a(gate27inter0), .b(s_178), .O(gate27inter1));
  and2  gate1795(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1796(.a(s_178), .O(gate27inter3));
  inv1  gate1797(.a(s_179), .O(gate27inter4));
  nand2 gate1798(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1799(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1800(.a(G2), .O(gate27inter7));
  inv1  gate1801(.a(G6), .O(gate27inter8));
  nand2 gate1802(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1803(.a(s_179), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1804(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1805(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1806(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2129(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2130(.a(gate33inter0), .b(s_226), .O(gate33inter1));
  and2  gate2131(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2132(.a(s_226), .O(gate33inter3));
  inv1  gate2133(.a(s_227), .O(gate33inter4));
  nand2 gate2134(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2135(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2136(.a(G17), .O(gate33inter7));
  inv1  gate2137(.a(G21), .O(gate33inter8));
  nand2 gate2138(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2139(.a(s_227), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2140(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2141(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2142(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate2073(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2074(.a(gate35inter0), .b(s_218), .O(gate35inter1));
  and2  gate2075(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2076(.a(s_218), .O(gate35inter3));
  inv1  gate2077(.a(s_219), .O(gate35inter4));
  nand2 gate2078(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2079(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2080(.a(G18), .O(gate35inter7));
  inv1  gate2081(.a(G22), .O(gate35inter8));
  nand2 gate2082(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2083(.a(s_219), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2084(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2085(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2086(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1429(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1430(.a(gate36inter0), .b(s_126), .O(gate36inter1));
  and2  gate1431(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1432(.a(s_126), .O(gate36inter3));
  inv1  gate1433(.a(s_127), .O(gate36inter4));
  nand2 gate1434(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1435(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1436(.a(G26), .O(gate36inter7));
  inv1  gate1437(.a(G30), .O(gate36inter8));
  nand2 gate1438(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1439(.a(s_127), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1440(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1441(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1442(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1023(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1024(.a(gate38inter0), .b(s_68), .O(gate38inter1));
  and2  gate1025(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1026(.a(s_68), .O(gate38inter3));
  inv1  gate1027(.a(s_69), .O(gate38inter4));
  nand2 gate1028(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1029(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1030(.a(G27), .O(gate38inter7));
  inv1  gate1031(.a(G31), .O(gate38inter8));
  nand2 gate1032(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1033(.a(s_69), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1034(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1035(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1036(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1233(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1234(.a(gate39inter0), .b(s_98), .O(gate39inter1));
  and2  gate1235(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1236(.a(s_98), .O(gate39inter3));
  inv1  gate1237(.a(s_99), .O(gate39inter4));
  nand2 gate1238(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1239(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1240(.a(G20), .O(gate39inter7));
  inv1  gate1241(.a(G24), .O(gate39inter8));
  nand2 gate1242(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1243(.a(s_99), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1244(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1245(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1246(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2241(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2242(.a(gate42inter0), .b(s_242), .O(gate42inter1));
  and2  gate2243(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2244(.a(s_242), .O(gate42inter3));
  inv1  gate2245(.a(s_243), .O(gate42inter4));
  nand2 gate2246(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2247(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2248(.a(G2), .O(gate42inter7));
  inv1  gate2249(.a(G266), .O(gate42inter8));
  nand2 gate2250(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2251(.a(s_243), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2252(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2253(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2254(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1527(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1528(.a(gate44inter0), .b(s_140), .O(gate44inter1));
  and2  gate1529(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1530(.a(s_140), .O(gate44inter3));
  inv1  gate1531(.a(s_141), .O(gate44inter4));
  nand2 gate1532(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1533(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1534(.a(G4), .O(gate44inter7));
  inv1  gate1535(.a(G269), .O(gate44inter8));
  nand2 gate1536(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1537(.a(s_141), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1538(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1539(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1540(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2031(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2032(.a(gate45inter0), .b(s_212), .O(gate45inter1));
  and2  gate2033(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2034(.a(s_212), .O(gate45inter3));
  inv1  gate2035(.a(s_213), .O(gate45inter4));
  nand2 gate2036(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2037(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2038(.a(G5), .O(gate45inter7));
  inv1  gate2039(.a(G272), .O(gate45inter8));
  nand2 gate2040(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2041(.a(s_213), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2042(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2043(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2044(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2185(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2186(.a(gate48inter0), .b(s_234), .O(gate48inter1));
  and2  gate2187(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2188(.a(s_234), .O(gate48inter3));
  inv1  gate2189(.a(s_235), .O(gate48inter4));
  nand2 gate2190(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2191(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2192(.a(G8), .O(gate48inter7));
  inv1  gate2193(.a(G275), .O(gate48inter8));
  nand2 gate2194(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2195(.a(s_235), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2196(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2197(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2198(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate981(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate982(.a(gate53inter0), .b(s_62), .O(gate53inter1));
  and2  gate983(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate984(.a(s_62), .O(gate53inter3));
  inv1  gate985(.a(s_63), .O(gate53inter4));
  nand2 gate986(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate987(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate988(.a(G13), .O(gate53inter7));
  inv1  gate989(.a(G284), .O(gate53inter8));
  nand2 gate990(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate991(.a(s_63), .b(gate53inter3), .O(gate53inter10));
  nor2  gate992(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate993(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate994(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate603(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate604(.a(gate62inter0), .b(s_8), .O(gate62inter1));
  and2  gate605(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate606(.a(s_8), .O(gate62inter3));
  inv1  gate607(.a(s_9), .O(gate62inter4));
  nand2 gate608(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate609(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate610(.a(G22), .O(gate62inter7));
  inv1  gate611(.a(G296), .O(gate62inter8));
  nand2 gate612(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate613(.a(s_9), .b(gate62inter3), .O(gate62inter10));
  nor2  gate614(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate615(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate616(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2325(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2326(.a(gate66inter0), .b(s_254), .O(gate66inter1));
  and2  gate2327(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2328(.a(s_254), .O(gate66inter3));
  inv1  gate2329(.a(s_255), .O(gate66inter4));
  nand2 gate2330(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2331(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2332(.a(G26), .O(gate66inter7));
  inv1  gate2333(.a(G302), .O(gate66inter8));
  nand2 gate2334(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2335(.a(s_255), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2336(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2337(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2338(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate687(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate688(.a(gate67inter0), .b(s_20), .O(gate67inter1));
  and2  gate689(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate690(.a(s_20), .O(gate67inter3));
  inv1  gate691(.a(s_21), .O(gate67inter4));
  nand2 gate692(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate693(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate694(.a(G27), .O(gate67inter7));
  inv1  gate695(.a(G305), .O(gate67inter8));
  nand2 gate696(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate697(.a(s_21), .b(gate67inter3), .O(gate67inter10));
  nor2  gate698(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate699(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate700(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate715(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate716(.a(gate71inter0), .b(s_24), .O(gate71inter1));
  and2  gate717(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate718(.a(s_24), .O(gate71inter3));
  inv1  gate719(.a(s_25), .O(gate71inter4));
  nand2 gate720(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate721(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate722(.a(G31), .O(gate71inter7));
  inv1  gate723(.a(G311), .O(gate71inter8));
  nand2 gate724(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate725(.a(s_25), .b(gate71inter3), .O(gate71inter10));
  nor2  gate726(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate727(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate728(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2283(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2284(.a(gate72inter0), .b(s_248), .O(gate72inter1));
  and2  gate2285(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2286(.a(s_248), .O(gate72inter3));
  inv1  gate2287(.a(s_249), .O(gate72inter4));
  nand2 gate2288(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2289(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2290(.a(G32), .O(gate72inter7));
  inv1  gate2291(.a(G311), .O(gate72inter8));
  nand2 gate2292(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2293(.a(s_249), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2294(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2295(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2296(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate771(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate772(.a(gate73inter0), .b(s_32), .O(gate73inter1));
  and2  gate773(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate774(.a(s_32), .O(gate73inter3));
  inv1  gate775(.a(s_33), .O(gate73inter4));
  nand2 gate776(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate777(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate778(.a(G1), .O(gate73inter7));
  inv1  gate779(.a(G314), .O(gate73inter8));
  nand2 gate780(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate781(.a(s_33), .b(gate73inter3), .O(gate73inter10));
  nor2  gate782(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate783(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate784(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate561(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate562(.a(gate74inter0), .b(s_2), .O(gate74inter1));
  and2  gate563(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate564(.a(s_2), .O(gate74inter3));
  inv1  gate565(.a(s_3), .O(gate74inter4));
  nand2 gate566(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate567(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate568(.a(G5), .O(gate74inter7));
  inv1  gate569(.a(G314), .O(gate74inter8));
  nand2 gate570(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate571(.a(s_3), .b(gate74inter3), .O(gate74inter10));
  nor2  gate572(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate573(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate574(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1765(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1766(.a(gate75inter0), .b(s_174), .O(gate75inter1));
  and2  gate1767(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1768(.a(s_174), .O(gate75inter3));
  inv1  gate1769(.a(s_175), .O(gate75inter4));
  nand2 gate1770(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1771(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1772(.a(G9), .O(gate75inter7));
  inv1  gate1773(.a(G317), .O(gate75inter8));
  nand2 gate1774(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1775(.a(s_175), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1776(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1777(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1778(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate645(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate646(.a(gate78inter0), .b(s_14), .O(gate78inter1));
  and2  gate647(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate648(.a(s_14), .O(gate78inter3));
  inv1  gate649(.a(s_15), .O(gate78inter4));
  nand2 gate650(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate651(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate652(.a(G6), .O(gate78inter7));
  inv1  gate653(.a(G320), .O(gate78inter8));
  nand2 gate654(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate655(.a(s_15), .b(gate78inter3), .O(gate78inter10));
  nor2  gate656(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate657(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate658(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1373(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1374(.a(gate79inter0), .b(s_118), .O(gate79inter1));
  and2  gate1375(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1376(.a(s_118), .O(gate79inter3));
  inv1  gate1377(.a(s_119), .O(gate79inter4));
  nand2 gate1378(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1379(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1380(.a(G10), .O(gate79inter7));
  inv1  gate1381(.a(G323), .O(gate79inter8));
  nand2 gate1382(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1383(.a(s_119), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1384(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1385(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1386(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1625(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1626(.a(gate94inter0), .b(s_154), .O(gate94inter1));
  and2  gate1627(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1628(.a(s_154), .O(gate94inter3));
  inv1  gate1629(.a(s_155), .O(gate94inter4));
  nand2 gate1630(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1631(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1632(.a(G22), .O(gate94inter7));
  inv1  gate1633(.a(G344), .O(gate94inter8));
  nand2 gate1634(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1635(.a(s_155), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1636(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1637(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1638(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1443(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1444(.a(gate98inter0), .b(s_128), .O(gate98inter1));
  and2  gate1445(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1446(.a(s_128), .O(gate98inter3));
  inv1  gate1447(.a(s_129), .O(gate98inter4));
  nand2 gate1448(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1449(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1450(.a(G23), .O(gate98inter7));
  inv1  gate1451(.a(G350), .O(gate98inter8));
  nand2 gate1452(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1453(.a(s_129), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1454(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1455(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1456(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1975(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1976(.a(gate104inter0), .b(s_204), .O(gate104inter1));
  and2  gate1977(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1978(.a(s_204), .O(gate104inter3));
  inv1  gate1979(.a(s_205), .O(gate104inter4));
  nand2 gate1980(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1981(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1982(.a(G32), .O(gate104inter7));
  inv1  gate1983(.a(G359), .O(gate104inter8));
  nand2 gate1984(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1985(.a(s_205), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1986(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1987(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1988(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2297(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2298(.a(gate106inter0), .b(s_250), .O(gate106inter1));
  and2  gate2299(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2300(.a(s_250), .O(gate106inter3));
  inv1  gate2301(.a(s_251), .O(gate106inter4));
  nand2 gate2302(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2303(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2304(.a(G364), .O(gate106inter7));
  inv1  gate2305(.a(G365), .O(gate106inter8));
  nand2 gate2306(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2307(.a(s_251), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2308(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2309(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2310(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1737(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1738(.a(gate108inter0), .b(s_170), .O(gate108inter1));
  and2  gate1739(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1740(.a(s_170), .O(gate108inter3));
  inv1  gate1741(.a(s_171), .O(gate108inter4));
  nand2 gate1742(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1743(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1744(.a(G368), .O(gate108inter7));
  inv1  gate1745(.a(G369), .O(gate108inter8));
  nand2 gate1746(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1747(.a(s_171), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1748(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1749(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1750(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1555(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1556(.a(gate119inter0), .b(s_144), .O(gate119inter1));
  and2  gate1557(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1558(.a(s_144), .O(gate119inter3));
  inv1  gate1559(.a(s_145), .O(gate119inter4));
  nand2 gate1560(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1561(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1562(.a(G390), .O(gate119inter7));
  inv1  gate1563(.a(G391), .O(gate119inter8));
  nand2 gate1564(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1565(.a(s_145), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1566(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1567(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1568(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate813(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate814(.a(gate120inter0), .b(s_38), .O(gate120inter1));
  and2  gate815(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate816(.a(s_38), .O(gate120inter3));
  inv1  gate817(.a(s_39), .O(gate120inter4));
  nand2 gate818(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate819(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate820(.a(G392), .O(gate120inter7));
  inv1  gate821(.a(G393), .O(gate120inter8));
  nand2 gate822(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate823(.a(s_39), .b(gate120inter3), .O(gate120inter10));
  nor2  gate824(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate825(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate826(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1051(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1052(.a(gate121inter0), .b(s_72), .O(gate121inter1));
  and2  gate1053(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1054(.a(s_72), .O(gate121inter3));
  inv1  gate1055(.a(s_73), .O(gate121inter4));
  nand2 gate1056(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1057(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1058(.a(G394), .O(gate121inter7));
  inv1  gate1059(.a(G395), .O(gate121inter8));
  nand2 gate1060(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1061(.a(s_73), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1062(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1063(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1064(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1933(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1934(.a(gate126inter0), .b(s_198), .O(gate126inter1));
  and2  gate1935(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1936(.a(s_198), .O(gate126inter3));
  inv1  gate1937(.a(s_199), .O(gate126inter4));
  nand2 gate1938(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1939(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1940(.a(G404), .O(gate126inter7));
  inv1  gate1941(.a(G405), .O(gate126inter8));
  nand2 gate1942(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1943(.a(s_199), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1944(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1945(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1946(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate995(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate996(.a(gate127inter0), .b(s_64), .O(gate127inter1));
  and2  gate997(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate998(.a(s_64), .O(gate127inter3));
  inv1  gate999(.a(s_65), .O(gate127inter4));
  nand2 gate1000(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1001(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1002(.a(G406), .O(gate127inter7));
  inv1  gate1003(.a(G407), .O(gate127inter8));
  nand2 gate1004(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1005(.a(s_65), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1006(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1007(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1008(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1317(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1318(.a(gate132inter0), .b(s_110), .O(gate132inter1));
  and2  gate1319(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1320(.a(s_110), .O(gate132inter3));
  inv1  gate1321(.a(s_111), .O(gate132inter4));
  nand2 gate1322(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1323(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1324(.a(G416), .O(gate132inter7));
  inv1  gate1325(.a(G417), .O(gate132inter8));
  nand2 gate1326(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1327(.a(s_111), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1328(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1329(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1330(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1107(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1108(.a(gate135inter0), .b(s_80), .O(gate135inter1));
  and2  gate1109(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1110(.a(s_80), .O(gate135inter3));
  inv1  gate1111(.a(s_81), .O(gate135inter4));
  nand2 gate1112(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1113(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1114(.a(G422), .O(gate135inter7));
  inv1  gate1115(.a(G423), .O(gate135inter8));
  nand2 gate1116(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1117(.a(s_81), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1118(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1119(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1120(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2339(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2340(.a(gate142inter0), .b(s_256), .O(gate142inter1));
  and2  gate2341(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2342(.a(s_256), .O(gate142inter3));
  inv1  gate2343(.a(s_257), .O(gate142inter4));
  nand2 gate2344(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2345(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2346(.a(G456), .O(gate142inter7));
  inv1  gate2347(.a(G459), .O(gate142inter8));
  nand2 gate2348(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2349(.a(s_257), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2350(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2351(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2352(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate2227(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2228(.a(gate143inter0), .b(s_240), .O(gate143inter1));
  and2  gate2229(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2230(.a(s_240), .O(gate143inter3));
  inv1  gate2231(.a(s_241), .O(gate143inter4));
  nand2 gate2232(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2233(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2234(.a(G462), .O(gate143inter7));
  inv1  gate2235(.a(G465), .O(gate143inter8));
  nand2 gate2236(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2237(.a(s_241), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2238(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2239(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2240(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1919(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1920(.a(gate146inter0), .b(s_196), .O(gate146inter1));
  and2  gate1921(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1922(.a(s_196), .O(gate146inter3));
  inv1  gate1923(.a(s_197), .O(gate146inter4));
  nand2 gate1924(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1925(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1926(.a(G480), .O(gate146inter7));
  inv1  gate1927(.a(G483), .O(gate146inter8));
  nand2 gate1928(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1929(.a(s_197), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1930(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1931(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1932(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1989(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1990(.a(gate147inter0), .b(s_206), .O(gate147inter1));
  and2  gate1991(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1992(.a(s_206), .O(gate147inter3));
  inv1  gate1993(.a(s_207), .O(gate147inter4));
  nand2 gate1994(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1995(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1996(.a(G486), .O(gate147inter7));
  inv1  gate1997(.a(G489), .O(gate147inter8));
  nand2 gate1998(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1999(.a(s_207), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2000(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2001(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2002(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate883(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate884(.a(gate150inter0), .b(s_48), .O(gate150inter1));
  and2  gate885(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate886(.a(s_48), .O(gate150inter3));
  inv1  gate887(.a(s_49), .O(gate150inter4));
  nand2 gate888(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate889(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate890(.a(G504), .O(gate150inter7));
  inv1  gate891(.a(G507), .O(gate150inter8));
  nand2 gate892(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate893(.a(s_49), .b(gate150inter3), .O(gate150inter10));
  nor2  gate894(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate895(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate896(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1359(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1360(.a(gate155inter0), .b(s_116), .O(gate155inter1));
  and2  gate1361(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1362(.a(s_116), .O(gate155inter3));
  inv1  gate1363(.a(s_117), .O(gate155inter4));
  nand2 gate1364(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1365(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1366(.a(G432), .O(gate155inter7));
  inv1  gate1367(.a(G525), .O(gate155inter8));
  nand2 gate1368(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1369(.a(s_117), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1370(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1371(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1372(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate659(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate660(.a(gate160inter0), .b(s_16), .O(gate160inter1));
  and2  gate661(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate662(.a(s_16), .O(gate160inter3));
  inv1  gate663(.a(s_17), .O(gate160inter4));
  nand2 gate664(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate665(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate666(.a(G447), .O(gate160inter7));
  inv1  gate667(.a(G531), .O(gate160inter8));
  nand2 gate668(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate669(.a(s_17), .b(gate160inter3), .O(gate160inter10));
  nor2  gate670(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate671(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate672(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2255(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2256(.a(gate162inter0), .b(s_244), .O(gate162inter1));
  and2  gate2257(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2258(.a(s_244), .O(gate162inter3));
  inv1  gate2259(.a(s_245), .O(gate162inter4));
  nand2 gate2260(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2261(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2262(.a(G453), .O(gate162inter7));
  inv1  gate2263(.a(G534), .O(gate162inter8));
  nand2 gate2264(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2265(.a(s_245), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2266(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2267(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2268(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1415(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1416(.a(gate168inter0), .b(s_124), .O(gate168inter1));
  and2  gate1417(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1418(.a(s_124), .O(gate168inter3));
  inv1  gate1419(.a(s_125), .O(gate168inter4));
  nand2 gate1420(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1421(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1422(.a(G471), .O(gate168inter7));
  inv1  gate1423(.a(G543), .O(gate168inter8));
  nand2 gate1424(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1425(.a(s_125), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1426(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1427(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1428(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate2213(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2214(.a(gate177inter0), .b(s_238), .O(gate177inter1));
  and2  gate2215(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2216(.a(s_238), .O(gate177inter3));
  inv1  gate2217(.a(s_239), .O(gate177inter4));
  nand2 gate2218(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2219(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2220(.a(G498), .O(gate177inter7));
  inv1  gate2221(.a(G558), .O(gate177inter8));
  nand2 gate2222(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2223(.a(s_239), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2224(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2225(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2226(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2367(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2368(.a(gate181inter0), .b(s_260), .O(gate181inter1));
  and2  gate2369(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2370(.a(s_260), .O(gate181inter3));
  inv1  gate2371(.a(s_261), .O(gate181inter4));
  nand2 gate2372(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2373(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2374(.a(G510), .O(gate181inter7));
  inv1  gate2375(.a(G564), .O(gate181inter8));
  nand2 gate2376(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2377(.a(s_261), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2378(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2379(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2380(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1807(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1808(.a(gate184inter0), .b(s_180), .O(gate184inter1));
  and2  gate1809(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1810(.a(s_180), .O(gate184inter3));
  inv1  gate1811(.a(s_181), .O(gate184inter4));
  nand2 gate1812(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1813(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1814(.a(G519), .O(gate184inter7));
  inv1  gate1815(.a(G567), .O(gate184inter8));
  nand2 gate1816(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1817(.a(s_181), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1818(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1819(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1820(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1471(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1472(.a(gate187inter0), .b(s_132), .O(gate187inter1));
  and2  gate1473(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1474(.a(s_132), .O(gate187inter3));
  inv1  gate1475(.a(s_133), .O(gate187inter4));
  nand2 gate1476(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1477(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1478(.a(G574), .O(gate187inter7));
  inv1  gate1479(.a(G575), .O(gate187inter8));
  nand2 gate1480(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1481(.a(s_133), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1482(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1483(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1484(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2087(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2088(.a(gate193inter0), .b(s_220), .O(gate193inter1));
  and2  gate2089(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2090(.a(s_220), .O(gate193inter3));
  inv1  gate2091(.a(s_221), .O(gate193inter4));
  nand2 gate2092(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2093(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2094(.a(G586), .O(gate193inter7));
  inv1  gate2095(.a(G587), .O(gate193inter8));
  nand2 gate2096(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2097(.a(s_221), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2098(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2099(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2100(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate2199(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2200(.a(gate194inter0), .b(s_236), .O(gate194inter1));
  and2  gate2201(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2202(.a(s_236), .O(gate194inter3));
  inv1  gate2203(.a(s_237), .O(gate194inter4));
  nand2 gate2204(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2205(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2206(.a(G588), .O(gate194inter7));
  inv1  gate2207(.a(G589), .O(gate194inter8));
  nand2 gate2208(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2209(.a(s_237), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2210(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2211(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2212(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1331(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1332(.a(gate196inter0), .b(s_112), .O(gate196inter1));
  and2  gate1333(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1334(.a(s_112), .O(gate196inter3));
  inv1  gate1335(.a(s_113), .O(gate196inter4));
  nand2 gate1336(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1337(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1338(.a(G592), .O(gate196inter7));
  inv1  gate1339(.a(G593), .O(gate196inter8));
  nand2 gate1340(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1341(.a(s_113), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1342(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1343(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1344(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate953(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate954(.a(gate202inter0), .b(s_58), .O(gate202inter1));
  and2  gate955(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate956(.a(s_58), .O(gate202inter3));
  inv1  gate957(.a(s_59), .O(gate202inter4));
  nand2 gate958(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate959(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate960(.a(G612), .O(gate202inter7));
  inv1  gate961(.a(G617), .O(gate202inter8));
  nand2 gate962(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate963(.a(s_59), .b(gate202inter3), .O(gate202inter10));
  nor2  gate964(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate965(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate966(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate743(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate744(.a(gate203inter0), .b(s_28), .O(gate203inter1));
  and2  gate745(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate746(.a(s_28), .O(gate203inter3));
  inv1  gate747(.a(s_29), .O(gate203inter4));
  nand2 gate748(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate749(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate750(.a(G602), .O(gate203inter7));
  inv1  gate751(.a(G612), .O(gate203inter8));
  nand2 gate752(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate753(.a(s_29), .b(gate203inter3), .O(gate203inter10));
  nor2  gate754(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate755(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate756(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate673(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate674(.a(gate204inter0), .b(s_18), .O(gate204inter1));
  and2  gate675(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate676(.a(s_18), .O(gate204inter3));
  inv1  gate677(.a(s_19), .O(gate204inter4));
  nand2 gate678(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate679(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate680(.a(G607), .O(gate204inter7));
  inv1  gate681(.a(G617), .O(gate204inter8));
  nand2 gate682(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate683(.a(s_19), .b(gate204inter3), .O(gate204inter10));
  nor2  gate684(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate685(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate686(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2157(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2158(.a(gate206inter0), .b(s_230), .O(gate206inter1));
  and2  gate2159(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2160(.a(s_230), .O(gate206inter3));
  inv1  gate2161(.a(s_231), .O(gate206inter4));
  nand2 gate2162(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2163(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2164(.a(G632), .O(gate206inter7));
  inv1  gate2165(.a(G637), .O(gate206inter8));
  nand2 gate2166(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2167(.a(s_231), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2168(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2169(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2170(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2101(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2102(.a(gate209inter0), .b(s_222), .O(gate209inter1));
  and2  gate2103(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2104(.a(s_222), .O(gate209inter3));
  inv1  gate2105(.a(s_223), .O(gate209inter4));
  nand2 gate2106(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2107(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2108(.a(G602), .O(gate209inter7));
  inv1  gate2109(.a(G666), .O(gate209inter8));
  nand2 gate2110(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2111(.a(s_223), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2112(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2113(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2114(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2143(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2144(.a(gate210inter0), .b(s_228), .O(gate210inter1));
  and2  gate2145(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2146(.a(s_228), .O(gate210inter3));
  inv1  gate2147(.a(s_229), .O(gate210inter4));
  nand2 gate2148(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2149(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2150(.a(G607), .O(gate210inter7));
  inv1  gate2151(.a(G666), .O(gate210inter8));
  nand2 gate2152(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2153(.a(s_229), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2154(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2155(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2156(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1611(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1612(.a(gate212inter0), .b(s_152), .O(gate212inter1));
  and2  gate1613(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1614(.a(s_152), .O(gate212inter3));
  inv1  gate1615(.a(s_153), .O(gate212inter4));
  nand2 gate1616(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1617(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1618(.a(G617), .O(gate212inter7));
  inv1  gate1619(.a(G669), .O(gate212inter8));
  nand2 gate1620(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1621(.a(s_153), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1622(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1623(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1624(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate2353(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2354(.a(gate213inter0), .b(s_258), .O(gate213inter1));
  and2  gate2355(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2356(.a(s_258), .O(gate213inter3));
  inv1  gate2357(.a(s_259), .O(gate213inter4));
  nand2 gate2358(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2359(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2360(.a(G602), .O(gate213inter7));
  inv1  gate2361(.a(G672), .O(gate213inter8));
  nand2 gate2362(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2363(.a(s_259), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2364(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2365(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2366(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate967(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate968(.a(gate215inter0), .b(s_60), .O(gate215inter1));
  and2  gate969(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate970(.a(s_60), .O(gate215inter3));
  inv1  gate971(.a(s_61), .O(gate215inter4));
  nand2 gate972(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate973(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate974(.a(G607), .O(gate215inter7));
  inv1  gate975(.a(G675), .O(gate215inter8));
  nand2 gate976(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate977(.a(s_61), .b(gate215inter3), .O(gate215inter10));
  nor2  gate978(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate979(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate980(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1009(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1010(.a(gate218inter0), .b(s_66), .O(gate218inter1));
  and2  gate1011(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1012(.a(s_66), .O(gate218inter3));
  inv1  gate1013(.a(s_67), .O(gate218inter4));
  nand2 gate1014(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1015(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1016(.a(G627), .O(gate218inter7));
  inv1  gate1017(.a(G678), .O(gate218inter8));
  nand2 gate1018(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1019(.a(s_67), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1020(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1021(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1022(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate631(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate632(.a(gate227inter0), .b(s_12), .O(gate227inter1));
  and2  gate633(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate634(.a(s_12), .O(gate227inter3));
  inv1  gate635(.a(s_13), .O(gate227inter4));
  nand2 gate636(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate637(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate638(.a(G694), .O(gate227inter7));
  inv1  gate639(.a(G695), .O(gate227inter8));
  nand2 gate640(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate641(.a(s_13), .b(gate227inter3), .O(gate227inter10));
  nor2  gate642(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate643(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate644(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate841(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate842(.a(gate229inter0), .b(s_42), .O(gate229inter1));
  and2  gate843(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate844(.a(s_42), .O(gate229inter3));
  inv1  gate845(.a(s_43), .O(gate229inter4));
  nand2 gate846(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate847(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate848(.a(G698), .O(gate229inter7));
  inv1  gate849(.a(G699), .O(gate229inter8));
  nand2 gate850(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate851(.a(s_43), .b(gate229inter3), .O(gate229inter10));
  nor2  gate852(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate853(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate854(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1065(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1066(.a(gate231inter0), .b(s_74), .O(gate231inter1));
  and2  gate1067(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1068(.a(s_74), .O(gate231inter3));
  inv1  gate1069(.a(s_75), .O(gate231inter4));
  nand2 gate1070(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1071(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1072(.a(G702), .O(gate231inter7));
  inv1  gate1073(.a(G703), .O(gate231inter8));
  nand2 gate1074(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1075(.a(s_75), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1076(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1077(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1078(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1905(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1906(.a(gate233inter0), .b(s_194), .O(gate233inter1));
  and2  gate1907(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1908(.a(s_194), .O(gate233inter3));
  inv1  gate1909(.a(s_195), .O(gate233inter4));
  nand2 gate1910(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1911(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1912(.a(G242), .O(gate233inter7));
  inv1  gate1913(.a(G718), .O(gate233inter8));
  nand2 gate1914(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1915(.a(s_195), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1916(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1917(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1918(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1863(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1864(.a(gate243inter0), .b(s_188), .O(gate243inter1));
  and2  gate1865(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1866(.a(s_188), .O(gate243inter3));
  inv1  gate1867(.a(s_189), .O(gate243inter4));
  nand2 gate1868(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1869(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1870(.a(G245), .O(gate243inter7));
  inv1  gate1871(.a(G733), .O(gate243inter8));
  nand2 gate1872(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1873(.a(s_189), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1874(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1875(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1876(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate869(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate870(.a(gate248inter0), .b(s_46), .O(gate248inter1));
  and2  gate871(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate872(.a(s_46), .O(gate248inter3));
  inv1  gate873(.a(s_47), .O(gate248inter4));
  nand2 gate874(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate875(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate876(.a(G727), .O(gate248inter7));
  inv1  gate877(.a(G739), .O(gate248inter8));
  nand2 gate878(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate879(.a(s_47), .b(gate248inter3), .O(gate248inter10));
  nor2  gate880(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate881(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate882(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate575(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate576(.a(gate249inter0), .b(s_4), .O(gate249inter1));
  and2  gate577(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate578(.a(s_4), .O(gate249inter3));
  inv1  gate579(.a(s_5), .O(gate249inter4));
  nand2 gate580(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate581(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate582(.a(G254), .O(gate249inter7));
  inv1  gate583(.a(G742), .O(gate249inter8));
  nand2 gate584(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate585(.a(s_5), .b(gate249inter3), .O(gate249inter10));
  nor2  gate586(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate587(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate588(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1947(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1948(.a(gate251inter0), .b(s_200), .O(gate251inter1));
  and2  gate1949(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1950(.a(s_200), .O(gate251inter3));
  inv1  gate1951(.a(s_201), .O(gate251inter4));
  nand2 gate1952(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1953(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1954(.a(G257), .O(gate251inter7));
  inv1  gate1955(.a(G745), .O(gate251inter8));
  nand2 gate1956(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1957(.a(s_201), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1958(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1959(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1960(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate2003(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2004(.a(gate252inter0), .b(s_208), .O(gate252inter1));
  and2  gate2005(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2006(.a(s_208), .O(gate252inter3));
  inv1  gate2007(.a(s_209), .O(gate252inter4));
  nand2 gate2008(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2009(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2010(.a(G709), .O(gate252inter7));
  inv1  gate2011(.a(G745), .O(gate252inter8));
  nand2 gate2012(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2013(.a(s_209), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2014(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2015(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2016(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2311(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2312(.a(gate264inter0), .b(s_252), .O(gate264inter1));
  and2  gate2313(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2314(.a(s_252), .O(gate264inter3));
  inv1  gate2315(.a(s_253), .O(gate264inter4));
  nand2 gate2316(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2317(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2318(.a(G768), .O(gate264inter7));
  inv1  gate2319(.a(G769), .O(gate264inter8));
  nand2 gate2320(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2321(.a(s_253), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2322(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2323(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2324(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate589(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate590(.a(gate267inter0), .b(s_6), .O(gate267inter1));
  and2  gate591(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate592(.a(s_6), .O(gate267inter3));
  inv1  gate593(.a(s_7), .O(gate267inter4));
  nand2 gate594(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate595(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate596(.a(G648), .O(gate267inter7));
  inv1  gate597(.a(G776), .O(gate267inter8));
  nand2 gate598(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate599(.a(s_7), .b(gate267inter3), .O(gate267inter10));
  nor2  gate600(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate601(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate602(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1835(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1836(.a(gate268inter0), .b(s_184), .O(gate268inter1));
  and2  gate1837(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1838(.a(s_184), .O(gate268inter3));
  inv1  gate1839(.a(s_185), .O(gate268inter4));
  nand2 gate1840(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1841(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1842(.a(G651), .O(gate268inter7));
  inv1  gate1843(.a(G779), .O(gate268inter8));
  nand2 gate1844(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1845(.a(s_185), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1846(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1847(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1848(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1191(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1192(.a(gate274inter0), .b(s_92), .O(gate274inter1));
  and2  gate1193(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1194(.a(s_92), .O(gate274inter3));
  inv1  gate1195(.a(s_93), .O(gate274inter4));
  nand2 gate1196(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1197(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1198(.a(G770), .O(gate274inter7));
  inv1  gate1199(.a(G794), .O(gate274inter8));
  nand2 gate1200(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1201(.a(s_93), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1202(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1203(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1204(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1821(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1822(.a(gate275inter0), .b(s_182), .O(gate275inter1));
  and2  gate1823(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1824(.a(s_182), .O(gate275inter3));
  inv1  gate1825(.a(s_183), .O(gate275inter4));
  nand2 gate1826(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1827(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1828(.a(G645), .O(gate275inter7));
  inv1  gate1829(.a(G797), .O(gate275inter8));
  nand2 gate1830(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1831(.a(s_183), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1832(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1833(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1834(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1891(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1892(.a(gate276inter0), .b(s_192), .O(gate276inter1));
  and2  gate1893(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1894(.a(s_192), .O(gate276inter3));
  inv1  gate1895(.a(s_193), .O(gate276inter4));
  nand2 gate1896(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1897(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1898(.a(G773), .O(gate276inter7));
  inv1  gate1899(.a(G797), .O(gate276inter8));
  nand2 gate1900(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1901(.a(s_193), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1902(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1903(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1904(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate827(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate828(.a(gate279inter0), .b(s_40), .O(gate279inter1));
  and2  gate829(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate830(.a(s_40), .O(gate279inter3));
  inv1  gate831(.a(s_41), .O(gate279inter4));
  nand2 gate832(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate833(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate834(.a(G651), .O(gate279inter7));
  inv1  gate835(.a(G803), .O(gate279inter8));
  nand2 gate836(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate837(.a(s_41), .b(gate279inter3), .O(gate279inter10));
  nor2  gate838(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate839(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate840(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1569(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1570(.a(gate283inter0), .b(s_146), .O(gate283inter1));
  and2  gate1571(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1572(.a(s_146), .O(gate283inter3));
  inv1  gate1573(.a(s_147), .O(gate283inter4));
  nand2 gate1574(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1575(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1576(.a(G657), .O(gate283inter7));
  inv1  gate1577(.a(G809), .O(gate283inter8));
  nand2 gate1578(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1579(.a(s_147), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1580(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1581(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1582(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2045(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2046(.a(gate287inter0), .b(s_214), .O(gate287inter1));
  and2  gate2047(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2048(.a(s_214), .O(gate287inter3));
  inv1  gate2049(.a(s_215), .O(gate287inter4));
  nand2 gate2050(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2051(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2052(.a(G663), .O(gate287inter7));
  inv1  gate2053(.a(G815), .O(gate287inter8));
  nand2 gate2054(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2055(.a(s_215), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2056(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2057(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2058(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1387(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1388(.a(gate288inter0), .b(s_120), .O(gate288inter1));
  and2  gate1389(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1390(.a(s_120), .O(gate288inter3));
  inv1  gate1391(.a(s_121), .O(gate288inter4));
  nand2 gate1392(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1393(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1394(.a(G791), .O(gate288inter7));
  inv1  gate1395(.a(G815), .O(gate288inter8));
  nand2 gate1396(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1397(.a(s_121), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1398(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1399(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1400(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1653(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1654(.a(gate289inter0), .b(s_158), .O(gate289inter1));
  and2  gate1655(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1656(.a(s_158), .O(gate289inter3));
  inv1  gate1657(.a(s_159), .O(gate289inter4));
  nand2 gate1658(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1659(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1660(.a(G818), .O(gate289inter7));
  inv1  gate1661(.a(G819), .O(gate289inter8));
  nand2 gate1662(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1663(.a(s_159), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1664(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1665(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1666(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1079(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1080(.a(gate290inter0), .b(s_76), .O(gate290inter1));
  and2  gate1081(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1082(.a(s_76), .O(gate290inter3));
  inv1  gate1083(.a(s_77), .O(gate290inter4));
  nand2 gate1084(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1085(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1086(.a(G820), .O(gate290inter7));
  inv1  gate1087(.a(G821), .O(gate290inter8));
  nand2 gate1088(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1089(.a(s_77), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1090(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1091(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1092(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1695(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1696(.a(gate292inter0), .b(s_164), .O(gate292inter1));
  and2  gate1697(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1698(.a(s_164), .O(gate292inter3));
  inv1  gate1699(.a(s_165), .O(gate292inter4));
  nand2 gate1700(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1701(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1702(.a(G824), .O(gate292inter7));
  inv1  gate1703(.a(G825), .O(gate292inter8));
  nand2 gate1704(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1705(.a(s_165), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1706(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1707(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1708(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1289(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1290(.a(gate294inter0), .b(s_106), .O(gate294inter1));
  and2  gate1291(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1292(.a(s_106), .O(gate294inter3));
  inv1  gate1293(.a(s_107), .O(gate294inter4));
  nand2 gate1294(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1295(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1296(.a(G832), .O(gate294inter7));
  inv1  gate1297(.a(G833), .O(gate294inter8));
  nand2 gate1298(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1299(.a(s_107), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1300(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1301(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1302(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1303(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1304(.a(gate296inter0), .b(s_108), .O(gate296inter1));
  and2  gate1305(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1306(.a(s_108), .O(gate296inter3));
  inv1  gate1307(.a(s_109), .O(gate296inter4));
  nand2 gate1308(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1309(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1310(.a(G826), .O(gate296inter7));
  inv1  gate1311(.a(G827), .O(gate296inter8));
  nand2 gate1312(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1313(.a(s_109), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1314(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1315(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1316(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1163(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1164(.a(gate387inter0), .b(s_88), .O(gate387inter1));
  and2  gate1165(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1166(.a(s_88), .O(gate387inter3));
  inv1  gate1167(.a(s_89), .O(gate387inter4));
  nand2 gate1168(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1169(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1170(.a(G1), .O(gate387inter7));
  inv1  gate1171(.a(G1036), .O(gate387inter8));
  nand2 gate1172(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1173(.a(s_89), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1174(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1175(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1176(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1261(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1262(.a(gate389inter0), .b(s_102), .O(gate389inter1));
  and2  gate1263(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1264(.a(s_102), .O(gate389inter3));
  inv1  gate1265(.a(s_103), .O(gate389inter4));
  nand2 gate1266(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1267(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1268(.a(G3), .O(gate389inter7));
  inv1  gate1269(.a(G1042), .O(gate389inter8));
  nand2 gate1270(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1271(.a(s_103), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1272(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1273(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1274(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate757(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate758(.a(gate390inter0), .b(s_30), .O(gate390inter1));
  and2  gate759(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate760(.a(s_30), .O(gate390inter3));
  inv1  gate761(.a(s_31), .O(gate390inter4));
  nand2 gate762(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate763(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate764(.a(G4), .O(gate390inter7));
  inv1  gate765(.a(G1045), .O(gate390inter8));
  nand2 gate766(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate767(.a(s_31), .b(gate390inter3), .O(gate390inter10));
  nor2  gate768(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate769(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate770(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1499(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1500(.a(gate393inter0), .b(s_136), .O(gate393inter1));
  and2  gate1501(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1502(.a(s_136), .O(gate393inter3));
  inv1  gate1503(.a(s_137), .O(gate393inter4));
  nand2 gate1504(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1505(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1506(.a(G7), .O(gate393inter7));
  inv1  gate1507(.a(G1054), .O(gate393inter8));
  nand2 gate1508(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1509(.a(s_137), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1510(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1511(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1512(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2171(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2172(.a(gate397inter0), .b(s_232), .O(gate397inter1));
  and2  gate2173(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2174(.a(s_232), .O(gate397inter3));
  inv1  gate2175(.a(s_233), .O(gate397inter4));
  nand2 gate2176(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2177(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2178(.a(G11), .O(gate397inter7));
  inv1  gate2179(.a(G1066), .O(gate397inter8));
  nand2 gate2180(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2181(.a(s_233), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2182(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2183(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2184(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1457(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1458(.a(gate398inter0), .b(s_130), .O(gate398inter1));
  and2  gate1459(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1460(.a(s_130), .O(gate398inter3));
  inv1  gate1461(.a(s_131), .O(gate398inter4));
  nand2 gate1462(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1463(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1464(.a(G12), .O(gate398inter7));
  inv1  gate1465(.a(G1069), .O(gate398inter8));
  nand2 gate1466(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1467(.a(s_131), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1468(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1469(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1470(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1247(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1248(.a(gate399inter0), .b(s_100), .O(gate399inter1));
  and2  gate1249(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1250(.a(s_100), .O(gate399inter3));
  inv1  gate1251(.a(s_101), .O(gate399inter4));
  nand2 gate1252(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1253(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1254(.a(G13), .O(gate399inter7));
  inv1  gate1255(.a(G1072), .O(gate399inter8));
  nand2 gate1256(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1257(.a(s_101), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1258(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1259(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1260(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2017(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2018(.a(gate400inter0), .b(s_210), .O(gate400inter1));
  and2  gate2019(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2020(.a(s_210), .O(gate400inter3));
  inv1  gate2021(.a(s_211), .O(gate400inter4));
  nand2 gate2022(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2023(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2024(.a(G14), .O(gate400inter7));
  inv1  gate2025(.a(G1075), .O(gate400inter8));
  nand2 gate2026(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2027(.a(s_211), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2028(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2029(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2030(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1583(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1584(.a(gate401inter0), .b(s_148), .O(gate401inter1));
  and2  gate1585(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1586(.a(s_148), .O(gate401inter3));
  inv1  gate1587(.a(s_149), .O(gate401inter4));
  nand2 gate1588(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1589(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1590(.a(G15), .O(gate401inter7));
  inv1  gate1591(.a(G1078), .O(gate401inter8));
  nand2 gate1592(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1593(.a(s_149), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1594(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1595(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1596(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1149(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1150(.a(gate404inter0), .b(s_86), .O(gate404inter1));
  and2  gate1151(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1152(.a(s_86), .O(gate404inter3));
  inv1  gate1153(.a(s_87), .O(gate404inter4));
  nand2 gate1154(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1155(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1156(.a(G18), .O(gate404inter7));
  inv1  gate1157(.a(G1087), .O(gate404inter8));
  nand2 gate1158(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1159(.a(s_87), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1160(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1161(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1162(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1205(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1206(.a(gate405inter0), .b(s_94), .O(gate405inter1));
  and2  gate1207(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1208(.a(s_94), .O(gate405inter3));
  inv1  gate1209(.a(s_95), .O(gate405inter4));
  nand2 gate1210(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1211(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1212(.a(G19), .O(gate405inter7));
  inv1  gate1213(.a(G1090), .O(gate405inter8));
  nand2 gate1214(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1215(.a(s_95), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1216(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1217(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1218(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1541(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1542(.a(gate408inter0), .b(s_142), .O(gate408inter1));
  and2  gate1543(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1544(.a(s_142), .O(gate408inter3));
  inv1  gate1545(.a(s_143), .O(gate408inter4));
  nand2 gate1546(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1547(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1548(.a(G22), .O(gate408inter7));
  inv1  gate1549(.a(G1099), .O(gate408inter8));
  nand2 gate1550(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1551(.a(s_143), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1552(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1553(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1554(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate617(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate618(.a(gate409inter0), .b(s_10), .O(gate409inter1));
  and2  gate619(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate620(.a(s_10), .O(gate409inter3));
  inv1  gate621(.a(s_11), .O(gate409inter4));
  nand2 gate622(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate623(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate624(.a(G23), .O(gate409inter7));
  inv1  gate625(.a(G1102), .O(gate409inter8));
  nand2 gate626(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate627(.a(s_11), .b(gate409inter3), .O(gate409inter10));
  nor2  gate628(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate629(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate630(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1681(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1682(.a(gate414inter0), .b(s_162), .O(gate414inter1));
  and2  gate1683(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1684(.a(s_162), .O(gate414inter3));
  inv1  gate1685(.a(s_163), .O(gate414inter4));
  nand2 gate1686(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1687(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1688(.a(G28), .O(gate414inter7));
  inv1  gate1689(.a(G1117), .O(gate414inter8));
  nand2 gate1690(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1691(.a(s_163), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1692(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1693(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1694(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate799(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate800(.a(gate418inter0), .b(s_36), .O(gate418inter1));
  and2  gate801(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate802(.a(s_36), .O(gate418inter3));
  inv1  gate803(.a(s_37), .O(gate418inter4));
  nand2 gate804(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate805(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate806(.a(G32), .O(gate418inter7));
  inv1  gate807(.a(G1129), .O(gate418inter8));
  nand2 gate808(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate809(.a(s_37), .b(gate418inter3), .O(gate418inter10));
  nor2  gate810(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate811(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate812(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate785(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate786(.a(gate419inter0), .b(s_34), .O(gate419inter1));
  and2  gate787(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate788(.a(s_34), .O(gate419inter3));
  inv1  gate789(.a(s_35), .O(gate419inter4));
  nand2 gate790(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate791(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate792(.a(G1), .O(gate419inter7));
  inv1  gate793(.a(G1132), .O(gate419inter8));
  nand2 gate794(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate795(.a(s_35), .b(gate419inter3), .O(gate419inter10));
  nor2  gate796(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate797(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate798(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1037(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1038(.a(gate421inter0), .b(s_70), .O(gate421inter1));
  and2  gate1039(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1040(.a(s_70), .O(gate421inter3));
  inv1  gate1041(.a(s_71), .O(gate421inter4));
  nand2 gate1042(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1043(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1044(.a(G2), .O(gate421inter7));
  inv1  gate1045(.a(G1135), .O(gate421inter8));
  nand2 gate1046(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1047(.a(s_71), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1048(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1049(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1050(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1961(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1962(.a(gate425inter0), .b(s_202), .O(gate425inter1));
  and2  gate1963(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1964(.a(s_202), .O(gate425inter3));
  inv1  gate1965(.a(s_203), .O(gate425inter4));
  nand2 gate1966(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1967(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1968(.a(G4), .O(gate425inter7));
  inv1  gate1969(.a(G1141), .O(gate425inter8));
  nand2 gate1970(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1971(.a(s_203), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1972(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1973(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1974(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate855(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate856(.a(gate432inter0), .b(s_44), .O(gate432inter1));
  and2  gate857(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate858(.a(s_44), .O(gate432inter3));
  inv1  gate859(.a(s_45), .O(gate432inter4));
  nand2 gate860(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate861(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate862(.a(G1054), .O(gate432inter7));
  inv1  gate863(.a(G1150), .O(gate432inter8));
  nand2 gate864(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate865(.a(s_45), .b(gate432inter3), .O(gate432inter10));
  nor2  gate866(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate867(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate868(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1709(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1710(.a(gate441inter0), .b(s_166), .O(gate441inter1));
  and2  gate1711(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1712(.a(s_166), .O(gate441inter3));
  inv1  gate1713(.a(s_167), .O(gate441inter4));
  nand2 gate1714(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1715(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1716(.a(G12), .O(gate441inter7));
  inv1  gate1717(.a(G1165), .O(gate441inter8));
  nand2 gate1718(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1719(.a(s_167), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1720(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1721(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1722(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate925(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate926(.a(gate452inter0), .b(s_54), .O(gate452inter1));
  and2  gate927(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate928(.a(s_54), .O(gate452inter3));
  inv1  gate929(.a(s_55), .O(gate452inter4));
  nand2 gate930(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate931(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate932(.a(G1084), .O(gate452inter7));
  inv1  gate933(.a(G1180), .O(gate452inter8));
  nand2 gate934(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate935(.a(s_55), .b(gate452inter3), .O(gate452inter10));
  nor2  gate936(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate937(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate938(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1093(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1094(.a(gate454inter0), .b(s_78), .O(gate454inter1));
  and2  gate1095(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1096(.a(s_78), .O(gate454inter3));
  inv1  gate1097(.a(s_79), .O(gate454inter4));
  nand2 gate1098(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1099(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1100(.a(G1087), .O(gate454inter7));
  inv1  gate1101(.a(G1183), .O(gate454inter8));
  nand2 gate1102(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1103(.a(s_79), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1104(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1105(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1106(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2269(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2270(.a(gate457inter0), .b(s_246), .O(gate457inter1));
  and2  gate2271(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2272(.a(s_246), .O(gate457inter3));
  inv1  gate2273(.a(s_247), .O(gate457inter4));
  nand2 gate2274(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2275(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2276(.a(G20), .O(gate457inter7));
  inv1  gate2277(.a(G1189), .O(gate457inter8));
  nand2 gate2278(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2279(.a(s_247), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2280(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2281(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2282(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1121(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1122(.a(gate459inter0), .b(s_82), .O(gate459inter1));
  and2  gate1123(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1124(.a(s_82), .O(gate459inter3));
  inv1  gate1125(.a(s_83), .O(gate459inter4));
  nand2 gate1126(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1127(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1128(.a(G21), .O(gate459inter7));
  inv1  gate1129(.a(G1192), .O(gate459inter8));
  nand2 gate1130(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1131(.a(s_83), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1132(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1133(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1134(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1723(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1724(.a(gate467inter0), .b(s_168), .O(gate467inter1));
  and2  gate1725(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1726(.a(s_168), .O(gate467inter3));
  inv1  gate1727(.a(s_169), .O(gate467inter4));
  nand2 gate1728(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1729(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1730(.a(G25), .O(gate467inter7));
  inv1  gate1731(.a(G1204), .O(gate467inter8));
  nand2 gate1732(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1733(.a(s_169), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1734(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1735(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1736(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1849(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1850(.a(gate468inter0), .b(s_186), .O(gate468inter1));
  and2  gate1851(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1852(.a(s_186), .O(gate468inter3));
  inv1  gate1853(.a(s_187), .O(gate468inter4));
  nand2 gate1854(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1855(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1856(.a(G1108), .O(gate468inter7));
  inv1  gate1857(.a(G1204), .O(gate468inter8));
  nand2 gate1858(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1859(.a(s_187), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1860(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1861(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1862(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate729(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate730(.a(gate469inter0), .b(s_26), .O(gate469inter1));
  and2  gate731(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate732(.a(s_26), .O(gate469inter3));
  inv1  gate733(.a(s_27), .O(gate469inter4));
  nand2 gate734(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate735(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate736(.a(G26), .O(gate469inter7));
  inv1  gate737(.a(G1207), .O(gate469inter8));
  nand2 gate738(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate739(.a(s_27), .b(gate469inter3), .O(gate469inter10));
  nor2  gate740(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate741(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate742(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate897(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate898(.a(gate474inter0), .b(s_50), .O(gate474inter1));
  and2  gate899(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate900(.a(s_50), .O(gate474inter3));
  inv1  gate901(.a(s_51), .O(gate474inter4));
  nand2 gate902(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate903(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate904(.a(G1117), .O(gate474inter7));
  inv1  gate905(.a(G1213), .O(gate474inter8));
  nand2 gate906(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate907(.a(s_51), .b(gate474inter3), .O(gate474inter10));
  nor2  gate908(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate909(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate910(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1485(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1486(.a(gate478inter0), .b(s_134), .O(gate478inter1));
  and2  gate1487(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1488(.a(s_134), .O(gate478inter3));
  inv1  gate1489(.a(s_135), .O(gate478inter4));
  nand2 gate1490(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1491(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1492(.a(G1123), .O(gate478inter7));
  inv1  gate1493(.a(G1219), .O(gate478inter8));
  nand2 gate1494(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1495(.a(s_135), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1496(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1497(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1498(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2115(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2116(.a(gate479inter0), .b(s_224), .O(gate479inter1));
  and2  gate2117(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2118(.a(s_224), .O(gate479inter3));
  inv1  gate2119(.a(s_225), .O(gate479inter4));
  nand2 gate2120(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2121(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2122(.a(G31), .O(gate479inter7));
  inv1  gate2123(.a(G1222), .O(gate479inter8));
  nand2 gate2124(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2125(.a(s_225), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2126(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2127(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2128(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1135(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1136(.a(gate481inter0), .b(s_84), .O(gate481inter1));
  and2  gate1137(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1138(.a(s_84), .O(gate481inter3));
  inv1  gate1139(.a(s_85), .O(gate481inter4));
  nand2 gate1140(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1141(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1142(.a(G32), .O(gate481inter7));
  inv1  gate1143(.a(G1225), .O(gate481inter8));
  nand2 gate1144(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1145(.a(s_85), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1146(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1147(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1148(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1177(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1178(.a(gate482inter0), .b(s_90), .O(gate482inter1));
  and2  gate1179(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1180(.a(s_90), .O(gate482inter3));
  inv1  gate1181(.a(s_91), .O(gate482inter4));
  nand2 gate1182(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1183(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1184(.a(G1129), .O(gate482inter7));
  inv1  gate1185(.a(G1225), .O(gate482inter8));
  nand2 gate1186(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1187(.a(s_91), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1188(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1189(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1190(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1639(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1640(.a(gate483inter0), .b(s_156), .O(gate483inter1));
  and2  gate1641(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1642(.a(s_156), .O(gate483inter3));
  inv1  gate1643(.a(s_157), .O(gate483inter4));
  nand2 gate1644(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1645(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1646(.a(G1228), .O(gate483inter7));
  inv1  gate1647(.a(G1229), .O(gate483inter8));
  nand2 gate1648(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1649(.a(s_157), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1650(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1651(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1652(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1219(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1220(.a(gate484inter0), .b(s_96), .O(gate484inter1));
  and2  gate1221(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1222(.a(s_96), .O(gate484inter3));
  inv1  gate1223(.a(s_97), .O(gate484inter4));
  nand2 gate1224(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1225(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1226(.a(G1230), .O(gate484inter7));
  inv1  gate1227(.a(G1231), .O(gate484inter8));
  nand2 gate1228(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1229(.a(s_97), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1230(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1231(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1232(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1667(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1668(.a(gate490inter0), .b(s_160), .O(gate490inter1));
  and2  gate1669(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1670(.a(s_160), .O(gate490inter3));
  inv1  gate1671(.a(s_161), .O(gate490inter4));
  nand2 gate1672(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1673(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1674(.a(G1242), .O(gate490inter7));
  inv1  gate1675(.a(G1243), .O(gate490inter8));
  nand2 gate1676(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1677(.a(s_161), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1678(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1679(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1680(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1345(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1346(.a(gate491inter0), .b(s_114), .O(gate491inter1));
  and2  gate1347(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1348(.a(s_114), .O(gate491inter3));
  inv1  gate1349(.a(s_115), .O(gate491inter4));
  nand2 gate1350(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1351(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1352(.a(G1244), .O(gate491inter7));
  inv1  gate1353(.a(G1245), .O(gate491inter8));
  nand2 gate1354(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1355(.a(s_115), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1356(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1357(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1358(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1401(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1402(.a(gate494inter0), .b(s_122), .O(gate494inter1));
  and2  gate1403(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1404(.a(s_122), .O(gate494inter3));
  inv1  gate1405(.a(s_123), .O(gate494inter4));
  nand2 gate1406(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1407(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1408(.a(G1250), .O(gate494inter7));
  inv1  gate1409(.a(G1251), .O(gate494inter8));
  nand2 gate1410(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1411(.a(s_123), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1412(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1413(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1414(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate911(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate912(.a(gate496inter0), .b(s_52), .O(gate496inter1));
  and2  gate913(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate914(.a(s_52), .O(gate496inter3));
  inv1  gate915(.a(s_53), .O(gate496inter4));
  nand2 gate916(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate917(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate918(.a(G1254), .O(gate496inter7));
  inv1  gate919(.a(G1255), .O(gate496inter8));
  nand2 gate920(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate921(.a(s_53), .b(gate496inter3), .O(gate496inter10));
  nor2  gate922(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate923(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate924(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1597(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1598(.a(gate497inter0), .b(s_150), .O(gate497inter1));
  and2  gate1599(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1600(.a(s_150), .O(gate497inter3));
  inv1  gate1601(.a(s_151), .O(gate497inter4));
  nand2 gate1602(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1603(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1604(.a(G1256), .O(gate497inter7));
  inv1  gate1605(.a(G1257), .O(gate497inter8));
  nand2 gate1606(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1607(.a(s_151), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1608(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1609(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1610(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1877(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1878(.a(gate499inter0), .b(s_190), .O(gate499inter1));
  and2  gate1879(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1880(.a(s_190), .O(gate499inter3));
  inv1  gate1881(.a(s_191), .O(gate499inter4));
  nand2 gate1882(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1883(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1884(.a(G1260), .O(gate499inter7));
  inv1  gate1885(.a(G1261), .O(gate499inter8));
  nand2 gate1886(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1887(.a(s_191), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1888(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1889(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1890(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate939(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate940(.a(gate502inter0), .b(s_56), .O(gate502inter1));
  and2  gate941(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate942(.a(s_56), .O(gate502inter3));
  inv1  gate943(.a(s_57), .O(gate502inter4));
  nand2 gate944(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate945(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate946(.a(G1266), .O(gate502inter7));
  inv1  gate947(.a(G1267), .O(gate502inter8));
  nand2 gate948(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate949(.a(s_57), .b(gate502inter3), .O(gate502inter10));
  nor2  gate950(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate951(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate952(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate547(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate548(.a(gate509inter0), .b(s_0), .O(gate509inter1));
  and2  gate549(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate550(.a(s_0), .O(gate509inter3));
  inv1  gate551(.a(s_1), .O(gate509inter4));
  nand2 gate552(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate553(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate554(.a(G1280), .O(gate509inter7));
  inv1  gate555(.a(G1281), .O(gate509inter8));
  nand2 gate556(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate557(.a(s_1), .b(gate509inter3), .O(gate509inter10));
  nor2  gate558(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate559(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate560(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule