module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;
wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate310inter0, gate310inter1, gate310inter2, gate310inter3, gate310inter4, gate310inter5, gate310inter6, gate310inter7, gate310inter8, gate310inter9, gate310inter10, gate310inter11, gate310inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate333inter0, gate333inter1, gate333inter2, gate333inter3, gate333inter4, gate333inter5, gate333inter6, gate333inter7, gate333inter8, gate333inter9, gate333inter10, gate333inter11, gate333inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12;


nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );

  xor2  gate678(.a(N68), .b(N29), .O(gate8inter0));
  nand2 gate679(.a(gate8inter0), .b(s_42), .O(gate8inter1));
  and2  gate680(.a(N68), .b(N29), .O(gate8inter2));
  inv1  gate681(.a(s_42), .O(gate8inter3));
  inv1  gate682(.a(s_43), .O(gate8inter4));
  nand2 gate683(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate684(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate685(.a(N29), .O(gate8inter7));
  inv1  gate686(.a(N68), .O(gate8inter8));
  nand2 gate687(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate688(.a(s_43), .b(gate8inter3), .O(gate8inter10));
  nor2  gate689(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate690(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate691(.a(gate8inter12), .b(gate8inter1), .O(N285));
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );
nand2 gate20( .a(N91), .b(N96), .O(N301) );
or2 gate21( .a(N91), .b(N96), .O(N302) );
nand2 gate22( .a(N101), .b(N106), .O(N303) );
or2 gate23( .a(N101), .b(N106), .O(N304) );
nand2 gate24( .a(N111), .b(N116), .O(N305) );
or2 gate25( .a(N111), .b(N116), .O(N306) );
nand2 gate26( .a(N121), .b(N126), .O(N307) );
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );
nand2 gate33( .a(N59), .b(N156), .O(N319) );
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17), .b(N42), .O(N323) );
nand2 gate36( .a(N159), .b(N165), .O(N324) );
or2 gate37( .a(N159), .b(N165), .O(N325) );
nand2 gate38( .a(N171), .b(N177), .O(N326) );
or2 gate39( .a(N171), .b(N177), .O(N327) );
nand2 gate40( .a(N183), .b(N189), .O(N328) );
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
and2 gate49( .a(N255), .b(N259), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );
nor2 gate60( .a(N280), .b(N284), .O(N348) );
or2 gate61( .a(N280), .b(N285), .O(N349) );
or2 gate62( .a(N280), .b(N286), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );

  xor2  gate664(.a(N298), .b(N89), .O(gate67inter0));
  nand2 gate665(.a(gate67inter0), .b(s_40), .O(gate67inter1));
  and2  gate666(.a(N298), .b(N89), .O(gate67inter2));
  inv1  gate667(.a(s_40), .O(gate67inter3));
  inv1  gate668(.a(s_41), .O(gate67inter4));
  nand2 gate669(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate670(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate671(.a(N89), .O(gate67inter7));
  inv1  gate672(.a(N298), .O(gate67inter8));
  nand2 gate673(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate674(.a(s_41), .b(gate67inter3), .O(gate67inter10));
  nor2  gate675(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate676(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate677(.a(gate67inter12), .b(gate67inter1), .O(N355));
and2 gate68( .a(N90), .b(N298), .O(N356) );

  xor2  gate734(.a(N302), .b(N301), .O(gate69inter0));
  nand2 gate735(.a(gate69inter0), .b(s_50), .O(gate69inter1));
  and2  gate736(.a(N302), .b(N301), .O(gate69inter2));
  inv1  gate737(.a(s_50), .O(gate69inter3));
  inv1  gate738(.a(s_51), .O(gate69inter4));
  nand2 gate739(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate740(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate741(.a(N301), .O(gate69inter7));
  inv1  gate742(.a(N302), .O(gate69inter8));
  nand2 gate743(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate744(.a(s_51), .b(gate69inter3), .O(gate69inter10));
  nor2  gate745(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate746(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate747(.a(gate69inter12), .b(gate69inter1), .O(N357));
nand2 gate70( .a(N303), .b(N304), .O(N360) );
nand2 gate71( .a(N305), .b(N306), .O(N363) );

  xor2  gate762(.a(N308), .b(N307), .O(gate72inter0));
  nand2 gate763(.a(gate72inter0), .b(s_54), .O(gate72inter1));
  and2  gate764(.a(N308), .b(N307), .O(gate72inter2));
  inv1  gate765(.a(s_54), .O(gate72inter3));
  inv1  gate766(.a(s_55), .O(gate72inter4));
  nand2 gate767(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate768(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate769(.a(N307), .O(gate72inter7));
  inv1  gate770(.a(N308), .O(gate72inter8));
  nand2 gate771(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate772(.a(s_55), .b(gate72inter3), .O(gate72inter10));
  nor2  gate773(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate774(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate775(.a(gate72inter12), .b(gate72inter1), .O(N366));
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );
nand2 gate76( .a(N326), .b(N327), .O(N379) );

  xor2  gate636(.a(N329), .b(N328), .O(gate77inter0));
  nand2 gate637(.a(gate77inter0), .b(s_36), .O(gate77inter1));
  and2  gate638(.a(N329), .b(N328), .O(gate77inter2));
  inv1  gate639(.a(s_36), .O(gate77inter3));
  inv1  gate640(.a(s_37), .O(gate77inter4));
  nand2 gate641(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate642(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate643(.a(N328), .O(gate77inter7));
  inv1  gate644(.a(N329), .O(gate77inter8));
  nand2 gate645(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate646(.a(s_37), .b(gate77inter3), .O(gate77inter10));
  nor2  gate647(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate648(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate649(.a(gate77inter12), .b(gate77inter1), .O(N382));
nand2 gate78( .a(N330), .b(N331), .O(N385) );
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );

  xor2  gate790(.a(N352), .b(N347), .O(gate96inter0));
  nand2 gate791(.a(gate96inter0), .b(s_58), .O(gate96inter1));
  and2  gate792(.a(N352), .b(N347), .O(gate96inter2));
  inv1  gate793(.a(s_58), .O(gate96inter3));
  inv1  gate794(.a(s_59), .O(gate96inter4));
  nand2 gate795(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate796(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate797(.a(N347), .O(gate96inter7));
  inv1  gate798(.a(N352), .O(gate96inter8));
  nand2 gate799(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate800(.a(s_59), .b(gate96inter3), .O(gate96inter10));
  nor2  gate801(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate802(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate803(.a(gate96inter12), .b(gate96inter1), .O(N410));
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );
nor2 gate126( .a(N406), .b(N425), .O(N460) );

  xor2  gate384(.a(N426), .b(N409), .O(gate127inter0));
  nand2 gate385(.a(gate127inter0), .b(s_0), .O(gate127inter1));
  and2  gate386(.a(N426), .b(N409), .O(gate127inter2));
  inv1  gate387(.a(s_0), .O(gate127inter3));
  inv1  gate388(.a(s_1), .O(gate127inter4));
  nand2 gate389(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate390(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate391(.a(N409), .O(gate127inter7));
  inv1  gate392(.a(N426), .O(gate127inter8));
  nand2 gate393(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate394(.a(s_1), .b(gate127inter3), .O(gate127inter10));
  nor2  gate395(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate396(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate397(.a(gate127inter12), .b(gate127inter1), .O(N463));
nand2 gate128( .a(N442), .b(N410), .O(N466) );
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );
nand2 gate137( .a(N443), .b(N1), .O(N483) );
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );
nor2 gate142( .a(N413), .b(N444), .O(N492) );
nor2 gate143( .a(N416), .b(N445), .O(N495) );

  xor2  gate426(.a(N460), .b(N130), .O(gate144inter0));
  nand2 gate427(.a(gate144inter0), .b(s_6), .O(gate144inter1));
  and2  gate428(.a(N460), .b(N130), .O(gate144inter2));
  inv1  gate429(.a(s_6), .O(gate144inter3));
  inv1  gate430(.a(s_7), .O(gate144inter4));
  nand2 gate431(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate432(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate433(.a(N130), .O(gate144inter7));
  inv1  gate434(.a(N460), .O(gate144inter8));
  nand2 gate435(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate436(.a(s_7), .b(gate144inter3), .O(gate144inter10));
  nor2  gate437(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate438(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate439(.a(gate144inter12), .b(gate144inter1), .O(N498));
or2 gate145( .a(N130), .b(N460), .O(N499) );
nand2 gate146( .a(N463), .b(N135), .O(N500) );
or2 gate147( .a(N463), .b(N135), .O(N501) );
and2 gate148( .a(N91), .b(N466), .O(N502) );
nor2 gate149( .a(N475), .b(N476), .O(N503) );
and2 gate150( .a(N96), .b(N466), .O(N504) );
nor2 gate151( .a(N477), .b(N478), .O(N505) );
and2 gate152( .a(N101), .b(N466), .O(N506) );
nor2 gate153( .a(N479), .b(N480), .O(N507) );
and2 gate154( .a(N106), .b(N466), .O(N508) );
nor2 gate155( .a(N481), .b(N482), .O(N509) );
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );

  xor2  gate510(.a(N492), .b(N130), .O(gate164inter0));
  nand2 gate511(.a(gate164inter0), .b(s_18), .O(gate164inter1));
  and2  gate512(.a(N492), .b(N130), .O(gate164inter2));
  inv1  gate513(.a(s_18), .O(gate164inter3));
  inv1  gate514(.a(s_19), .O(gate164inter4));
  nand2 gate515(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate516(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate517(.a(N130), .O(gate164inter7));
  inv1  gate518(.a(N492), .O(gate164inter8));
  nand2 gate519(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate520(.a(s_19), .b(gate164inter3), .O(gate164inter10));
  nor2  gate521(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate522(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate523(.a(gate164inter12), .b(gate164inter1), .O(N518));
or2 gate165( .a(N130), .b(N492), .O(N519) );
nand2 gate166( .a(N495), .b(N207), .O(N520) );
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
and2 gate170( .a(N451), .b(N171), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );
nand2 gate173( .a(N451), .b(N189), .O(N527) );
nand2 gate174( .a(N451), .b(N195), .O(N528) );
nand2 gate175( .a(N451), .b(N201), .O(N529) );

  xor2  gate832(.a(N499), .b(N498), .O(gate176inter0));
  nand2 gate833(.a(gate176inter0), .b(s_64), .O(gate176inter1));
  and2  gate834(.a(N499), .b(N498), .O(gate176inter2));
  inv1  gate835(.a(s_64), .O(gate176inter3));
  inv1  gate836(.a(s_65), .O(gate176inter4));
  nand2 gate837(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate838(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate839(.a(N498), .O(gate176inter7));
  inv1  gate840(.a(N499), .O(gate176inter8));
  nand2 gate841(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate842(.a(s_65), .b(gate176inter3), .O(gate176inter10));
  nor2  gate843(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate844(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate845(.a(gate176inter12), .b(gate176inter1), .O(N530));
nand2 gate177( .a(N500), .b(N501), .O(N533) );
nor2 gate178( .a(N309), .b(N502), .O(N536) );
nor2 gate179( .a(N316), .b(N504), .O(N537) );

  xor2  gate440(.a(N506), .b(N317), .O(gate180inter0));
  nand2 gate441(.a(gate180inter0), .b(s_8), .O(gate180inter1));
  and2  gate442(.a(N506), .b(N317), .O(gate180inter2));
  inv1  gate443(.a(s_8), .O(gate180inter3));
  inv1  gate444(.a(s_9), .O(gate180inter4));
  nand2 gate445(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate446(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate447(.a(N317), .O(gate180inter7));
  inv1  gate448(.a(N506), .O(gate180inter8));
  nand2 gate449(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate450(.a(s_9), .b(gate180inter3), .O(gate180inter10));
  nor2  gate451(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate452(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate453(.a(gate180inter12), .b(gate180inter1), .O(N538));
nor2 gate181( .a(N318), .b(N508), .O(N539) );

  xor2  gate706(.a(N511), .b(N510), .O(gate182inter0));
  nand2 gate707(.a(gate182inter0), .b(s_46), .O(gate182inter1));
  and2  gate708(.a(N511), .b(N510), .O(gate182inter2));
  inv1  gate709(.a(s_46), .O(gate182inter3));
  inv1  gate710(.a(s_47), .O(gate182inter4));
  nand2 gate711(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate712(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate713(.a(N510), .O(gate182inter7));
  inv1  gate714(.a(N511), .O(gate182inter8));
  nand2 gate715(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate716(.a(s_47), .b(gate182inter3), .O(gate182inter10));
  nor2  gate717(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate718(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate719(.a(gate182inter12), .b(gate182inter1), .O(N540));

  xor2  gate608(.a(N513), .b(N512), .O(gate183inter0));
  nand2 gate609(.a(gate183inter0), .b(s_32), .O(gate183inter1));
  and2  gate610(.a(N513), .b(N512), .O(gate183inter2));
  inv1  gate611(.a(s_32), .O(gate183inter3));
  inv1  gate612(.a(s_33), .O(gate183inter4));
  nand2 gate613(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate614(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate615(.a(N512), .O(gate183inter7));
  inv1  gate616(.a(N513), .O(gate183inter8));
  nand2 gate617(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate618(.a(s_33), .b(gate183inter3), .O(gate183inter10));
  nor2  gate619(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate620(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate621(.a(gate183inter12), .b(gate183inter1), .O(N541));
nor2 gate184( .a(N514), .b(N515), .O(N542) );

  xor2  gate846(.a(N517), .b(N516), .O(gate185inter0));
  nand2 gate847(.a(gate185inter0), .b(s_66), .O(gate185inter1));
  and2  gate848(.a(N517), .b(N516), .O(gate185inter2));
  inv1  gate849(.a(s_66), .O(gate185inter3));
  inv1  gate850(.a(s_67), .O(gate185inter4));
  nand2 gate851(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate852(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate853(.a(N516), .O(gate185inter7));
  inv1  gate854(.a(N517), .O(gate185inter8));
  nand2 gate855(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate856(.a(s_67), .b(gate185inter3), .O(gate185inter10));
  nor2  gate857(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate858(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate859(.a(gate185inter12), .b(gate185inter1), .O(N543));
nand2 gate186( .a(N518), .b(N519), .O(N544) );
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );

  xor2  gate482(.a(N503), .b(N536), .O(gate191inter0));
  nand2 gate483(.a(gate191inter0), .b(s_14), .O(gate191inter1));
  and2  gate484(.a(N503), .b(N536), .O(gate191inter2));
  inv1  gate485(.a(s_14), .O(gate191inter3));
  inv1  gate486(.a(s_15), .O(gate191inter4));
  nand2 gate487(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate488(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate489(.a(N536), .O(gate191inter7));
  inv1  gate490(.a(N503), .O(gate191inter8));
  nand2 gate491(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate492(.a(s_15), .b(gate191inter3), .O(gate191inter10));
  nor2  gate493(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate494(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate495(.a(gate191inter12), .b(gate191inter1), .O(N553));
nand2 gate192( .a(N537), .b(N505), .O(N557) );

  xor2  gate874(.a(N507), .b(N538), .O(gate193inter0));
  nand2 gate875(.a(gate193inter0), .b(s_70), .O(gate193inter1));
  and2  gate876(.a(N507), .b(N538), .O(gate193inter2));
  inv1  gate877(.a(s_70), .O(gate193inter3));
  inv1  gate878(.a(s_71), .O(gate193inter4));
  nand2 gate879(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate880(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate881(.a(N538), .O(gate193inter7));
  inv1  gate882(.a(N507), .O(gate193inter8));
  nand2 gate883(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate884(.a(s_71), .b(gate193inter3), .O(gate193inter10));
  nor2  gate885(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate886(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate887(.a(gate193inter12), .b(gate193inter1), .O(N561));
nand2 gate194( .a(N539), .b(N509), .O(N565) );
nand2 gate195( .a(N488), .b(N540), .O(N569) );
nand2 gate196( .a(N489), .b(N541), .O(N573) );

  xor2  gate748(.a(N542), .b(N490), .O(gate197inter0));
  nand2 gate749(.a(gate197inter0), .b(s_52), .O(gate197inter1));
  and2  gate750(.a(N542), .b(N490), .O(gate197inter2));
  inv1  gate751(.a(s_52), .O(gate197inter3));
  inv1  gate752(.a(s_53), .O(gate197inter4));
  nand2 gate753(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate754(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate755(.a(N490), .O(gate197inter7));
  inv1  gate756(.a(N542), .O(gate197inter8));
  nand2 gate757(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate758(.a(s_53), .b(gate197inter3), .O(gate197inter10));
  nor2  gate759(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate760(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate761(.a(gate197inter12), .b(gate197inter1), .O(N577));
nand2 gate198( .a(N491), .b(N543), .O(N581) );
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );

  xor2  gate496(.a(N159), .b(N553), .O(gate204inter0));
  nand2 gate497(.a(gate204inter0), .b(s_16), .O(gate204inter1));
  and2  gate498(.a(N159), .b(N553), .O(gate204inter2));
  inv1  gate499(.a(s_16), .O(gate204inter3));
  inv1  gate500(.a(s_17), .O(gate204inter4));
  nand2 gate501(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate502(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate503(.a(N553), .O(gate204inter7));
  inv1  gate504(.a(N159), .O(gate204inter8));
  nand2 gate505(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate506(.a(s_17), .b(gate204inter3), .O(gate204inter10));
  nor2  gate507(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate508(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate509(.a(gate204inter12), .b(gate204inter1), .O(N590));
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );

  xor2  gate818(.a(N165), .b(N557), .O(gate207inter0));
  nand2 gate819(.a(gate207inter0), .b(s_62), .O(gate207inter1));
  and2  gate820(.a(N165), .b(N557), .O(gate207inter2));
  inv1  gate821(.a(s_62), .O(gate207inter3));
  inv1  gate822(.a(s_63), .O(gate207inter4));
  nand2 gate823(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate824(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate825(.a(N557), .O(gate207inter7));
  inv1  gate826(.a(N165), .O(gate207inter8));
  nand2 gate827(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate828(.a(s_63), .b(gate207inter3), .O(gate207inter10));
  nor2  gate829(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate830(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate831(.a(gate207inter12), .b(gate207inter1), .O(N597));
or2 gate208( .a(N557), .b(N165), .O(N600) );
and2 gate209( .a(N246), .b(N557), .O(N605) );

  xor2  gate538(.a(N171), .b(N561), .O(gate210inter0));
  nand2 gate539(.a(gate210inter0), .b(s_22), .O(gate210inter1));
  and2  gate540(.a(N171), .b(N561), .O(gate210inter2));
  inv1  gate541(.a(s_22), .O(gate210inter3));
  inv1  gate542(.a(s_23), .O(gate210inter4));
  nand2 gate543(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate544(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate545(.a(N561), .O(gate210inter7));
  inv1  gate546(.a(N171), .O(gate210inter8));
  nand2 gate547(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate548(.a(s_23), .b(gate210inter3), .O(gate210inter10));
  nor2  gate549(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate550(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate551(.a(gate210inter12), .b(gate210inter1), .O(N606));
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );
nand2 gate213( .a(N565), .b(N177), .O(N616) );
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );

  xor2  gate454(.a(N183), .b(N569), .O(gate216inter0));
  nand2 gate455(.a(gate216inter0), .b(s_10), .O(gate216inter1));
  and2  gate456(.a(N183), .b(N569), .O(gate216inter2));
  inv1  gate457(.a(s_10), .O(gate216inter3));
  inv1  gate458(.a(s_11), .O(gate216inter4));
  nand2 gate459(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate460(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate461(.a(N569), .O(gate216inter7));
  inv1  gate462(.a(N183), .O(gate216inter8));
  nand2 gate463(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate464(.a(s_11), .b(gate216inter3), .O(gate216inter10));
  nor2  gate465(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate466(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate467(.a(gate216inter12), .b(gate216inter1), .O(N625));
or2 gate217( .a(N569), .b(N183), .O(N628) );
and2 gate218( .a(N246), .b(N569), .O(N631) );

  xor2  gate594(.a(N189), .b(N573), .O(gate219inter0));
  nand2 gate595(.a(gate219inter0), .b(s_30), .O(gate219inter1));
  and2  gate596(.a(N189), .b(N573), .O(gate219inter2));
  inv1  gate597(.a(s_30), .O(gate219inter3));
  inv1  gate598(.a(s_31), .O(gate219inter4));
  nand2 gate599(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate600(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate601(.a(N573), .O(gate219inter7));
  inv1  gate602(.a(N189), .O(gate219inter8));
  nand2 gate603(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate604(.a(s_31), .b(gate219inter3), .O(gate219inter10));
  nor2  gate605(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate606(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate607(.a(gate219inter12), .b(gate219inter1), .O(N632));
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );

  xor2  gate650(.a(N195), .b(N577), .O(gate222inter0));
  nand2 gate651(.a(gate222inter0), .b(s_38), .O(gate222inter1));
  and2  gate652(.a(N195), .b(N577), .O(gate222inter2));
  inv1  gate653(.a(s_38), .O(gate222inter3));
  inv1  gate654(.a(s_39), .O(gate222inter4));
  nand2 gate655(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate656(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate657(.a(N577), .O(gate222inter7));
  inv1  gate658(.a(N195), .O(gate222inter8));
  nand2 gate659(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate660(.a(s_39), .b(gate222inter3), .O(gate222inter10));
  nor2  gate661(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate662(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate663(.a(gate222inter12), .b(gate222inter1), .O(N641));
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );
nand2 gate225( .a(N581), .b(N201), .O(N651) );
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );
nor2 gate228( .a(N552), .b(N588), .O(N660) );
nor2 gate229( .a(N587), .b(N589), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
and2 gate231( .a(N593), .b(N590), .O(N665) );
nor2 gate232( .a(N596), .b(N522), .O(N669) );
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );
nor2 gate235( .a(N605), .b(N523), .O(N677) );
inv1 gate236( .a(N606), .O(N678) );
and2 gate237( .a(N609), .b(N606), .O(N682) );
nor2 gate238( .a(N615), .b(N524), .O(N686) );
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );

  xor2  gate692(.a(N525), .b(N624), .O(gate241inter0));
  nand2 gate693(.a(gate241inter0), .b(s_44), .O(gate241inter1));
  and2  gate694(.a(N525), .b(N624), .O(gate241inter2));
  inv1  gate695(.a(s_44), .O(gate241inter3));
  inv1  gate696(.a(s_45), .O(gate241inter4));
  nand2 gate697(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate698(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate699(.a(N624), .O(gate241inter7));
  inv1  gate700(.a(N525), .O(gate241inter8));
  nand2 gate701(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate702(.a(s_45), .b(gate241inter3), .O(gate241inter10));
  nor2  gate703(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate704(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate705(.a(gate241inter12), .b(gate241inter1), .O(N696));
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );
nor2 gate244( .a(N631), .b(N526), .O(N704) );
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );

  xor2  gate552(.a(N640), .b(N337), .O(gate247inter0));
  nand2 gate553(.a(gate247inter0), .b(s_24), .O(gate247inter1));
  and2  gate554(.a(N640), .b(N337), .O(gate247inter2));
  inv1  gate555(.a(s_24), .O(gate247inter3));
  inv1  gate556(.a(s_25), .O(gate247inter4));
  nand2 gate557(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate558(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate559(.a(N337), .O(gate247inter7));
  inv1  gate560(.a(N640), .O(gate247inter8));
  nand2 gate561(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate562(.a(s_25), .b(gate247inter3), .O(gate247inter10));
  nor2  gate563(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate564(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate565(.a(gate247inter12), .b(gate247inter1), .O(N712));
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );

  xor2  gate720(.a(N650), .b(N339), .O(gate250inter0));
  nand2 gate721(.a(gate250inter0), .b(s_48), .O(gate250inter1));
  and2  gate722(.a(N650), .b(N339), .O(gate250inter2));
  inv1  gate723(.a(s_48), .O(gate250inter3));
  inv1  gate724(.a(s_49), .O(gate250inter4));
  nand2 gate725(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate726(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate727(.a(N339), .O(gate250inter7));
  inv1  gate728(.a(N650), .O(gate250inter8));
  nand2 gate729(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate730(.a(s_49), .b(gate250inter3), .O(gate250inter10));
  nor2  gate731(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate732(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate733(.a(gate250inter12), .b(gate250inter1), .O(N721));
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );

  xor2  gate580(.a(N659), .b(N341), .O(gate253inter0));
  nand2 gate581(.a(gate253inter0), .b(s_28), .O(gate253inter1));
  and2  gate582(.a(N659), .b(N341), .O(gate253inter2));
  inv1  gate583(.a(s_28), .O(gate253inter3));
  inv1  gate584(.a(s_29), .O(gate253inter4));
  nand2 gate585(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate586(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate587(.a(N341), .O(gate253inter7));
  inv1  gate588(.a(N659), .O(gate253inter8));
  nand2 gate589(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate590(.a(s_29), .b(gate253inter3), .O(gate253inter10));
  nor2  gate591(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate592(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate593(.a(gate253inter12), .b(gate253inter1), .O(N731));
nand2 gate254( .a(N654), .b(N261), .O(N732) );
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
and2 gate273( .a(N228), .b(N708), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );

  xor2  gate776(.a(N261), .b(N727), .O(gate279inter0));
  nand2 gate777(.a(gate279inter0), .b(s_56), .O(gate279inter1));
  and2  gate778(.a(N261), .b(N727), .O(gate279inter2));
  inv1  gate779(.a(s_56), .O(gate279inter3));
  inv1  gate780(.a(s_57), .O(gate279inter4));
  nand2 gate781(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate782(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate783(.a(N727), .O(gate279inter7));
  inv1  gate784(.a(N261), .O(gate279inter8));
  nand2 gate785(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate786(.a(s_57), .b(gate279inter3), .O(gate279inter10));
  nor2  gate787(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate788(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate789(.a(gate279inter12), .b(gate279inter1), .O(N757));
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );
nand2 gate284( .a(N635), .b(N713), .O(N762) );
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );

  xor2  gate622(.a(N737), .b(N736), .O(gate291inter0));
  nand2 gate623(.a(gate291inter0), .b(s_34), .O(gate291inter1));
  and2  gate624(.a(N737), .b(N736), .O(gate291inter2));
  inv1  gate625(.a(s_34), .O(gate291inter3));
  inv1  gate626(.a(s_35), .O(gate291inter4));
  nand2 gate627(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate628(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate629(.a(N736), .O(gate291inter7));
  inv1  gate630(.a(N737), .O(gate291inter8));
  nand2 gate631(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate632(.a(s_35), .b(gate291inter3), .O(gate291inter10));
  nor2  gate633(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate634(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate635(.a(gate291inter12), .b(gate291inter1), .O(N769));
nor2 gate292( .a(N739), .b(N740), .O(N770) );
nor2 gate293( .a(N742), .b(N743), .O(N771) );
nor2 gate294( .a(N745), .b(N746), .O(N772) );
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );

  xor2  gate566(.a(N749), .b(N748), .O(gate296inter0));
  nand2 gate567(.a(gate296inter0), .b(s_26), .O(gate296inter1));
  and2  gate568(.a(N749), .b(N748), .O(gate296inter2));
  inv1  gate569(.a(s_26), .O(gate296inter3));
  inv1  gate570(.a(s_27), .O(gate296inter4));
  nand2 gate571(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate572(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate573(.a(N748), .O(gate296inter7));
  inv1  gate574(.a(N749), .O(gate296inter8));
  nand2 gate575(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate576(.a(s_27), .b(gate296inter3), .O(gate296inter10));
  nor2  gate577(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate578(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate579(.a(gate296inter12), .b(gate296inter1), .O(N777));
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );
nor2 gate298( .a(N751), .b(N752), .O(N781) );
nand2 gate299( .a(N756), .b(N732), .O(N782) );

  xor2  gate524(.a(N755), .b(N754), .O(gate300inter0));
  nand2 gate525(.a(gate300inter0), .b(s_20), .O(gate300inter1));
  and2  gate526(.a(N755), .b(N754), .O(gate300inter2));
  inv1  gate527(.a(s_20), .O(gate300inter3));
  inv1  gate528(.a(s_21), .O(gate300inter4));
  nand2 gate529(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate530(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate531(.a(N754), .O(gate300inter7));
  inv1  gate532(.a(N755), .O(gate300inter8));
  nand2 gate533(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate534(.a(s_21), .b(gate300inter3), .O(gate300inter10));
  nor2  gate535(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate536(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate537(.a(gate300inter12), .b(gate300inter1), .O(N785));
nor2 gate301( .a(N757), .b(N758), .O(N786) );
nor2 gate302( .a(N759), .b(N760), .O(N787) );
nor2 gate303( .a(N700), .b(N773), .O(N788) );
and2 gate304( .a(N700), .b(N773), .O(N789) );
nor2 gate305( .a(N708), .b(N778), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );
nor2 gate307( .a(N717), .b(N782), .O(N792) );
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );

  xor2  gate468(.a(N773), .b(N628), .O(gate310inter0));
  nand2 gate469(.a(gate310inter0), .b(s_12), .O(gate310inter1));
  and2  gate470(.a(N773), .b(N628), .O(gate310inter2));
  inv1  gate471(.a(s_12), .O(gate310inter3));
  inv1  gate472(.a(s_13), .O(gate310inter4));
  nand2 gate473(.a(gate310inter4), .b(gate310inter3), .O(gate310inter5));
  nor2  gate474(.a(gate310inter5), .b(gate310inter2), .O(gate310inter6));
  inv1  gate475(.a(N628), .O(gate310inter7));
  inv1  gate476(.a(N773), .O(gate310inter8));
  nand2 gate477(.a(gate310inter8), .b(gate310inter7), .O(gate310inter9));
  nand2 gate478(.a(s_13), .b(gate310inter3), .O(gate310inter10));
  nor2  gate479(.a(gate310inter10), .b(gate310inter9), .O(gate310inter11));
  nor2  gate480(.a(gate310inter11), .b(gate310inter6), .O(gate310inter12));
  nand2 gate481(.a(gate310inter12), .b(gate310inter1), .O(N795));
nand2 gate311( .a(N795), .b(N747), .O(N796) );
nor2 gate312( .a(N788), .b(N789), .O(N802) );

  xor2  gate412(.a(N791), .b(N790), .O(gate313inter0));
  nand2 gate413(.a(gate313inter0), .b(s_4), .O(gate313inter1));
  and2  gate414(.a(N791), .b(N790), .O(gate313inter2));
  inv1  gate415(.a(s_4), .O(gate313inter3));
  inv1  gate416(.a(s_5), .O(gate313inter4));
  nand2 gate417(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate418(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate419(.a(N790), .O(gate313inter7));
  inv1  gate420(.a(N791), .O(gate313inter8));
  nand2 gate421(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate422(.a(s_5), .b(gate313inter3), .O(gate313inter10));
  nor2  gate423(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate424(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate425(.a(gate313inter12), .b(gate313inter1), .O(N803));
nor2 gate314( .a(N792), .b(N793), .O(N804) );
nor2 gate315( .a(N340), .b(N794), .O(N805) );

  xor2  gate804(.a(N796), .b(N692), .O(gate316inter0));
  nand2 gate805(.a(gate316inter0), .b(s_60), .O(gate316inter1));
  and2  gate806(.a(N796), .b(N692), .O(gate316inter2));
  inv1  gate807(.a(s_60), .O(gate316inter3));
  inv1  gate808(.a(s_61), .O(gate316inter4));
  nand2 gate809(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate810(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate811(.a(N692), .O(gate316inter7));
  inv1  gate812(.a(N796), .O(gate316inter8));
  nand2 gate813(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate814(.a(s_61), .b(gate316inter3), .O(gate316inter10));
  nor2  gate815(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate816(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate817(.a(gate316inter12), .b(gate316inter1), .O(N806));
and2 gate317( .a(N692), .b(N796), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );

  xor2  gate398(.a(N796), .b(N619), .O(gate322inter0));
  nand2 gate399(.a(gate322inter0), .b(s_2), .O(gate322inter1));
  and2  gate400(.a(N796), .b(N619), .O(gate322inter2));
  inv1  gate401(.a(s_2), .O(gate322inter3));
  inv1  gate402(.a(s_3), .O(gate322inter4));
  nand2 gate403(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate404(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate405(.a(N619), .O(gate322inter7));
  inv1  gate406(.a(N796), .O(gate322inter8));
  nand2 gate407(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate408(.a(s_3), .b(gate322inter3), .O(gate322inter10));
  nor2  gate409(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate410(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate411(.a(gate322inter12), .b(gate322inter1), .O(N812));
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );
nand2 gate327( .a(N744), .b(N812), .O(N822) );
nor2 gate328( .a(N806), .b(N807), .O(N825) );
nor2 gate329( .a(N335), .b(N808), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );

  xor2  gate860(.a(N815), .b(N665), .O(gate333inter0));
  nand2 gate861(.a(gate333inter0), .b(s_68), .O(gate333inter1));
  and2  gate862(.a(N815), .b(N665), .O(gate333inter2));
  inv1  gate863(.a(s_68), .O(gate333inter3));
  inv1  gate864(.a(s_69), .O(gate333inter4));
  nand2 gate865(.a(gate333inter4), .b(gate333inter3), .O(gate333inter5));
  nor2  gate866(.a(gate333inter5), .b(gate333inter2), .O(gate333inter6));
  inv1  gate867(.a(N665), .O(gate333inter7));
  inv1  gate868(.a(N815), .O(gate333inter8));
  nand2 gate869(.a(gate333inter8), .b(gate333inter7), .O(gate333inter9));
  nand2 gate870(.a(s_69), .b(gate333inter3), .O(gate333inter10));
  nor2  gate871(.a(gate333inter10), .b(gate333inter9), .O(gate333inter11));
  nor2  gate872(.a(gate333inter11), .b(gate333inter6), .O(gate333inter12));
  nand2 gate873(.a(gate333inter12), .b(gate333inter1), .O(N830));
and2 gate334( .a(N665), .b(N815), .O(N831) );
nor2 gate335( .a(N673), .b(N819), .O(N832) );
and2 gate336( .a(N673), .b(N819), .O(N833) );
nor2 gate337( .a(N682), .b(N822), .O(N834) );
and2 gate338( .a(N682), .b(N822), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
nand2 gate344( .a(N815), .b(N593), .O(N841) );
nor2 gate345( .a(N830), .b(N831), .O(N842) );
nor2 gate346( .a(N832), .b(N833), .O(N843) );
nor2 gate347( .a(N834), .b(N835), .O(N844) );
nor2 gate348( .a(N334), .b(N836), .O(N845) );
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
and2 gate354( .a(N219), .b(N842), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );
nor2 gate362( .a(N417), .b(N851), .O(N859) );
nor2 gate363( .a(N332), .b(N852), .O(N860) );
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

endmodule