module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1975(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1976(.a(gate9inter0), .b(s_204), .O(gate9inter1));
  and2  gate1977(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1978(.a(s_204), .O(gate9inter3));
  inv1  gate1979(.a(s_205), .O(gate9inter4));
  nand2 gate1980(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1981(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1982(.a(G1), .O(gate9inter7));
  inv1  gate1983(.a(G2), .O(gate9inter8));
  nand2 gate1984(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1985(.a(s_205), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1986(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1987(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1988(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1555(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1556(.a(gate12inter0), .b(s_144), .O(gate12inter1));
  and2  gate1557(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1558(.a(s_144), .O(gate12inter3));
  inv1  gate1559(.a(s_145), .O(gate12inter4));
  nand2 gate1560(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1561(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1562(.a(G7), .O(gate12inter7));
  inv1  gate1563(.a(G8), .O(gate12inter8));
  nand2 gate1564(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1565(.a(s_145), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1566(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1567(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1568(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1933(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1934(.a(gate13inter0), .b(s_198), .O(gate13inter1));
  and2  gate1935(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1936(.a(s_198), .O(gate13inter3));
  inv1  gate1937(.a(s_199), .O(gate13inter4));
  nand2 gate1938(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1939(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1940(.a(G9), .O(gate13inter7));
  inv1  gate1941(.a(G10), .O(gate13inter8));
  nand2 gate1942(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1943(.a(s_199), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1944(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1945(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1946(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1471(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1472(.a(gate15inter0), .b(s_132), .O(gate15inter1));
  and2  gate1473(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1474(.a(s_132), .O(gate15inter3));
  inv1  gate1475(.a(s_133), .O(gate15inter4));
  nand2 gate1476(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1477(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1478(.a(G13), .O(gate15inter7));
  inv1  gate1479(.a(G14), .O(gate15inter8));
  nand2 gate1480(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1481(.a(s_133), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1482(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1483(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1484(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1331(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1332(.a(gate18inter0), .b(s_112), .O(gate18inter1));
  and2  gate1333(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1334(.a(s_112), .O(gate18inter3));
  inv1  gate1335(.a(s_113), .O(gate18inter4));
  nand2 gate1336(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1337(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1338(.a(G19), .O(gate18inter7));
  inv1  gate1339(.a(G20), .O(gate18inter8));
  nand2 gate1340(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1341(.a(s_113), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1342(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1343(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1344(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1065(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1066(.a(gate19inter0), .b(s_74), .O(gate19inter1));
  and2  gate1067(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1068(.a(s_74), .O(gate19inter3));
  inv1  gate1069(.a(s_75), .O(gate19inter4));
  nand2 gate1070(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1071(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1072(.a(G21), .O(gate19inter7));
  inv1  gate1073(.a(G22), .O(gate19inter8));
  nand2 gate1074(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1075(.a(s_75), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1076(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1077(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1078(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1989(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1990(.a(gate21inter0), .b(s_206), .O(gate21inter1));
  and2  gate1991(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1992(.a(s_206), .O(gate21inter3));
  inv1  gate1993(.a(s_207), .O(gate21inter4));
  nand2 gate1994(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1995(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1996(.a(G25), .O(gate21inter7));
  inv1  gate1997(.a(G26), .O(gate21inter8));
  nand2 gate1998(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1999(.a(s_207), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2000(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2001(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2002(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1765(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1766(.a(gate30inter0), .b(s_174), .O(gate30inter1));
  and2  gate1767(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1768(.a(s_174), .O(gate30inter3));
  inv1  gate1769(.a(s_175), .O(gate30inter4));
  nand2 gate1770(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1771(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1772(.a(G11), .O(gate30inter7));
  inv1  gate1773(.a(G15), .O(gate30inter8));
  nand2 gate1774(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1775(.a(s_175), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1776(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1777(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1778(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1177(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1178(.a(gate34inter0), .b(s_90), .O(gate34inter1));
  and2  gate1179(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1180(.a(s_90), .O(gate34inter3));
  inv1  gate1181(.a(s_91), .O(gate34inter4));
  nand2 gate1182(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1183(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1184(.a(G25), .O(gate34inter7));
  inv1  gate1185(.a(G29), .O(gate34inter8));
  nand2 gate1186(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1187(.a(s_91), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1188(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1189(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1190(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1191(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1192(.a(gate51inter0), .b(s_92), .O(gate51inter1));
  and2  gate1193(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1194(.a(s_92), .O(gate51inter3));
  inv1  gate1195(.a(s_93), .O(gate51inter4));
  nand2 gate1196(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1197(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1198(.a(G11), .O(gate51inter7));
  inv1  gate1199(.a(G281), .O(gate51inter8));
  nand2 gate1200(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1201(.a(s_93), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1202(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1203(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1204(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1905(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1906(.a(gate54inter0), .b(s_194), .O(gate54inter1));
  and2  gate1907(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1908(.a(s_194), .O(gate54inter3));
  inv1  gate1909(.a(s_195), .O(gate54inter4));
  nand2 gate1910(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1911(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1912(.a(G14), .O(gate54inter7));
  inv1  gate1913(.a(G284), .O(gate54inter8));
  nand2 gate1914(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1915(.a(s_195), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1916(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1917(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1918(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1849(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1850(.a(gate60inter0), .b(s_186), .O(gate60inter1));
  and2  gate1851(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1852(.a(s_186), .O(gate60inter3));
  inv1  gate1853(.a(s_187), .O(gate60inter4));
  nand2 gate1854(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1855(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1856(.a(G20), .O(gate60inter7));
  inv1  gate1857(.a(G293), .O(gate60inter8));
  nand2 gate1858(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1859(.a(s_187), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1860(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1861(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1862(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1639(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1640(.a(gate61inter0), .b(s_156), .O(gate61inter1));
  and2  gate1641(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1642(.a(s_156), .O(gate61inter3));
  inv1  gate1643(.a(s_157), .O(gate61inter4));
  nand2 gate1644(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1645(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1646(.a(G21), .O(gate61inter7));
  inv1  gate1647(.a(G296), .O(gate61inter8));
  nand2 gate1648(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1649(.a(s_157), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1650(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1651(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1652(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1667(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1668(.a(gate62inter0), .b(s_160), .O(gate62inter1));
  and2  gate1669(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1670(.a(s_160), .O(gate62inter3));
  inv1  gate1671(.a(s_161), .O(gate62inter4));
  nand2 gate1672(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1673(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1674(.a(G22), .O(gate62inter7));
  inv1  gate1675(.a(G296), .O(gate62inter8));
  nand2 gate1676(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1677(.a(s_161), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1678(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1679(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1680(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1485(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1486(.a(gate63inter0), .b(s_134), .O(gate63inter1));
  and2  gate1487(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1488(.a(s_134), .O(gate63inter3));
  inv1  gate1489(.a(s_135), .O(gate63inter4));
  nand2 gate1490(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1491(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1492(.a(G23), .O(gate63inter7));
  inv1  gate1493(.a(G299), .O(gate63inter8));
  nand2 gate1494(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1495(.a(s_135), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1496(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1497(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1498(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate869(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate870(.a(gate76inter0), .b(s_46), .O(gate76inter1));
  and2  gate871(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate872(.a(s_46), .O(gate76inter3));
  inv1  gate873(.a(s_47), .O(gate76inter4));
  nand2 gate874(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate875(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate876(.a(G13), .O(gate76inter7));
  inv1  gate877(.a(G317), .O(gate76inter8));
  nand2 gate878(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate879(.a(s_47), .b(gate76inter3), .O(gate76inter10));
  nor2  gate880(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate881(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate882(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1961(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1962(.a(gate78inter0), .b(s_202), .O(gate78inter1));
  and2  gate1963(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1964(.a(s_202), .O(gate78inter3));
  inv1  gate1965(.a(s_203), .O(gate78inter4));
  nand2 gate1966(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1967(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1968(.a(G6), .O(gate78inter7));
  inv1  gate1969(.a(G320), .O(gate78inter8));
  nand2 gate1970(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1971(.a(s_203), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1972(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1973(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1974(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate729(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate730(.a(gate79inter0), .b(s_26), .O(gate79inter1));
  and2  gate731(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate732(.a(s_26), .O(gate79inter3));
  inv1  gate733(.a(s_27), .O(gate79inter4));
  nand2 gate734(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate735(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate736(.a(G10), .O(gate79inter7));
  inv1  gate737(.a(G323), .O(gate79inter8));
  nand2 gate738(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate739(.a(s_27), .b(gate79inter3), .O(gate79inter10));
  nor2  gate740(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate741(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate742(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1681(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1682(.a(gate80inter0), .b(s_162), .O(gate80inter1));
  and2  gate1683(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1684(.a(s_162), .O(gate80inter3));
  inv1  gate1685(.a(s_163), .O(gate80inter4));
  nand2 gate1686(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1687(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1688(.a(G14), .O(gate80inter7));
  inv1  gate1689(.a(G323), .O(gate80inter8));
  nand2 gate1690(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1691(.a(s_163), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1692(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1693(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1694(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate925(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate926(.a(gate86inter0), .b(s_54), .O(gate86inter1));
  and2  gate927(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate928(.a(s_54), .O(gate86inter3));
  inv1  gate929(.a(s_55), .O(gate86inter4));
  nand2 gate930(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate931(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate932(.a(G8), .O(gate86inter7));
  inv1  gate933(.a(G332), .O(gate86inter8));
  nand2 gate934(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate935(.a(s_55), .b(gate86inter3), .O(gate86inter10));
  nor2  gate936(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate937(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate938(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate701(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate702(.a(gate97inter0), .b(s_22), .O(gate97inter1));
  and2  gate703(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate704(.a(s_22), .O(gate97inter3));
  inv1  gate705(.a(s_23), .O(gate97inter4));
  nand2 gate706(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate707(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate708(.a(G19), .O(gate97inter7));
  inv1  gate709(.a(G350), .O(gate97inter8));
  nand2 gate710(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate711(.a(s_23), .b(gate97inter3), .O(gate97inter10));
  nor2  gate712(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate713(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate714(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate813(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate814(.a(gate98inter0), .b(s_38), .O(gate98inter1));
  and2  gate815(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate816(.a(s_38), .O(gate98inter3));
  inv1  gate817(.a(s_39), .O(gate98inter4));
  nand2 gate818(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate819(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate820(.a(G23), .O(gate98inter7));
  inv1  gate821(.a(G350), .O(gate98inter8));
  nand2 gate822(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate823(.a(s_39), .b(gate98inter3), .O(gate98inter10));
  nor2  gate824(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate825(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate826(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1821(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1822(.a(gate100inter0), .b(s_182), .O(gate100inter1));
  and2  gate1823(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1824(.a(s_182), .O(gate100inter3));
  inv1  gate1825(.a(s_183), .O(gate100inter4));
  nand2 gate1826(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1827(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1828(.a(G31), .O(gate100inter7));
  inv1  gate1829(.a(G353), .O(gate100inter8));
  nand2 gate1830(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1831(.a(s_183), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1832(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1833(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1834(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1611(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1612(.a(gate101inter0), .b(s_152), .O(gate101inter1));
  and2  gate1613(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1614(.a(s_152), .O(gate101inter3));
  inv1  gate1615(.a(s_153), .O(gate101inter4));
  nand2 gate1616(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1617(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1618(.a(G20), .O(gate101inter7));
  inv1  gate1619(.a(G356), .O(gate101inter8));
  nand2 gate1620(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1621(.a(s_153), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1622(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1623(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1624(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1051(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1052(.a(gate103inter0), .b(s_72), .O(gate103inter1));
  and2  gate1053(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1054(.a(s_72), .O(gate103inter3));
  inv1  gate1055(.a(s_73), .O(gate103inter4));
  nand2 gate1056(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1057(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1058(.a(G28), .O(gate103inter7));
  inv1  gate1059(.a(G359), .O(gate103inter8));
  nand2 gate1060(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1061(.a(s_73), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1062(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1063(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1064(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1345(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1346(.a(gate104inter0), .b(s_114), .O(gate104inter1));
  and2  gate1347(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1348(.a(s_114), .O(gate104inter3));
  inv1  gate1349(.a(s_115), .O(gate104inter4));
  nand2 gate1350(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1351(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1352(.a(G32), .O(gate104inter7));
  inv1  gate1353(.a(G359), .O(gate104inter8));
  nand2 gate1354(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1355(.a(s_115), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1356(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1357(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1358(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1695(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1696(.a(gate105inter0), .b(s_164), .O(gate105inter1));
  and2  gate1697(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1698(.a(s_164), .O(gate105inter3));
  inv1  gate1699(.a(s_165), .O(gate105inter4));
  nand2 gate1700(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1701(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1702(.a(G362), .O(gate105inter7));
  inv1  gate1703(.a(G363), .O(gate105inter8));
  nand2 gate1704(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1705(.a(s_165), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1706(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1707(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1708(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1093(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1094(.a(gate107inter0), .b(s_78), .O(gate107inter1));
  and2  gate1095(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1096(.a(s_78), .O(gate107inter3));
  inv1  gate1097(.a(s_79), .O(gate107inter4));
  nand2 gate1098(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1099(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1100(.a(G366), .O(gate107inter7));
  inv1  gate1101(.a(G367), .O(gate107inter8));
  nand2 gate1102(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1103(.a(s_79), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1104(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1105(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1106(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1289(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1290(.a(gate116inter0), .b(s_106), .O(gate116inter1));
  and2  gate1291(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1292(.a(s_106), .O(gate116inter3));
  inv1  gate1293(.a(s_107), .O(gate116inter4));
  nand2 gate1294(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1295(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1296(.a(G384), .O(gate116inter7));
  inv1  gate1297(.a(G385), .O(gate116inter8));
  nand2 gate1298(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1299(.a(s_107), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1300(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1301(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1302(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate659(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate660(.a(gate117inter0), .b(s_16), .O(gate117inter1));
  and2  gate661(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate662(.a(s_16), .O(gate117inter3));
  inv1  gate663(.a(s_17), .O(gate117inter4));
  nand2 gate664(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate665(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate666(.a(G386), .O(gate117inter7));
  inv1  gate667(.a(G387), .O(gate117inter8));
  nand2 gate668(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate669(.a(s_17), .b(gate117inter3), .O(gate117inter10));
  nor2  gate670(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate671(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate672(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1023(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1024(.a(gate121inter0), .b(s_68), .O(gate121inter1));
  and2  gate1025(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1026(.a(s_68), .O(gate121inter3));
  inv1  gate1027(.a(s_69), .O(gate121inter4));
  nand2 gate1028(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1029(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1030(.a(G394), .O(gate121inter7));
  inv1  gate1031(.a(G395), .O(gate121inter8));
  nand2 gate1032(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1033(.a(s_69), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1034(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1035(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1036(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2073(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2074(.a(gate123inter0), .b(s_218), .O(gate123inter1));
  and2  gate2075(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2076(.a(s_218), .O(gate123inter3));
  inv1  gate2077(.a(s_219), .O(gate123inter4));
  nand2 gate2078(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2079(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2080(.a(G398), .O(gate123inter7));
  inv1  gate2081(.a(G399), .O(gate123inter8));
  nand2 gate2082(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2083(.a(s_219), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2084(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2085(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2086(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1247(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1248(.a(gate124inter0), .b(s_100), .O(gate124inter1));
  and2  gate1249(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1250(.a(s_100), .O(gate124inter3));
  inv1  gate1251(.a(s_101), .O(gate124inter4));
  nand2 gate1252(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1253(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1254(.a(G400), .O(gate124inter7));
  inv1  gate1255(.a(G401), .O(gate124inter8));
  nand2 gate1256(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1257(.a(s_101), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1258(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1259(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1260(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate589(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate590(.a(gate127inter0), .b(s_6), .O(gate127inter1));
  and2  gate591(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate592(.a(s_6), .O(gate127inter3));
  inv1  gate593(.a(s_7), .O(gate127inter4));
  nand2 gate594(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate595(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate596(.a(G406), .O(gate127inter7));
  inv1  gate597(.a(G407), .O(gate127inter8));
  nand2 gate598(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate599(.a(s_7), .b(gate127inter3), .O(gate127inter10));
  nor2  gate600(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate601(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate602(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1205(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1206(.a(gate134inter0), .b(s_94), .O(gate134inter1));
  and2  gate1207(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1208(.a(s_94), .O(gate134inter3));
  inv1  gate1209(.a(s_95), .O(gate134inter4));
  nand2 gate1210(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1211(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1212(.a(G420), .O(gate134inter7));
  inv1  gate1213(.a(G421), .O(gate134inter8));
  nand2 gate1214(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1215(.a(s_95), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1216(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1217(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1218(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1835(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1836(.a(gate138inter0), .b(s_184), .O(gate138inter1));
  and2  gate1837(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1838(.a(s_184), .O(gate138inter3));
  inv1  gate1839(.a(s_185), .O(gate138inter4));
  nand2 gate1840(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1841(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1842(.a(G432), .O(gate138inter7));
  inv1  gate1843(.a(G435), .O(gate138inter8));
  nand2 gate1844(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1845(.a(s_185), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1846(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1847(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1848(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate757(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate758(.a(gate139inter0), .b(s_30), .O(gate139inter1));
  and2  gate759(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate760(.a(s_30), .O(gate139inter3));
  inv1  gate761(.a(s_31), .O(gate139inter4));
  nand2 gate762(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate763(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate764(.a(G438), .O(gate139inter7));
  inv1  gate765(.a(G441), .O(gate139inter8));
  nand2 gate766(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate767(.a(s_31), .b(gate139inter3), .O(gate139inter10));
  nor2  gate768(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate769(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate770(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1303(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1304(.a(gate145inter0), .b(s_108), .O(gate145inter1));
  and2  gate1305(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1306(.a(s_108), .O(gate145inter3));
  inv1  gate1307(.a(s_109), .O(gate145inter4));
  nand2 gate1308(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1309(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1310(.a(G474), .O(gate145inter7));
  inv1  gate1311(.a(G477), .O(gate145inter8));
  nand2 gate1312(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1313(.a(s_109), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1314(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1315(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1316(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate645(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate646(.a(gate146inter0), .b(s_14), .O(gate146inter1));
  and2  gate647(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate648(.a(s_14), .O(gate146inter3));
  inv1  gate649(.a(s_15), .O(gate146inter4));
  nand2 gate650(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate651(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate652(.a(G480), .O(gate146inter7));
  inv1  gate653(.a(G483), .O(gate146inter8));
  nand2 gate654(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate655(.a(s_15), .b(gate146inter3), .O(gate146inter10));
  nor2  gate656(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate657(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate658(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1597(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1598(.a(gate150inter0), .b(s_150), .O(gate150inter1));
  and2  gate1599(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1600(.a(s_150), .O(gate150inter3));
  inv1  gate1601(.a(s_151), .O(gate150inter4));
  nand2 gate1602(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1603(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1604(.a(G504), .O(gate150inter7));
  inv1  gate1605(.a(G507), .O(gate150inter8));
  nand2 gate1606(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1607(.a(s_151), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1608(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1609(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1610(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1457(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1458(.a(gate151inter0), .b(s_130), .O(gate151inter1));
  and2  gate1459(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1460(.a(s_130), .O(gate151inter3));
  inv1  gate1461(.a(s_131), .O(gate151inter4));
  nand2 gate1462(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1463(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1464(.a(G510), .O(gate151inter7));
  inv1  gate1465(.a(G513), .O(gate151inter8));
  nand2 gate1466(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1467(.a(s_131), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1468(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1469(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1470(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate743(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate744(.a(gate155inter0), .b(s_28), .O(gate155inter1));
  and2  gate745(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate746(.a(s_28), .O(gate155inter3));
  inv1  gate747(.a(s_29), .O(gate155inter4));
  nand2 gate748(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate749(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate750(.a(G432), .O(gate155inter7));
  inv1  gate751(.a(G525), .O(gate155inter8));
  nand2 gate752(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate753(.a(s_29), .b(gate155inter3), .O(gate155inter10));
  nor2  gate754(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate755(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate756(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1751(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1752(.a(gate156inter0), .b(s_172), .O(gate156inter1));
  and2  gate1753(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1754(.a(s_172), .O(gate156inter3));
  inv1  gate1755(.a(s_173), .O(gate156inter4));
  nand2 gate1756(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1757(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1758(.a(G435), .O(gate156inter7));
  inv1  gate1759(.a(G525), .O(gate156inter8));
  nand2 gate1760(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1761(.a(s_173), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1762(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1763(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1764(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1527(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1528(.a(gate158inter0), .b(s_140), .O(gate158inter1));
  and2  gate1529(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1530(.a(s_140), .O(gate158inter3));
  inv1  gate1531(.a(s_141), .O(gate158inter4));
  nand2 gate1532(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1533(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1534(.a(G441), .O(gate158inter7));
  inv1  gate1535(.a(G528), .O(gate158inter8));
  nand2 gate1536(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1537(.a(s_141), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1538(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1539(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1540(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate981(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate982(.a(gate160inter0), .b(s_62), .O(gate160inter1));
  and2  gate983(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate984(.a(s_62), .O(gate160inter3));
  inv1  gate985(.a(s_63), .O(gate160inter4));
  nand2 gate986(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate987(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate988(.a(G447), .O(gate160inter7));
  inv1  gate989(.a(G531), .O(gate160inter8));
  nand2 gate990(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate991(.a(s_63), .b(gate160inter3), .O(gate160inter10));
  nor2  gate992(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate993(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate994(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1947(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1948(.a(gate161inter0), .b(s_200), .O(gate161inter1));
  and2  gate1949(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1950(.a(s_200), .O(gate161inter3));
  inv1  gate1951(.a(s_201), .O(gate161inter4));
  nand2 gate1952(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1953(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1954(.a(G450), .O(gate161inter7));
  inv1  gate1955(.a(G534), .O(gate161inter8));
  nand2 gate1956(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1957(.a(s_201), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1958(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1959(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1960(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate603(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate604(.a(gate163inter0), .b(s_8), .O(gate163inter1));
  and2  gate605(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate606(.a(s_8), .O(gate163inter3));
  inv1  gate607(.a(s_9), .O(gate163inter4));
  nand2 gate608(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate609(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate610(.a(G456), .O(gate163inter7));
  inv1  gate611(.a(G537), .O(gate163inter8));
  nand2 gate612(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate613(.a(s_9), .b(gate163inter3), .O(gate163inter10));
  nor2  gate614(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate615(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate616(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1709(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1710(.a(gate172inter0), .b(s_166), .O(gate172inter1));
  and2  gate1711(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1712(.a(s_166), .O(gate172inter3));
  inv1  gate1713(.a(s_167), .O(gate172inter4));
  nand2 gate1714(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1715(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1716(.a(G483), .O(gate172inter7));
  inv1  gate1717(.a(G549), .O(gate172inter8));
  nand2 gate1718(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1719(.a(s_167), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1720(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1721(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1722(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate967(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate968(.a(gate181inter0), .b(s_60), .O(gate181inter1));
  and2  gate969(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate970(.a(s_60), .O(gate181inter3));
  inv1  gate971(.a(s_61), .O(gate181inter4));
  nand2 gate972(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate973(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate974(.a(G510), .O(gate181inter7));
  inv1  gate975(.a(G564), .O(gate181inter8));
  nand2 gate976(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate977(.a(s_61), .b(gate181inter3), .O(gate181inter10));
  nor2  gate978(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate979(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate980(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1429(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1430(.a(gate182inter0), .b(s_126), .O(gate182inter1));
  and2  gate1431(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1432(.a(s_126), .O(gate182inter3));
  inv1  gate1433(.a(s_127), .O(gate182inter4));
  nand2 gate1434(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1435(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1436(.a(G513), .O(gate182inter7));
  inv1  gate1437(.a(G564), .O(gate182inter8));
  nand2 gate1438(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1439(.a(s_127), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1440(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1441(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1442(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate2101(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2102(.a(gate183inter0), .b(s_222), .O(gate183inter1));
  and2  gate2103(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2104(.a(s_222), .O(gate183inter3));
  inv1  gate2105(.a(s_223), .O(gate183inter4));
  nand2 gate2106(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2107(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2108(.a(G516), .O(gate183inter7));
  inv1  gate2109(.a(G567), .O(gate183inter8));
  nand2 gate2110(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2111(.a(s_223), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2112(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2113(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2114(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1723(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1724(.a(gate187inter0), .b(s_168), .O(gate187inter1));
  and2  gate1725(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1726(.a(s_168), .O(gate187inter3));
  inv1  gate1727(.a(s_169), .O(gate187inter4));
  nand2 gate1728(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1729(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1730(.a(G574), .O(gate187inter7));
  inv1  gate1731(.a(G575), .O(gate187inter8));
  nand2 gate1732(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1733(.a(s_169), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1734(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1735(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1736(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate953(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate954(.a(gate190inter0), .b(s_58), .O(gate190inter1));
  and2  gate955(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate956(.a(s_58), .O(gate190inter3));
  inv1  gate957(.a(s_59), .O(gate190inter4));
  nand2 gate958(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate959(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate960(.a(G580), .O(gate190inter7));
  inv1  gate961(.a(G581), .O(gate190inter8));
  nand2 gate962(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate963(.a(s_59), .b(gate190inter3), .O(gate190inter10));
  nor2  gate964(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate965(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate966(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate883(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate884(.a(gate191inter0), .b(s_48), .O(gate191inter1));
  and2  gate885(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate886(.a(s_48), .O(gate191inter3));
  inv1  gate887(.a(s_49), .O(gate191inter4));
  nand2 gate888(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate889(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate890(.a(G582), .O(gate191inter7));
  inv1  gate891(.a(G583), .O(gate191inter8));
  nand2 gate892(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate893(.a(s_49), .b(gate191inter3), .O(gate191inter10));
  nor2  gate894(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate895(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate896(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2045(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2046(.a(gate194inter0), .b(s_214), .O(gate194inter1));
  and2  gate2047(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2048(.a(s_214), .O(gate194inter3));
  inv1  gate2049(.a(s_215), .O(gate194inter4));
  nand2 gate2050(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2051(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2052(.a(G588), .O(gate194inter7));
  inv1  gate2053(.a(G589), .O(gate194inter8));
  nand2 gate2054(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2055(.a(s_215), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2056(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2057(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2058(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate2087(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2088(.a(gate196inter0), .b(s_220), .O(gate196inter1));
  and2  gate2089(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2090(.a(s_220), .O(gate196inter3));
  inv1  gate2091(.a(s_221), .O(gate196inter4));
  nand2 gate2092(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2093(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2094(.a(G592), .O(gate196inter7));
  inv1  gate2095(.a(G593), .O(gate196inter8));
  nand2 gate2096(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2097(.a(s_221), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2098(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2099(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2100(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1737(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1738(.a(gate200inter0), .b(s_170), .O(gate200inter1));
  and2  gate1739(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1740(.a(s_170), .O(gate200inter3));
  inv1  gate1741(.a(s_171), .O(gate200inter4));
  nand2 gate1742(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1743(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1744(.a(G600), .O(gate200inter7));
  inv1  gate1745(.a(G601), .O(gate200inter8));
  nand2 gate1746(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1747(.a(s_171), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1748(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1749(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1750(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1653(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1654(.a(gate201inter0), .b(s_158), .O(gate201inter1));
  and2  gate1655(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1656(.a(s_158), .O(gate201inter3));
  inv1  gate1657(.a(s_159), .O(gate201inter4));
  nand2 gate1658(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1659(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1660(.a(G602), .O(gate201inter7));
  inv1  gate1661(.a(G607), .O(gate201inter8));
  nand2 gate1662(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1663(.a(s_159), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1664(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1665(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1666(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1121(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1122(.a(gate203inter0), .b(s_82), .O(gate203inter1));
  and2  gate1123(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1124(.a(s_82), .O(gate203inter3));
  inv1  gate1125(.a(s_83), .O(gate203inter4));
  nand2 gate1126(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1127(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1128(.a(G602), .O(gate203inter7));
  inv1  gate1129(.a(G612), .O(gate203inter8));
  nand2 gate1130(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1131(.a(s_83), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1132(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1133(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1134(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1891(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1892(.a(gate209inter0), .b(s_192), .O(gate209inter1));
  and2  gate1893(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1894(.a(s_192), .O(gate209inter3));
  inv1  gate1895(.a(s_193), .O(gate209inter4));
  nand2 gate1896(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1897(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1898(.a(G602), .O(gate209inter7));
  inv1  gate1899(.a(G666), .O(gate209inter8));
  nand2 gate1900(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1901(.a(s_193), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1902(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1903(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1904(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1793(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1794(.a(gate213inter0), .b(s_178), .O(gate213inter1));
  and2  gate1795(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1796(.a(s_178), .O(gate213inter3));
  inv1  gate1797(.a(s_179), .O(gate213inter4));
  nand2 gate1798(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1799(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1800(.a(G602), .O(gate213inter7));
  inv1  gate1801(.a(G672), .O(gate213inter8));
  nand2 gate1802(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1803(.a(s_179), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1804(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1805(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1806(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1779(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1780(.a(gate221inter0), .b(s_176), .O(gate221inter1));
  and2  gate1781(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1782(.a(s_176), .O(gate221inter3));
  inv1  gate1783(.a(s_177), .O(gate221inter4));
  nand2 gate1784(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1785(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1786(.a(G622), .O(gate221inter7));
  inv1  gate1787(.a(G684), .O(gate221inter8));
  nand2 gate1788(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1789(.a(s_177), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1790(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1791(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1792(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate897(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate898(.a(gate226inter0), .b(s_50), .O(gate226inter1));
  and2  gate899(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate900(.a(s_50), .O(gate226inter3));
  inv1  gate901(.a(s_51), .O(gate226inter4));
  nand2 gate902(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate903(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate904(.a(G692), .O(gate226inter7));
  inv1  gate905(.a(G693), .O(gate226inter8));
  nand2 gate906(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate907(.a(s_51), .b(gate226inter3), .O(gate226inter10));
  nor2  gate908(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate909(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate910(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2017(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2018(.a(gate228inter0), .b(s_210), .O(gate228inter1));
  and2  gate2019(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2020(.a(s_210), .O(gate228inter3));
  inv1  gate2021(.a(s_211), .O(gate228inter4));
  nand2 gate2022(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2023(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2024(.a(G696), .O(gate228inter7));
  inv1  gate2025(.a(G697), .O(gate228inter8));
  nand2 gate2026(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2027(.a(s_211), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2028(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2029(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2030(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate911(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate912(.a(gate231inter0), .b(s_52), .O(gate231inter1));
  and2  gate913(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate914(.a(s_52), .O(gate231inter3));
  inv1  gate915(.a(s_53), .O(gate231inter4));
  nand2 gate916(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate917(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate918(.a(G702), .O(gate231inter7));
  inv1  gate919(.a(G703), .O(gate231inter8));
  nand2 gate920(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate921(.a(s_53), .b(gate231inter3), .O(gate231inter10));
  nor2  gate922(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate923(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate924(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1359(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1360(.a(gate234inter0), .b(s_116), .O(gate234inter1));
  and2  gate1361(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1362(.a(s_116), .O(gate234inter3));
  inv1  gate1363(.a(s_117), .O(gate234inter4));
  nand2 gate1364(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1365(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1366(.a(G245), .O(gate234inter7));
  inv1  gate1367(.a(G721), .O(gate234inter8));
  nand2 gate1368(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1369(.a(s_117), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1370(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1371(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1372(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1863(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1864(.a(gate242inter0), .b(s_188), .O(gate242inter1));
  and2  gate1865(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1866(.a(s_188), .O(gate242inter3));
  inv1  gate1867(.a(s_189), .O(gate242inter4));
  nand2 gate1868(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1869(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1870(.a(G718), .O(gate242inter7));
  inv1  gate1871(.a(G730), .O(gate242inter8));
  nand2 gate1872(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1873(.a(s_189), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1874(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1875(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1876(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate575(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate576(.a(gate246inter0), .b(s_4), .O(gate246inter1));
  and2  gate577(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate578(.a(s_4), .O(gate246inter3));
  inv1  gate579(.a(s_5), .O(gate246inter4));
  nand2 gate580(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate581(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate582(.a(G724), .O(gate246inter7));
  inv1  gate583(.a(G736), .O(gate246inter8));
  nand2 gate584(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate585(.a(s_5), .b(gate246inter3), .O(gate246inter10));
  nor2  gate586(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate587(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate588(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1919(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1920(.a(gate248inter0), .b(s_196), .O(gate248inter1));
  and2  gate1921(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1922(.a(s_196), .O(gate248inter3));
  inv1  gate1923(.a(s_197), .O(gate248inter4));
  nand2 gate1924(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1925(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1926(.a(G727), .O(gate248inter7));
  inv1  gate1927(.a(G739), .O(gate248inter8));
  nand2 gate1928(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1929(.a(s_197), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1930(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1931(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1932(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1219(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1220(.a(gate249inter0), .b(s_96), .O(gate249inter1));
  and2  gate1221(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1222(.a(s_96), .O(gate249inter3));
  inv1  gate1223(.a(s_97), .O(gate249inter4));
  nand2 gate1224(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1225(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1226(.a(G254), .O(gate249inter7));
  inv1  gate1227(.a(G742), .O(gate249inter8));
  nand2 gate1228(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1229(.a(s_97), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1230(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1231(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1232(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1625(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1626(.a(gate252inter0), .b(s_154), .O(gate252inter1));
  and2  gate1627(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1628(.a(s_154), .O(gate252inter3));
  inv1  gate1629(.a(s_155), .O(gate252inter4));
  nand2 gate1630(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1631(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1632(.a(G709), .O(gate252inter7));
  inv1  gate1633(.a(G745), .O(gate252inter8));
  nand2 gate1634(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1635(.a(s_155), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1636(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1637(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1638(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1373(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1374(.a(gate254inter0), .b(s_118), .O(gate254inter1));
  and2  gate1375(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1376(.a(s_118), .O(gate254inter3));
  inv1  gate1377(.a(s_119), .O(gate254inter4));
  nand2 gate1378(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1379(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1380(.a(G712), .O(gate254inter7));
  inv1  gate1381(.a(G748), .O(gate254inter8));
  nand2 gate1382(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1383(.a(s_119), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1384(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1385(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1386(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1261(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1262(.a(gate258inter0), .b(s_102), .O(gate258inter1));
  and2  gate1263(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1264(.a(s_102), .O(gate258inter3));
  inv1  gate1265(.a(s_103), .O(gate258inter4));
  nand2 gate1266(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1267(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1268(.a(G756), .O(gate258inter7));
  inv1  gate1269(.a(G757), .O(gate258inter8));
  nand2 gate1270(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1271(.a(s_103), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1272(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1273(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1274(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2059(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2060(.a(gate263inter0), .b(s_216), .O(gate263inter1));
  and2  gate2061(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2062(.a(s_216), .O(gate263inter3));
  inv1  gate2063(.a(s_217), .O(gate263inter4));
  nand2 gate2064(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2065(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2066(.a(G766), .O(gate263inter7));
  inv1  gate2067(.a(G767), .O(gate263inter8));
  nand2 gate2068(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2069(.a(s_217), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2070(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2071(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2072(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1037(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1038(.a(gate271inter0), .b(s_70), .O(gate271inter1));
  and2  gate1039(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1040(.a(s_70), .O(gate271inter3));
  inv1  gate1041(.a(s_71), .O(gate271inter4));
  nand2 gate1042(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1043(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1044(.a(G660), .O(gate271inter7));
  inv1  gate1045(.a(G788), .O(gate271inter8));
  nand2 gate1046(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1047(.a(s_71), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1048(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1049(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1050(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate827(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate828(.a(gate274inter0), .b(s_40), .O(gate274inter1));
  and2  gate829(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate830(.a(s_40), .O(gate274inter3));
  inv1  gate831(.a(s_41), .O(gate274inter4));
  nand2 gate832(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate833(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate834(.a(G770), .O(gate274inter7));
  inv1  gate835(.a(G794), .O(gate274inter8));
  nand2 gate836(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate837(.a(s_41), .b(gate274inter3), .O(gate274inter10));
  nor2  gate838(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate839(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate840(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate995(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate996(.a(gate286inter0), .b(s_64), .O(gate286inter1));
  and2  gate997(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate998(.a(s_64), .O(gate286inter3));
  inv1  gate999(.a(s_65), .O(gate286inter4));
  nand2 gate1000(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1001(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1002(.a(G788), .O(gate286inter7));
  inv1  gate1003(.a(G812), .O(gate286inter8));
  nand2 gate1004(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1005(.a(s_65), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1006(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1007(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1008(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2129(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2130(.a(gate288inter0), .b(s_226), .O(gate288inter1));
  and2  gate2131(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2132(.a(s_226), .O(gate288inter3));
  inv1  gate2133(.a(s_227), .O(gate288inter4));
  nand2 gate2134(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2135(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2136(.a(G791), .O(gate288inter7));
  inv1  gate2137(.a(G815), .O(gate288inter8));
  nand2 gate2138(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2139(.a(s_227), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2140(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2141(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2142(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate855(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate856(.a(gate289inter0), .b(s_44), .O(gate289inter1));
  and2  gate857(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate858(.a(s_44), .O(gate289inter3));
  inv1  gate859(.a(s_45), .O(gate289inter4));
  nand2 gate860(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate861(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate862(.a(G818), .O(gate289inter7));
  inv1  gate863(.a(G819), .O(gate289inter8));
  nand2 gate864(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate865(.a(s_45), .b(gate289inter3), .O(gate289inter10));
  nor2  gate866(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate867(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate868(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate939(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate940(.a(gate292inter0), .b(s_56), .O(gate292inter1));
  and2  gate941(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate942(.a(s_56), .O(gate292inter3));
  inv1  gate943(.a(s_57), .O(gate292inter4));
  nand2 gate944(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate945(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate946(.a(G824), .O(gate292inter7));
  inv1  gate947(.a(G825), .O(gate292inter8));
  nand2 gate948(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate949(.a(s_57), .b(gate292inter3), .O(gate292inter10));
  nor2  gate950(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate951(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate952(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate561(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate562(.a(gate293inter0), .b(s_2), .O(gate293inter1));
  and2  gate563(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate564(.a(s_2), .O(gate293inter3));
  inv1  gate565(.a(s_3), .O(gate293inter4));
  nand2 gate566(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate567(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate568(.a(G828), .O(gate293inter7));
  inv1  gate569(.a(G829), .O(gate293inter8));
  nand2 gate570(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate571(.a(s_3), .b(gate293inter3), .O(gate293inter10));
  nor2  gate572(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate573(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate574(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate687(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate688(.a(gate295inter0), .b(s_20), .O(gate295inter1));
  and2  gate689(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate690(.a(s_20), .O(gate295inter3));
  inv1  gate691(.a(s_21), .O(gate295inter4));
  nand2 gate692(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate693(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate694(.a(G830), .O(gate295inter7));
  inv1  gate695(.a(G831), .O(gate295inter8));
  nand2 gate696(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate697(.a(s_21), .b(gate295inter3), .O(gate295inter10));
  nor2  gate698(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate699(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate700(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate547(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate548(.a(gate296inter0), .b(s_0), .O(gate296inter1));
  and2  gate549(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate550(.a(s_0), .O(gate296inter3));
  inv1  gate551(.a(s_1), .O(gate296inter4));
  nand2 gate552(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate553(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate554(.a(G826), .O(gate296inter7));
  inv1  gate555(.a(G827), .O(gate296inter8));
  nand2 gate556(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate557(.a(s_1), .b(gate296inter3), .O(gate296inter10));
  nor2  gate558(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate559(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate560(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2003(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2004(.a(gate389inter0), .b(s_208), .O(gate389inter1));
  and2  gate2005(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2006(.a(s_208), .O(gate389inter3));
  inv1  gate2007(.a(s_209), .O(gate389inter4));
  nand2 gate2008(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2009(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2010(.a(G3), .O(gate389inter7));
  inv1  gate2011(.a(G1042), .O(gate389inter8));
  nand2 gate2012(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2013(.a(s_209), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2014(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2015(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2016(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate715(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate716(.a(gate390inter0), .b(s_24), .O(gate390inter1));
  and2  gate717(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate718(.a(s_24), .O(gate390inter3));
  inv1  gate719(.a(s_25), .O(gate390inter4));
  nand2 gate720(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate721(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate722(.a(G4), .O(gate390inter7));
  inv1  gate723(.a(G1045), .O(gate390inter8));
  nand2 gate724(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate725(.a(s_25), .b(gate390inter3), .O(gate390inter10));
  nor2  gate726(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate727(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate728(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1163(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1164(.a(gate391inter0), .b(s_88), .O(gate391inter1));
  and2  gate1165(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1166(.a(s_88), .O(gate391inter3));
  inv1  gate1167(.a(s_89), .O(gate391inter4));
  nand2 gate1168(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1169(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1170(.a(G5), .O(gate391inter7));
  inv1  gate1171(.a(G1048), .O(gate391inter8));
  nand2 gate1172(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1173(.a(s_89), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1174(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1175(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1176(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1443(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1444(.a(gate393inter0), .b(s_128), .O(gate393inter1));
  and2  gate1445(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1446(.a(s_128), .O(gate393inter3));
  inv1  gate1447(.a(s_129), .O(gate393inter4));
  nand2 gate1448(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1449(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1450(.a(G7), .O(gate393inter7));
  inv1  gate1451(.a(G1054), .O(gate393inter8));
  nand2 gate1452(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1453(.a(s_129), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1454(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1455(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1456(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1877(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1878(.a(gate395inter0), .b(s_190), .O(gate395inter1));
  and2  gate1879(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1880(.a(s_190), .O(gate395inter3));
  inv1  gate1881(.a(s_191), .O(gate395inter4));
  nand2 gate1882(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1883(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1884(.a(G9), .O(gate395inter7));
  inv1  gate1885(.a(G1060), .O(gate395inter8));
  nand2 gate1886(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1887(.a(s_191), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1888(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1889(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1890(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate785(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate786(.a(gate398inter0), .b(s_34), .O(gate398inter1));
  and2  gate787(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate788(.a(s_34), .O(gate398inter3));
  inv1  gate789(.a(s_35), .O(gate398inter4));
  nand2 gate790(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate791(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate792(.a(G12), .O(gate398inter7));
  inv1  gate793(.a(G1069), .O(gate398inter8));
  nand2 gate794(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate795(.a(s_35), .b(gate398inter3), .O(gate398inter10));
  nor2  gate796(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate797(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate798(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1317(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1318(.a(gate401inter0), .b(s_110), .O(gate401inter1));
  and2  gate1319(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1320(.a(s_110), .O(gate401inter3));
  inv1  gate1321(.a(s_111), .O(gate401inter4));
  nand2 gate1322(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1323(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1324(.a(G15), .O(gate401inter7));
  inv1  gate1325(.a(G1078), .O(gate401inter8));
  nand2 gate1326(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1327(.a(s_111), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1328(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1329(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1330(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate841(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate842(.a(gate409inter0), .b(s_42), .O(gate409inter1));
  and2  gate843(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate844(.a(s_42), .O(gate409inter3));
  inv1  gate845(.a(s_43), .O(gate409inter4));
  nand2 gate846(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate847(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate848(.a(G23), .O(gate409inter7));
  inv1  gate849(.a(G1102), .O(gate409inter8));
  nand2 gate850(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate851(.a(s_43), .b(gate409inter3), .O(gate409inter10));
  nor2  gate852(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate853(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate854(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2143(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2144(.a(gate410inter0), .b(s_228), .O(gate410inter1));
  and2  gate2145(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2146(.a(s_228), .O(gate410inter3));
  inv1  gate2147(.a(s_229), .O(gate410inter4));
  nand2 gate2148(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2149(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2150(.a(G24), .O(gate410inter7));
  inv1  gate2151(.a(G1105), .O(gate410inter8));
  nand2 gate2152(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2153(.a(s_229), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2154(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2155(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2156(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1569(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1570(.a(gate413inter0), .b(s_146), .O(gate413inter1));
  and2  gate1571(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1572(.a(s_146), .O(gate413inter3));
  inv1  gate1573(.a(s_147), .O(gate413inter4));
  nand2 gate1574(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1575(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1576(.a(G27), .O(gate413inter7));
  inv1  gate1577(.a(G1114), .O(gate413inter8));
  nand2 gate1578(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1579(.a(s_147), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1580(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1581(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1582(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1275(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1276(.a(gate416inter0), .b(s_104), .O(gate416inter1));
  and2  gate1277(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1278(.a(s_104), .O(gate416inter3));
  inv1  gate1279(.a(s_105), .O(gate416inter4));
  nand2 gate1280(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1281(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1282(.a(G30), .O(gate416inter7));
  inv1  gate1283(.a(G1123), .O(gate416inter8));
  nand2 gate1284(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1285(.a(s_105), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1286(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1287(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1288(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1513(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1514(.a(gate420inter0), .b(s_138), .O(gate420inter1));
  and2  gate1515(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1516(.a(s_138), .O(gate420inter3));
  inv1  gate1517(.a(s_139), .O(gate420inter4));
  nand2 gate1518(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1519(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1520(.a(G1036), .O(gate420inter7));
  inv1  gate1521(.a(G1132), .O(gate420inter8));
  nand2 gate1522(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1523(.a(s_139), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1524(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1525(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1526(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2115(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2116(.a(gate422inter0), .b(s_224), .O(gate422inter1));
  and2  gate2117(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2118(.a(s_224), .O(gate422inter3));
  inv1  gate2119(.a(s_225), .O(gate422inter4));
  nand2 gate2120(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2121(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2122(.a(G1039), .O(gate422inter7));
  inv1  gate2123(.a(G1135), .O(gate422inter8));
  nand2 gate2124(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2125(.a(s_225), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2126(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2127(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2128(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate617(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate618(.a(gate424inter0), .b(s_10), .O(gate424inter1));
  and2  gate619(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate620(.a(s_10), .O(gate424inter3));
  inv1  gate621(.a(s_11), .O(gate424inter4));
  nand2 gate622(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate623(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate624(.a(G1042), .O(gate424inter7));
  inv1  gate625(.a(G1138), .O(gate424inter8));
  nand2 gate626(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate627(.a(s_11), .b(gate424inter3), .O(gate424inter10));
  nor2  gate628(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate629(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate630(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1541(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1542(.a(gate445inter0), .b(s_142), .O(gate445inter1));
  and2  gate1543(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1544(.a(s_142), .O(gate445inter3));
  inv1  gate1545(.a(s_143), .O(gate445inter4));
  nand2 gate1546(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1547(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1548(.a(G14), .O(gate445inter7));
  inv1  gate1549(.a(G1171), .O(gate445inter8));
  nand2 gate1550(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1551(.a(s_143), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1552(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1553(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1554(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1807(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1808(.a(gate450inter0), .b(s_180), .O(gate450inter1));
  and2  gate1809(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1810(.a(s_180), .O(gate450inter3));
  inv1  gate1811(.a(s_181), .O(gate450inter4));
  nand2 gate1812(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1813(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1814(.a(G1081), .O(gate450inter7));
  inv1  gate1815(.a(G1177), .O(gate450inter8));
  nand2 gate1816(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1817(.a(s_181), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1818(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1819(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1820(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1149(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1150(.a(gate455inter0), .b(s_86), .O(gate455inter1));
  and2  gate1151(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1152(.a(s_86), .O(gate455inter3));
  inv1  gate1153(.a(s_87), .O(gate455inter4));
  nand2 gate1154(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1155(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1156(.a(G19), .O(gate455inter7));
  inv1  gate1157(.a(G1186), .O(gate455inter8));
  nand2 gate1158(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1159(.a(s_87), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1160(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1161(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1162(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1583(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1584(.a(gate465inter0), .b(s_148), .O(gate465inter1));
  and2  gate1585(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1586(.a(s_148), .O(gate465inter3));
  inv1  gate1587(.a(s_149), .O(gate465inter4));
  nand2 gate1588(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1589(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1590(.a(G24), .O(gate465inter7));
  inv1  gate1591(.a(G1201), .O(gate465inter8));
  nand2 gate1592(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1593(.a(s_149), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1594(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1595(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1596(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1079(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1080(.a(gate466inter0), .b(s_76), .O(gate466inter1));
  and2  gate1081(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1082(.a(s_76), .O(gate466inter3));
  inv1  gate1083(.a(s_77), .O(gate466inter4));
  nand2 gate1084(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1085(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1086(.a(G1105), .O(gate466inter7));
  inv1  gate1087(.a(G1201), .O(gate466inter8));
  nand2 gate1088(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1089(.a(s_77), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1090(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1091(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1092(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1233(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1234(.a(gate468inter0), .b(s_98), .O(gate468inter1));
  and2  gate1235(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1236(.a(s_98), .O(gate468inter3));
  inv1  gate1237(.a(s_99), .O(gate468inter4));
  nand2 gate1238(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1239(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1240(.a(G1108), .O(gate468inter7));
  inv1  gate1241(.a(G1204), .O(gate468inter8));
  nand2 gate1242(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1243(.a(s_99), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1244(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1245(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1246(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1387(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1388(.a(gate470inter0), .b(s_120), .O(gate470inter1));
  and2  gate1389(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1390(.a(s_120), .O(gate470inter3));
  inv1  gate1391(.a(s_121), .O(gate470inter4));
  nand2 gate1392(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1393(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1394(.a(G1111), .O(gate470inter7));
  inv1  gate1395(.a(G1207), .O(gate470inter8));
  nand2 gate1396(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1397(.a(s_121), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1398(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1399(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1400(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1415(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1416(.a(gate471inter0), .b(s_124), .O(gate471inter1));
  and2  gate1417(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1418(.a(s_124), .O(gate471inter3));
  inv1  gate1419(.a(s_125), .O(gate471inter4));
  nand2 gate1420(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1421(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1422(.a(G27), .O(gate471inter7));
  inv1  gate1423(.a(G1210), .O(gate471inter8));
  nand2 gate1424(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1425(.a(s_125), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1426(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1427(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1428(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1009(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1010(.a(gate475inter0), .b(s_66), .O(gate475inter1));
  and2  gate1011(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1012(.a(s_66), .O(gate475inter3));
  inv1  gate1013(.a(s_67), .O(gate475inter4));
  nand2 gate1014(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1015(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1016(.a(G29), .O(gate475inter7));
  inv1  gate1017(.a(G1216), .O(gate475inter8));
  nand2 gate1018(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1019(.a(s_67), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1020(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1021(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1022(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate673(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate674(.a(gate478inter0), .b(s_18), .O(gate478inter1));
  and2  gate675(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate676(.a(s_18), .O(gate478inter3));
  inv1  gate677(.a(s_19), .O(gate478inter4));
  nand2 gate678(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate679(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate680(.a(G1123), .O(gate478inter7));
  inv1  gate681(.a(G1219), .O(gate478inter8));
  nand2 gate682(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate683(.a(s_19), .b(gate478inter3), .O(gate478inter10));
  nor2  gate684(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate685(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate686(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1499(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1500(.a(gate480inter0), .b(s_136), .O(gate480inter1));
  and2  gate1501(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1502(.a(s_136), .O(gate480inter3));
  inv1  gate1503(.a(s_137), .O(gate480inter4));
  nand2 gate1504(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1505(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1506(.a(G1126), .O(gate480inter7));
  inv1  gate1507(.a(G1222), .O(gate480inter8));
  nand2 gate1508(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1509(.a(s_137), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1510(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1511(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1512(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate799(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate800(.a(gate484inter0), .b(s_36), .O(gate484inter1));
  and2  gate801(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate802(.a(s_36), .O(gate484inter3));
  inv1  gate803(.a(s_37), .O(gate484inter4));
  nand2 gate804(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate805(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate806(.a(G1230), .O(gate484inter7));
  inv1  gate807(.a(G1231), .O(gate484inter8));
  nand2 gate808(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate809(.a(s_37), .b(gate484inter3), .O(gate484inter10));
  nor2  gate810(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate811(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate812(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate631(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate632(.a(gate486inter0), .b(s_12), .O(gate486inter1));
  and2  gate633(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate634(.a(s_12), .O(gate486inter3));
  inv1  gate635(.a(s_13), .O(gate486inter4));
  nand2 gate636(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate637(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate638(.a(G1234), .O(gate486inter7));
  inv1  gate639(.a(G1235), .O(gate486inter8));
  nand2 gate640(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate641(.a(s_13), .b(gate486inter3), .O(gate486inter10));
  nor2  gate642(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate643(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate644(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2031(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2032(.a(gate496inter0), .b(s_212), .O(gate496inter1));
  and2  gate2033(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2034(.a(s_212), .O(gate496inter3));
  inv1  gate2035(.a(s_213), .O(gate496inter4));
  nand2 gate2036(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2037(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2038(.a(G1254), .O(gate496inter7));
  inv1  gate2039(.a(G1255), .O(gate496inter8));
  nand2 gate2040(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2041(.a(s_213), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2042(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2043(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2044(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1107(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1108(.a(gate497inter0), .b(s_80), .O(gate497inter1));
  and2  gate1109(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1110(.a(s_80), .O(gate497inter3));
  inv1  gate1111(.a(s_81), .O(gate497inter4));
  nand2 gate1112(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1113(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1114(.a(G1256), .O(gate497inter7));
  inv1  gate1115(.a(G1257), .O(gate497inter8));
  nand2 gate1116(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1117(.a(s_81), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1118(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1119(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1120(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2157(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2158(.a(gate501inter0), .b(s_230), .O(gate501inter1));
  and2  gate2159(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2160(.a(s_230), .O(gate501inter3));
  inv1  gate2161(.a(s_231), .O(gate501inter4));
  nand2 gate2162(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2163(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2164(.a(G1264), .O(gate501inter7));
  inv1  gate2165(.a(G1265), .O(gate501inter8));
  nand2 gate2166(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2167(.a(s_231), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2168(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2169(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2170(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1135(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1136(.a(gate504inter0), .b(s_84), .O(gate504inter1));
  and2  gate1137(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1138(.a(s_84), .O(gate504inter3));
  inv1  gate1139(.a(s_85), .O(gate504inter4));
  nand2 gate1140(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1141(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1142(.a(G1270), .O(gate504inter7));
  inv1  gate1143(.a(G1271), .O(gate504inter8));
  nand2 gate1144(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1145(.a(s_85), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1146(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1147(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1148(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1401(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1402(.a(gate508inter0), .b(s_122), .O(gate508inter1));
  and2  gate1403(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1404(.a(s_122), .O(gate508inter3));
  inv1  gate1405(.a(s_123), .O(gate508inter4));
  nand2 gate1406(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1407(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1408(.a(G1278), .O(gate508inter7));
  inv1  gate1409(.a(G1279), .O(gate508inter8));
  nand2 gate1410(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1411(.a(s_123), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1412(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1413(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1414(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate771(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate772(.a(gate514inter0), .b(s_32), .O(gate514inter1));
  and2  gate773(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate774(.a(s_32), .O(gate514inter3));
  inv1  gate775(.a(s_33), .O(gate514inter4));
  nand2 gate776(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate777(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate778(.a(G1290), .O(gate514inter7));
  inv1  gate779(.a(G1291), .O(gate514inter8));
  nand2 gate780(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate781(.a(s_33), .b(gate514inter3), .O(gate514inter10));
  nor2  gate782(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate783(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate784(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule