module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate743(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate744(.a(gate9inter0), .b(s_28), .O(gate9inter1));
  and2  gate745(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate746(.a(s_28), .O(gate9inter3));
  inv1  gate747(.a(s_29), .O(gate9inter4));
  nand2 gate748(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate749(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate750(.a(G1), .O(gate9inter7));
  inv1  gate751(.a(G2), .O(gate9inter8));
  nand2 gate752(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate753(.a(s_29), .b(gate9inter3), .O(gate9inter10));
  nor2  gate754(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate755(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate756(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1317(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1318(.a(gate10inter0), .b(s_110), .O(gate10inter1));
  and2  gate1319(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1320(.a(s_110), .O(gate10inter3));
  inv1  gate1321(.a(s_111), .O(gate10inter4));
  nand2 gate1322(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1323(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1324(.a(G3), .O(gate10inter7));
  inv1  gate1325(.a(G4), .O(gate10inter8));
  nand2 gate1326(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1327(.a(s_111), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1328(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1329(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1330(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1639(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1640(.a(gate17inter0), .b(s_156), .O(gate17inter1));
  and2  gate1641(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1642(.a(s_156), .O(gate17inter3));
  inv1  gate1643(.a(s_157), .O(gate17inter4));
  nand2 gate1644(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1645(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1646(.a(G17), .O(gate17inter7));
  inv1  gate1647(.a(G18), .O(gate17inter8));
  nand2 gate1648(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1649(.a(s_157), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1650(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1651(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1652(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1107(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1108(.a(gate20inter0), .b(s_80), .O(gate20inter1));
  and2  gate1109(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1110(.a(s_80), .O(gate20inter3));
  inv1  gate1111(.a(s_81), .O(gate20inter4));
  nand2 gate1112(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1113(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1114(.a(G23), .O(gate20inter7));
  inv1  gate1115(.a(G24), .O(gate20inter8));
  nand2 gate1116(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1117(.a(s_81), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1118(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1119(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1120(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate589(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate590(.a(gate21inter0), .b(s_6), .O(gate21inter1));
  and2  gate591(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate592(.a(s_6), .O(gate21inter3));
  inv1  gate593(.a(s_7), .O(gate21inter4));
  nand2 gate594(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate595(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate596(.a(G25), .O(gate21inter7));
  inv1  gate597(.a(G26), .O(gate21inter8));
  nand2 gate598(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate599(.a(s_7), .b(gate21inter3), .O(gate21inter10));
  nor2  gate600(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate601(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate602(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1289(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1290(.a(gate25inter0), .b(s_106), .O(gate25inter1));
  and2  gate1291(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1292(.a(s_106), .O(gate25inter3));
  inv1  gate1293(.a(s_107), .O(gate25inter4));
  nand2 gate1294(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1295(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1296(.a(G1), .O(gate25inter7));
  inv1  gate1297(.a(G5), .O(gate25inter8));
  nand2 gate1298(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1299(.a(s_107), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1300(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1301(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1302(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2003(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2004(.a(gate27inter0), .b(s_208), .O(gate27inter1));
  and2  gate2005(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2006(.a(s_208), .O(gate27inter3));
  inv1  gate2007(.a(s_209), .O(gate27inter4));
  nand2 gate2008(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2009(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2010(.a(G2), .O(gate27inter7));
  inv1  gate2011(.a(G6), .O(gate27inter8));
  nand2 gate2012(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2013(.a(s_209), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2014(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2015(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2016(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1807(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1808(.a(gate30inter0), .b(s_180), .O(gate30inter1));
  and2  gate1809(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1810(.a(s_180), .O(gate30inter3));
  inv1  gate1811(.a(s_181), .O(gate30inter4));
  nand2 gate1812(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1813(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1814(.a(G11), .O(gate30inter7));
  inv1  gate1815(.a(G15), .O(gate30inter8));
  nand2 gate1816(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1817(.a(s_181), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1818(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1819(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1820(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate841(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate842(.a(gate36inter0), .b(s_42), .O(gate36inter1));
  and2  gate843(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate844(.a(s_42), .O(gate36inter3));
  inv1  gate845(.a(s_43), .O(gate36inter4));
  nand2 gate846(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate847(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate848(.a(G26), .O(gate36inter7));
  inv1  gate849(.a(G30), .O(gate36inter8));
  nand2 gate850(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate851(.a(s_43), .b(gate36inter3), .O(gate36inter10));
  nor2  gate852(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate853(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate854(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate659(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate660(.a(gate44inter0), .b(s_16), .O(gate44inter1));
  and2  gate661(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate662(.a(s_16), .O(gate44inter3));
  inv1  gate663(.a(s_17), .O(gate44inter4));
  nand2 gate664(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate665(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate666(.a(G4), .O(gate44inter7));
  inv1  gate667(.a(G269), .O(gate44inter8));
  nand2 gate668(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate669(.a(s_17), .b(gate44inter3), .O(gate44inter10));
  nor2  gate670(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate671(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate672(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1849(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1850(.a(gate49inter0), .b(s_186), .O(gate49inter1));
  and2  gate1851(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1852(.a(s_186), .O(gate49inter3));
  inv1  gate1853(.a(s_187), .O(gate49inter4));
  nand2 gate1854(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1855(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1856(.a(G9), .O(gate49inter7));
  inv1  gate1857(.a(G278), .O(gate49inter8));
  nand2 gate1858(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1859(.a(s_187), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1860(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1861(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1862(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate575(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate576(.a(gate54inter0), .b(s_4), .O(gate54inter1));
  and2  gate577(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate578(.a(s_4), .O(gate54inter3));
  inv1  gate579(.a(s_5), .O(gate54inter4));
  nand2 gate580(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate581(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate582(.a(G14), .O(gate54inter7));
  inv1  gate583(.a(G284), .O(gate54inter8));
  nand2 gate584(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate585(.a(s_5), .b(gate54inter3), .O(gate54inter10));
  nor2  gate586(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate587(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate588(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate715(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate716(.a(gate58inter0), .b(s_24), .O(gate58inter1));
  and2  gate717(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate718(.a(s_24), .O(gate58inter3));
  inv1  gate719(.a(s_25), .O(gate58inter4));
  nand2 gate720(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate721(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate722(.a(G18), .O(gate58inter7));
  inv1  gate723(.a(G290), .O(gate58inter8));
  nand2 gate724(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate725(.a(s_25), .b(gate58inter3), .O(gate58inter10));
  nor2  gate726(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate727(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate728(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1079(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1080(.a(gate61inter0), .b(s_76), .O(gate61inter1));
  and2  gate1081(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1082(.a(s_76), .O(gate61inter3));
  inv1  gate1083(.a(s_77), .O(gate61inter4));
  nand2 gate1084(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1085(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1086(.a(G21), .O(gate61inter7));
  inv1  gate1087(.a(G296), .O(gate61inter8));
  nand2 gate1088(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1089(.a(s_77), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1090(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1091(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1092(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1975(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1976(.a(gate62inter0), .b(s_204), .O(gate62inter1));
  and2  gate1977(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1978(.a(s_204), .O(gate62inter3));
  inv1  gate1979(.a(s_205), .O(gate62inter4));
  nand2 gate1980(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1981(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1982(.a(G22), .O(gate62inter7));
  inv1  gate1983(.a(G296), .O(gate62inter8));
  nand2 gate1984(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1985(.a(s_205), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1986(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1987(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1988(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1653(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1654(.a(gate68inter0), .b(s_158), .O(gate68inter1));
  and2  gate1655(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1656(.a(s_158), .O(gate68inter3));
  inv1  gate1657(.a(s_159), .O(gate68inter4));
  nand2 gate1658(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1659(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1660(.a(G28), .O(gate68inter7));
  inv1  gate1661(.a(G305), .O(gate68inter8));
  nand2 gate1662(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1663(.a(s_159), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1664(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1665(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1666(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate561(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate562(.a(gate69inter0), .b(s_2), .O(gate69inter1));
  and2  gate563(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate564(.a(s_2), .O(gate69inter3));
  inv1  gate565(.a(s_3), .O(gate69inter4));
  nand2 gate566(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate567(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate568(.a(G29), .O(gate69inter7));
  inv1  gate569(.a(G308), .O(gate69inter8));
  nand2 gate570(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate571(.a(s_3), .b(gate69inter3), .O(gate69inter10));
  nor2  gate572(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate573(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate574(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1709(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1710(.a(gate70inter0), .b(s_166), .O(gate70inter1));
  and2  gate1711(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1712(.a(s_166), .O(gate70inter3));
  inv1  gate1713(.a(s_167), .O(gate70inter4));
  nand2 gate1714(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1715(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1716(.a(G30), .O(gate70inter7));
  inv1  gate1717(.a(G308), .O(gate70inter8));
  nand2 gate1718(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1719(.a(s_167), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1720(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1721(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1722(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1037(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1038(.a(gate72inter0), .b(s_70), .O(gate72inter1));
  and2  gate1039(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1040(.a(s_70), .O(gate72inter3));
  inv1  gate1041(.a(s_71), .O(gate72inter4));
  nand2 gate1042(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1043(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1044(.a(G32), .O(gate72inter7));
  inv1  gate1045(.a(G311), .O(gate72inter8));
  nand2 gate1046(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1047(.a(s_71), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1048(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1049(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1050(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1163(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1164(.a(gate74inter0), .b(s_88), .O(gate74inter1));
  and2  gate1165(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1166(.a(s_88), .O(gate74inter3));
  inv1  gate1167(.a(s_89), .O(gate74inter4));
  nand2 gate1168(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1169(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1170(.a(G5), .O(gate74inter7));
  inv1  gate1171(.a(G314), .O(gate74inter8));
  nand2 gate1172(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1173(.a(s_89), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1174(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1175(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1176(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate869(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate870(.a(gate75inter0), .b(s_46), .O(gate75inter1));
  and2  gate871(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate872(.a(s_46), .O(gate75inter3));
  inv1  gate873(.a(s_47), .O(gate75inter4));
  nand2 gate874(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate875(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate876(.a(G9), .O(gate75inter7));
  inv1  gate877(.a(G317), .O(gate75inter8));
  nand2 gate878(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate879(.a(s_47), .b(gate75inter3), .O(gate75inter10));
  nor2  gate880(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate881(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate882(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1359(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1360(.a(gate77inter0), .b(s_116), .O(gate77inter1));
  and2  gate1361(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1362(.a(s_116), .O(gate77inter3));
  inv1  gate1363(.a(s_117), .O(gate77inter4));
  nand2 gate1364(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1365(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1366(.a(G2), .O(gate77inter7));
  inv1  gate1367(.a(G320), .O(gate77inter8));
  nand2 gate1368(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1369(.a(s_117), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1370(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1371(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1372(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1261(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1262(.a(gate80inter0), .b(s_102), .O(gate80inter1));
  and2  gate1263(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1264(.a(s_102), .O(gate80inter3));
  inv1  gate1265(.a(s_103), .O(gate80inter4));
  nand2 gate1266(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1267(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1268(.a(G14), .O(gate80inter7));
  inv1  gate1269(.a(G323), .O(gate80inter8));
  nand2 gate1270(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1271(.a(s_103), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1272(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1273(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1274(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1401(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1402(.a(gate86inter0), .b(s_122), .O(gate86inter1));
  and2  gate1403(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1404(.a(s_122), .O(gate86inter3));
  inv1  gate1405(.a(s_123), .O(gate86inter4));
  nand2 gate1406(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1407(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1408(.a(G8), .O(gate86inter7));
  inv1  gate1409(.a(G332), .O(gate86inter8));
  nand2 gate1410(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1411(.a(s_123), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1412(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1413(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1414(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1737(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1738(.a(gate87inter0), .b(s_170), .O(gate87inter1));
  and2  gate1739(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1740(.a(s_170), .O(gate87inter3));
  inv1  gate1741(.a(s_171), .O(gate87inter4));
  nand2 gate1742(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1743(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1744(.a(G12), .O(gate87inter7));
  inv1  gate1745(.a(G335), .O(gate87inter8));
  nand2 gate1746(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1747(.a(s_171), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1748(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1749(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1750(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1723(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1724(.a(gate99inter0), .b(s_168), .O(gate99inter1));
  and2  gate1725(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1726(.a(s_168), .O(gate99inter3));
  inv1  gate1727(.a(s_169), .O(gate99inter4));
  nand2 gate1728(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1729(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1730(.a(G27), .O(gate99inter7));
  inv1  gate1731(.a(G353), .O(gate99inter8));
  nand2 gate1732(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1733(.a(s_169), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1734(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1735(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1736(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1121(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1122(.a(gate100inter0), .b(s_82), .O(gate100inter1));
  and2  gate1123(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1124(.a(s_82), .O(gate100inter3));
  inv1  gate1125(.a(s_83), .O(gate100inter4));
  nand2 gate1126(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1127(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1128(.a(G31), .O(gate100inter7));
  inv1  gate1129(.a(G353), .O(gate100inter8));
  nand2 gate1130(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1131(.a(s_83), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1132(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1133(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1134(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1443(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1444(.a(gate104inter0), .b(s_128), .O(gate104inter1));
  and2  gate1445(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1446(.a(s_128), .O(gate104inter3));
  inv1  gate1447(.a(s_129), .O(gate104inter4));
  nand2 gate1448(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1449(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1450(.a(G32), .O(gate104inter7));
  inv1  gate1451(.a(G359), .O(gate104inter8));
  nand2 gate1452(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1453(.a(s_129), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1454(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1455(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1456(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate771(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate772(.a(gate122inter0), .b(s_32), .O(gate122inter1));
  and2  gate773(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate774(.a(s_32), .O(gate122inter3));
  inv1  gate775(.a(s_33), .O(gate122inter4));
  nand2 gate776(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate777(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate778(.a(G396), .O(gate122inter7));
  inv1  gate779(.a(G397), .O(gate122inter8));
  nand2 gate780(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate781(.a(s_33), .b(gate122inter3), .O(gate122inter10));
  nor2  gate782(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate783(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate784(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate785(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate786(.a(gate127inter0), .b(s_34), .O(gate127inter1));
  and2  gate787(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate788(.a(s_34), .O(gate127inter3));
  inv1  gate789(.a(s_35), .O(gate127inter4));
  nand2 gate790(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate791(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate792(.a(G406), .O(gate127inter7));
  inv1  gate793(.a(G407), .O(gate127inter8));
  nand2 gate794(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate795(.a(s_35), .b(gate127inter3), .O(gate127inter10));
  nor2  gate796(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate797(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate798(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1415(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1416(.a(gate129inter0), .b(s_124), .O(gate129inter1));
  and2  gate1417(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1418(.a(s_124), .O(gate129inter3));
  inv1  gate1419(.a(s_125), .O(gate129inter4));
  nand2 gate1420(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1421(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1422(.a(G410), .O(gate129inter7));
  inv1  gate1423(.a(G411), .O(gate129inter8));
  nand2 gate1424(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1425(.a(s_125), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1426(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1427(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1428(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate799(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate800(.a(gate136inter0), .b(s_36), .O(gate136inter1));
  and2  gate801(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate802(.a(s_36), .O(gate136inter3));
  inv1  gate803(.a(s_37), .O(gate136inter4));
  nand2 gate804(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate805(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate806(.a(G424), .O(gate136inter7));
  inv1  gate807(.a(G425), .O(gate136inter8));
  nand2 gate808(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate809(.a(s_37), .b(gate136inter3), .O(gate136inter10));
  nor2  gate810(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate811(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate812(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1345(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1346(.a(gate137inter0), .b(s_114), .O(gate137inter1));
  and2  gate1347(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1348(.a(s_114), .O(gate137inter3));
  inv1  gate1349(.a(s_115), .O(gate137inter4));
  nand2 gate1350(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1351(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1352(.a(G426), .O(gate137inter7));
  inv1  gate1353(.a(G429), .O(gate137inter8));
  nand2 gate1354(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1355(.a(s_115), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1356(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1357(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1358(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1513(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1514(.a(gate142inter0), .b(s_138), .O(gate142inter1));
  and2  gate1515(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1516(.a(s_138), .O(gate142inter3));
  inv1  gate1517(.a(s_139), .O(gate142inter4));
  nand2 gate1518(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1519(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1520(.a(G456), .O(gate142inter7));
  inv1  gate1521(.a(G459), .O(gate142inter8));
  nand2 gate1522(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1523(.a(s_139), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1524(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1525(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1526(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1331(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1332(.a(gate145inter0), .b(s_112), .O(gate145inter1));
  and2  gate1333(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1334(.a(s_112), .O(gate145inter3));
  inv1  gate1335(.a(s_113), .O(gate145inter4));
  nand2 gate1336(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1337(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1338(.a(G474), .O(gate145inter7));
  inv1  gate1339(.a(G477), .O(gate145inter8));
  nand2 gate1340(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1341(.a(s_113), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1342(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1343(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1344(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate939(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate940(.a(gate146inter0), .b(s_56), .O(gate146inter1));
  and2  gate941(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate942(.a(s_56), .O(gate146inter3));
  inv1  gate943(.a(s_57), .O(gate146inter4));
  nand2 gate944(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate945(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate946(.a(G480), .O(gate146inter7));
  inv1  gate947(.a(G483), .O(gate146inter8));
  nand2 gate948(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate949(.a(s_57), .b(gate146inter3), .O(gate146inter10));
  nor2  gate950(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate951(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate952(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1233(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1234(.a(gate149inter0), .b(s_98), .O(gate149inter1));
  and2  gate1235(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1236(.a(s_98), .O(gate149inter3));
  inv1  gate1237(.a(s_99), .O(gate149inter4));
  nand2 gate1238(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1239(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1240(.a(G498), .O(gate149inter7));
  inv1  gate1241(.a(G501), .O(gate149inter8));
  nand2 gate1242(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1243(.a(s_99), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1244(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1245(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1246(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate953(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate954(.a(gate154inter0), .b(s_58), .O(gate154inter1));
  and2  gate955(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate956(.a(s_58), .O(gate154inter3));
  inv1  gate957(.a(s_59), .O(gate154inter4));
  nand2 gate958(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate959(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate960(.a(G429), .O(gate154inter7));
  inv1  gate961(.a(G522), .O(gate154inter8));
  nand2 gate962(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate963(.a(s_59), .b(gate154inter3), .O(gate154inter10));
  nor2  gate964(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate965(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate966(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1933(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1934(.a(gate156inter0), .b(s_198), .O(gate156inter1));
  and2  gate1935(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1936(.a(s_198), .O(gate156inter3));
  inv1  gate1937(.a(s_199), .O(gate156inter4));
  nand2 gate1938(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1939(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1940(.a(G435), .O(gate156inter7));
  inv1  gate1941(.a(G525), .O(gate156inter8));
  nand2 gate1942(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1943(.a(s_199), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1944(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1945(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1946(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate617(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate618(.a(gate159inter0), .b(s_10), .O(gate159inter1));
  and2  gate619(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate620(.a(s_10), .O(gate159inter3));
  inv1  gate621(.a(s_11), .O(gate159inter4));
  nand2 gate622(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate623(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate624(.a(G444), .O(gate159inter7));
  inv1  gate625(.a(G531), .O(gate159inter8));
  nand2 gate626(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate627(.a(s_11), .b(gate159inter3), .O(gate159inter10));
  nor2  gate628(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate629(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate630(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1625(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1626(.a(gate165inter0), .b(s_154), .O(gate165inter1));
  and2  gate1627(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1628(.a(s_154), .O(gate165inter3));
  inv1  gate1629(.a(s_155), .O(gate165inter4));
  nand2 gate1630(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1631(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1632(.a(G462), .O(gate165inter7));
  inv1  gate1633(.a(G540), .O(gate165inter8));
  nand2 gate1634(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1635(.a(s_155), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1636(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1637(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1638(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1177(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1178(.a(gate166inter0), .b(s_90), .O(gate166inter1));
  and2  gate1179(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1180(.a(s_90), .O(gate166inter3));
  inv1  gate1181(.a(s_91), .O(gate166inter4));
  nand2 gate1182(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1183(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1184(.a(G465), .O(gate166inter7));
  inv1  gate1185(.a(G540), .O(gate166inter8));
  nand2 gate1186(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1187(.a(s_91), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1188(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1189(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1190(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate995(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate996(.a(gate167inter0), .b(s_64), .O(gate167inter1));
  and2  gate997(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate998(.a(s_64), .O(gate167inter3));
  inv1  gate999(.a(s_65), .O(gate167inter4));
  nand2 gate1000(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1001(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1002(.a(G468), .O(gate167inter7));
  inv1  gate1003(.a(G543), .O(gate167inter8));
  nand2 gate1004(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1005(.a(s_65), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1006(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1007(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1008(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1765(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1766(.a(gate168inter0), .b(s_174), .O(gate168inter1));
  and2  gate1767(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1768(.a(s_174), .O(gate168inter3));
  inv1  gate1769(.a(s_175), .O(gate168inter4));
  nand2 gate1770(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1771(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1772(.a(G471), .O(gate168inter7));
  inv1  gate1773(.a(G543), .O(gate168inter8));
  nand2 gate1774(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1775(.a(s_175), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1776(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1777(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1778(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1065(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1066(.a(gate169inter0), .b(s_74), .O(gate169inter1));
  and2  gate1067(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1068(.a(s_74), .O(gate169inter3));
  inv1  gate1069(.a(s_75), .O(gate169inter4));
  nand2 gate1070(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1071(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1072(.a(G474), .O(gate169inter7));
  inv1  gate1073(.a(G546), .O(gate169inter8));
  nand2 gate1074(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1075(.a(s_75), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1076(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1077(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1078(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1835(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1836(.a(gate171inter0), .b(s_184), .O(gate171inter1));
  and2  gate1837(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1838(.a(s_184), .O(gate171inter3));
  inv1  gate1839(.a(s_185), .O(gate171inter4));
  nand2 gate1840(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1841(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1842(.a(G480), .O(gate171inter7));
  inv1  gate1843(.a(G549), .O(gate171inter8));
  nand2 gate1844(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1845(.a(s_185), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1846(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1847(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1848(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1779(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1780(.a(gate174inter0), .b(s_176), .O(gate174inter1));
  and2  gate1781(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1782(.a(s_176), .O(gate174inter3));
  inv1  gate1783(.a(s_177), .O(gate174inter4));
  nand2 gate1784(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1785(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1786(.a(G489), .O(gate174inter7));
  inv1  gate1787(.a(G552), .O(gate174inter8));
  nand2 gate1788(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1789(.a(s_177), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1790(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1791(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1792(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1275(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1276(.a(gate176inter0), .b(s_104), .O(gate176inter1));
  and2  gate1277(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1278(.a(s_104), .O(gate176inter3));
  inv1  gate1279(.a(s_105), .O(gate176inter4));
  nand2 gate1280(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1281(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1282(.a(G495), .O(gate176inter7));
  inv1  gate1283(.a(G555), .O(gate176inter8));
  nand2 gate1284(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1285(.a(s_105), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1286(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1287(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1288(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1555(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1556(.a(gate184inter0), .b(s_144), .O(gate184inter1));
  and2  gate1557(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1558(.a(s_144), .O(gate184inter3));
  inv1  gate1559(.a(s_145), .O(gate184inter4));
  nand2 gate1560(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1561(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1562(.a(G519), .O(gate184inter7));
  inv1  gate1563(.a(G567), .O(gate184inter8));
  nand2 gate1564(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1565(.a(s_145), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1566(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1567(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1568(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1891(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1892(.a(gate186inter0), .b(s_192), .O(gate186inter1));
  and2  gate1893(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1894(.a(s_192), .O(gate186inter3));
  inv1  gate1895(.a(s_193), .O(gate186inter4));
  nand2 gate1896(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1897(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1898(.a(G572), .O(gate186inter7));
  inv1  gate1899(.a(G573), .O(gate186inter8));
  nand2 gate1900(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1901(.a(s_193), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1902(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1903(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1904(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1947(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1948(.a(gate188inter0), .b(s_200), .O(gate188inter1));
  and2  gate1949(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1950(.a(s_200), .O(gate188inter3));
  inv1  gate1951(.a(s_201), .O(gate188inter4));
  nand2 gate1952(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1953(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1954(.a(G576), .O(gate188inter7));
  inv1  gate1955(.a(G577), .O(gate188inter8));
  nand2 gate1956(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1957(.a(s_201), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1958(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1959(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1960(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1499(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1500(.a(gate189inter0), .b(s_136), .O(gate189inter1));
  and2  gate1501(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1502(.a(s_136), .O(gate189inter3));
  inv1  gate1503(.a(s_137), .O(gate189inter4));
  nand2 gate1504(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1505(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1506(.a(G578), .O(gate189inter7));
  inv1  gate1507(.a(G579), .O(gate189inter8));
  nand2 gate1508(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1509(.a(s_137), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1510(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1511(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1512(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1597(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1598(.a(gate191inter0), .b(s_150), .O(gate191inter1));
  and2  gate1599(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1600(.a(s_150), .O(gate191inter3));
  inv1  gate1601(.a(s_151), .O(gate191inter4));
  nand2 gate1602(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1603(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1604(.a(G582), .O(gate191inter7));
  inv1  gate1605(.a(G583), .O(gate191inter8));
  nand2 gate1606(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1607(.a(s_151), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1608(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1609(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1610(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1821(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1822(.a(gate193inter0), .b(s_182), .O(gate193inter1));
  and2  gate1823(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1824(.a(s_182), .O(gate193inter3));
  inv1  gate1825(.a(s_183), .O(gate193inter4));
  nand2 gate1826(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1827(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1828(.a(G586), .O(gate193inter7));
  inv1  gate1829(.a(G587), .O(gate193inter8));
  nand2 gate1830(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1831(.a(s_183), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1832(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1833(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1834(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1611(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1612(.a(gate195inter0), .b(s_152), .O(gate195inter1));
  and2  gate1613(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1614(.a(s_152), .O(gate195inter3));
  inv1  gate1615(.a(s_153), .O(gate195inter4));
  nand2 gate1616(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1617(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1618(.a(G590), .O(gate195inter7));
  inv1  gate1619(.a(G591), .O(gate195inter8));
  nand2 gate1620(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1621(.a(s_153), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1622(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1623(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1624(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1751(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1752(.a(gate197inter0), .b(s_172), .O(gate197inter1));
  and2  gate1753(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1754(.a(s_172), .O(gate197inter3));
  inv1  gate1755(.a(s_173), .O(gate197inter4));
  nand2 gate1756(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1757(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1758(.a(G594), .O(gate197inter7));
  inv1  gate1759(.a(G595), .O(gate197inter8));
  nand2 gate1760(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1761(.a(s_173), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1762(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1763(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1764(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1009(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1010(.a(gate201inter0), .b(s_66), .O(gate201inter1));
  and2  gate1011(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1012(.a(s_66), .O(gate201inter3));
  inv1  gate1013(.a(s_67), .O(gate201inter4));
  nand2 gate1014(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1015(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1016(.a(G602), .O(gate201inter7));
  inv1  gate1017(.a(G607), .O(gate201inter8));
  nand2 gate1018(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1019(.a(s_67), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1020(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1021(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1022(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate925(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate926(.a(gate210inter0), .b(s_54), .O(gate210inter1));
  and2  gate927(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate928(.a(s_54), .O(gate210inter3));
  inv1  gate929(.a(s_55), .O(gate210inter4));
  nand2 gate930(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate931(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate932(.a(G607), .O(gate210inter7));
  inv1  gate933(.a(G666), .O(gate210inter8));
  nand2 gate934(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate935(.a(s_55), .b(gate210inter3), .O(gate210inter10));
  nor2  gate936(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate937(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate938(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1877(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1878(.a(gate214inter0), .b(s_190), .O(gate214inter1));
  and2  gate1879(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1880(.a(s_190), .O(gate214inter3));
  inv1  gate1881(.a(s_191), .O(gate214inter4));
  nand2 gate1882(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1883(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1884(.a(G612), .O(gate214inter7));
  inv1  gate1885(.a(G672), .O(gate214inter8));
  nand2 gate1886(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1887(.a(s_191), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1888(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1889(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1890(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1219(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1220(.a(gate220inter0), .b(s_96), .O(gate220inter1));
  and2  gate1221(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1222(.a(s_96), .O(gate220inter3));
  inv1  gate1223(.a(s_97), .O(gate220inter4));
  nand2 gate1224(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1225(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1226(.a(G637), .O(gate220inter7));
  inv1  gate1227(.a(G681), .O(gate220inter8));
  nand2 gate1228(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1229(.a(s_97), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1230(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1231(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1232(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate757(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate758(.a(gate224inter0), .b(s_30), .O(gate224inter1));
  and2  gate759(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate760(.a(s_30), .O(gate224inter3));
  inv1  gate761(.a(s_31), .O(gate224inter4));
  nand2 gate762(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate763(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate764(.a(G637), .O(gate224inter7));
  inv1  gate765(.a(G687), .O(gate224inter8));
  nand2 gate766(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate767(.a(s_31), .b(gate224inter3), .O(gate224inter10));
  nor2  gate768(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate769(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate770(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1429(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1430(.a(gate228inter0), .b(s_126), .O(gate228inter1));
  and2  gate1431(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1432(.a(s_126), .O(gate228inter3));
  inv1  gate1433(.a(s_127), .O(gate228inter4));
  nand2 gate1434(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1435(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1436(.a(G696), .O(gate228inter7));
  inv1  gate1437(.a(G697), .O(gate228inter8));
  nand2 gate1438(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1439(.a(s_127), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1440(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1441(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1442(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1863(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1864(.a(gate229inter0), .b(s_188), .O(gate229inter1));
  and2  gate1865(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1866(.a(s_188), .O(gate229inter3));
  inv1  gate1867(.a(s_189), .O(gate229inter4));
  nand2 gate1868(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1869(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1870(.a(G698), .O(gate229inter7));
  inv1  gate1871(.a(G699), .O(gate229inter8));
  nand2 gate1872(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1873(.a(s_189), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1874(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1875(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1876(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1051(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1052(.a(gate231inter0), .b(s_72), .O(gate231inter1));
  and2  gate1053(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1054(.a(s_72), .O(gate231inter3));
  inv1  gate1055(.a(s_73), .O(gate231inter4));
  nand2 gate1056(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1057(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1058(.a(G702), .O(gate231inter7));
  inv1  gate1059(.a(G703), .O(gate231inter8));
  nand2 gate1060(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1061(.a(s_73), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1062(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1063(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1064(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1247(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1248(.a(gate238inter0), .b(s_100), .O(gate238inter1));
  and2  gate1249(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1250(.a(s_100), .O(gate238inter3));
  inv1  gate1251(.a(s_101), .O(gate238inter4));
  nand2 gate1252(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1253(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1254(.a(G257), .O(gate238inter7));
  inv1  gate1255(.a(G709), .O(gate238inter8));
  nand2 gate1256(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1257(.a(s_101), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1258(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1259(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1260(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1919(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1920(.a(gate243inter0), .b(s_196), .O(gate243inter1));
  and2  gate1921(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1922(.a(s_196), .O(gate243inter3));
  inv1  gate1923(.a(s_197), .O(gate243inter4));
  nand2 gate1924(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1925(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1926(.a(G245), .O(gate243inter7));
  inv1  gate1927(.a(G733), .O(gate243inter8));
  nand2 gate1928(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1929(.a(s_197), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1930(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1931(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1932(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate603(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate604(.a(gate244inter0), .b(s_8), .O(gate244inter1));
  and2  gate605(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate606(.a(s_8), .O(gate244inter3));
  inv1  gate607(.a(s_9), .O(gate244inter4));
  nand2 gate608(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate609(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate610(.a(G721), .O(gate244inter7));
  inv1  gate611(.a(G733), .O(gate244inter8));
  nand2 gate612(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate613(.a(s_9), .b(gate244inter3), .O(gate244inter10));
  nor2  gate614(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate615(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate616(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate813(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate814(.a(gate245inter0), .b(s_38), .O(gate245inter1));
  and2  gate815(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate816(.a(s_38), .O(gate245inter3));
  inv1  gate817(.a(s_39), .O(gate245inter4));
  nand2 gate818(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate819(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate820(.a(G248), .O(gate245inter7));
  inv1  gate821(.a(G736), .O(gate245inter8));
  nand2 gate822(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate823(.a(s_39), .b(gate245inter3), .O(gate245inter10));
  nor2  gate824(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate825(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate826(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1135(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1136(.a(gate257inter0), .b(s_84), .O(gate257inter1));
  and2  gate1137(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1138(.a(s_84), .O(gate257inter3));
  inv1  gate1139(.a(s_85), .O(gate257inter4));
  nand2 gate1140(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1141(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1142(.a(G754), .O(gate257inter7));
  inv1  gate1143(.a(G755), .O(gate257inter8));
  nand2 gate1144(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1145(.a(s_85), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1146(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1147(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1148(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1961(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1962(.a(gate286inter0), .b(s_202), .O(gate286inter1));
  and2  gate1963(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1964(.a(s_202), .O(gate286inter3));
  inv1  gate1965(.a(s_203), .O(gate286inter4));
  nand2 gate1966(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1967(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1968(.a(G788), .O(gate286inter7));
  inv1  gate1969(.a(G812), .O(gate286inter8));
  nand2 gate1970(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1971(.a(s_203), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1972(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1973(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1974(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1989(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1990(.a(gate290inter0), .b(s_206), .O(gate290inter1));
  and2  gate1991(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1992(.a(s_206), .O(gate290inter3));
  inv1  gate1993(.a(s_207), .O(gate290inter4));
  nand2 gate1994(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1995(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1996(.a(G820), .O(gate290inter7));
  inv1  gate1997(.a(G821), .O(gate290inter8));
  nand2 gate1998(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1999(.a(s_207), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2000(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2001(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2002(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1205(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1206(.a(gate294inter0), .b(s_94), .O(gate294inter1));
  and2  gate1207(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1208(.a(s_94), .O(gate294inter3));
  inv1  gate1209(.a(s_95), .O(gate294inter4));
  nand2 gate1210(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1211(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1212(.a(G832), .O(gate294inter7));
  inv1  gate1213(.a(G833), .O(gate294inter8));
  nand2 gate1214(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1215(.a(s_95), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1216(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1217(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1218(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1583(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1584(.a(gate387inter0), .b(s_148), .O(gate387inter1));
  and2  gate1585(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1586(.a(s_148), .O(gate387inter3));
  inv1  gate1587(.a(s_149), .O(gate387inter4));
  nand2 gate1588(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1589(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1590(.a(G1), .O(gate387inter7));
  inv1  gate1591(.a(G1036), .O(gate387inter8));
  nand2 gate1592(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1593(.a(s_149), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1594(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1595(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1596(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate883(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate884(.a(gate393inter0), .b(s_48), .O(gate393inter1));
  and2  gate885(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate886(.a(s_48), .O(gate393inter3));
  inv1  gate887(.a(s_49), .O(gate393inter4));
  nand2 gate888(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate889(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate890(.a(G7), .O(gate393inter7));
  inv1  gate891(.a(G1054), .O(gate393inter8));
  nand2 gate892(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate893(.a(s_49), .b(gate393inter3), .O(gate393inter10));
  nor2  gate894(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate895(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate896(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate687(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate688(.a(gate395inter0), .b(s_20), .O(gate395inter1));
  and2  gate689(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate690(.a(s_20), .O(gate395inter3));
  inv1  gate691(.a(s_21), .O(gate395inter4));
  nand2 gate692(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate693(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate694(.a(G9), .O(gate395inter7));
  inv1  gate695(.a(G1060), .O(gate395inter8));
  nand2 gate696(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate697(.a(s_21), .b(gate395inter3), .O(gate395inter10));
  nor2  gate698(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate699(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate700(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate645(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate646(.a(gate399inter0), .b(s_14), .O(gate399inter1));
  and2  gate647(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate648(.a(s_14), .O(gate399inter3));
  inv1  gate649(.a(s_15), .O(gate399inter4));
  nand2 gate650(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate651(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate652(.a(G13), .O(gate399inter7));
  inv1  gate653(.a(G1072), .O(gate399inter8));
  nand2 gate654(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate655(.a(s_15), .b(gate399inter3), .O(gate399inter10));
  nor2  gate656(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate657(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate658(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1569(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1570(.a(gate401inter0), .b(s_146), .O(gate401inter1));
  and2  gate1571(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1572(.a(s_146), .O(gate401inter3));
  inv1  gate1573(.a(s_147), .O(gate401inter4));
  nand2 gate1574(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1575(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1576(.a(G15), .O(gate401inter7));
  inv1  gate1577(.a(G1078), .O(gate401inter8));
  nand2 gate1578(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1579(.a(s_147), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1580(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1581(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1582(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1793(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1794(.a(gate406inter0), .b(s_178), .O(gate406inter1));
  and2  gate1795(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1796(.a(s_178), .O(gate406inter3));
  inv1  gate1797(.a(s_179), .O(gate406inter4));
  nand2 gate1798(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1799(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1800(.a(G20), .O(gate406inter7));
  inv1  gate1801(.a(G1093), .O(gate406inter8));
  nand2 gate1802(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1803(.a(s_179), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1804(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1805(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1806(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate981(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate982(.a(gate411inter0), .b(s_62), .O(gate411inter1));
  and2  gate983(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate984(.a(s_62), .O(gate411inter3));
  inv1  gate985(.a(s_63), .O(gate411inter4));
  nand2 gate986(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate987(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate988(.a(G25), .O(gate411inter7));
  inv1  gate989(.a(G1108), .O(gate411inter8));
  nand2 gate990(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate991(.a(s_63), .b(gate411inter3), .O(gate411inter10));
  nor2  gate992(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate993(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate994(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1023(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1024(.a(gate412inter0), .b(s_68), .O(gate412inter1));
  and2  gate1025(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1026(.a(s_68), .O(gate412inter3));
  inv1  gate1027(.a(s_69), .O(gate412inter4));
  nand2 gate1028(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1029(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1030(.a(G26), .O(gate412inter7));
  inv1  gate1031(.a(G1111), .O(gate412inter8));
  nand2 gate1032(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1033(.a(s_69), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1034(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1035(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1036(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1387(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1388(.a(gate414inter0), .b(s_120), .O(gate414inter1));
  and2  gate1389(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1390(.a(s_120), .O(gate414inter3));
  inv1  gate1391(.a(s_121), .O(gate414inter4));
  nand2 gate1392(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1393(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1394(.a(G28), .O(gate414inter7));
  inv1  gate1395(.a(G1117), .O(gate414inter8));
  nand2 gate1396(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1397(.a(s_121), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1398(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1399(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1400(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate911(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate912(.a(gate416inter0), .b(s_52), .O(gate416inter1));
  and2  gate913(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate914(.a(s_52), .O(gate416inter3));
  inv1  gate915(.a(s_53), .O(gate416inter4));
  nand2 gate916(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate917(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate918(.a(G30), .O(gate416inter7));
  inv1  gate919(.a(G1123), .O(gate416inter8));
  nand2 gate920(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate921(.a(s_53), .b(gate416inter3), .O(gate416inter10));
  nor2  gate922(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate923(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate924(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1905(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1906(.a(gate418inter0), .b(s_194), .O(gate418inter1));
  and2  gate1907(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1908(.a(s_194), .O(gate418inter3));
  inv1  gate1909(.a(s_195), .O(gate418inter4));
  nand2 gate1910(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1911(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1912(.a(G32), .O(gate418inter7));
  inv1  gate1913(.a(G1129), .O(gate418inter8));
  nand2 gate1914(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1915(.a(s_195), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1916(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1917(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1918(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate701(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate702(.a(gate419inter0), .b(s_22), .O(gate419inter1));
  and2  gate703(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate704(.a(s_22), .O(gate419inter3));
  inv1  gate705(.a(s_23), .O(gate419inter4));
  nand2 gate706(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate707(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate708(.a(G1), .O(gate419inter7));
  inv1  gate709(.a(G1132), .O(gate419inter8));
  nand2 gate710(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate711(.a(s_23), .b(gate419inter3), .O(gate419inter10));
  nor2  gate712(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate713(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate714(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1541(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1542(.a(gate422inter0), .b(s_142), .O(gate422inter1));
  and2  gate1543(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1544(.a(s_142), .O(gate422inter3));
  inv1  gate1545(.a(s_143), .O(gate422inter4));
  nand2 gate1546(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1547(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1548(.a(G1039), .O(gate422inter7));
  inv1  gate1549(.a(G1135), .O(gate422inter8));
  nand2 gate1550(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1551(.a(s_143), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1552(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1553(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1554(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1191(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1192(.a(gate428inter0), .b(s_92), .O(gate428inter1));
  and2  gate1193(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1194(.a(s_92), .O(gate428inter3));
  inv1  gate1195(.a(s_93), .O(gate428inter4));
  nand2 gate1196(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1197(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1198(.a(G1048), .O(gate428inter7));
  inv1  gate1199(.a(G1144), .O(gate428inter8));
  nand2 gate1200(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1201(.a(s_93), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1202(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1203(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1204(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate631(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate632(.a(gate431inter0), .b(s_12), .O(gate431inter1));
  and2  gate633(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate634(.a(s_12), .O(gate431inter3));
  inv1  gate635(.a(s_13), .O(gate431inter4));
  nand2 gate636(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate637(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate638(.a(G7), .O(gate431inter7));
  inv1  gate639(.a(G1150), .O(gate431inter8));
  nand2 gate640(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate641(.a(s_13), .b(gate431inter3), .O(gate431inter10));
  nor2  gate642(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate643(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate644(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1457(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1458(.a(gate438inter0), .b(s_130), .O(gate438inter1));
  and2  gate1459(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1460(.a(s_130), .O(gate438inter3));
  inv1  gate1461(.a(s_131), .O(gate438inter4));
  nand2 gate1462(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1463(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1464(.a(G1063), .O(gate438inter7));
  inv1  gate1465(.a(G1159), .O(gate438inter8));
  nand2 gate1466(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1467(.a(s_131), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1468(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1469(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1470(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1149(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1150(.a(gate446inter0), .b(s_86), .O(gate446inter1));
  and2  gate1151(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1152(.a(s_86), .O(gate446inter3));
  inv1  gate1153(.a(s_87), .O(gate446inter4));
  nand2 gate1154(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1155(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1156(.a(G1075), .O(gate446inter7));
  inv1  gate1157(.a(G1171), .O(gate446inter8));
  nand2 gate1158(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1159(.a(s_87), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1160(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1161(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1162(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate897(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate898(.a(gate452inter0), .b(s_50), .O(gate452inter1));
  and2  gate899(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate900(.a(s_50), .O(gate452inter3));
  inv1  gate901(.a(s_51), .O(gate452inter4));
  nand2 gate902(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate903(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate904(.a(G1084), .O(gate452inter7));
  inv1  gate905(.a(G1180), .O(gate452inter8));
  nand2 gate906(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate907(.a(s_51), .b(gate452inter3), .O(gate452inter10));
  nor2  gate908(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate909(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate910(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1373(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1374(.a(gate457inter0), .b(s_118), .O(gate457inter1));
  and2  gate1375(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1376(.a(s_118), .O(gate457inter3));
  inv1  gate1377(.a(s_119), .O(gate457inter4));
  nand2 gate1378(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1379(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1380(.a(G20), .O(gate457inter7));
  inv1  gate1381(.a(G1189), .O(gate457inter8));
  nand2 gate1382(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1383(.a(s_119), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1384(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1385(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1386(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate855(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate856(.a(gate458inter0), .b(s_44), .O(gate458inter1));
  and2  gate857(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate858(.a(s_44), .O(gate458inter3));
  inv1  gate859(.a(s_45), .O(gate458inter4));
  nand2 gate860(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate861(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate862(.a(G1093), .O(gate458inter7));
  inv1  gate863(.a(G1189), .O(gate458inter8));
  nand2 gate864(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate865(.a(s_45), .b(gate458inter3), .O(gate458inter10));
  nor2  gate866(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate867(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate868(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1667(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1668(.a(gate460inter0), .b(s_160), .O(gate460inter1));
  and2  gate1669(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1670(.a(s_160), .O(gate460inter3));
  inv1  gate1671(.a(s_161), .O(gate460inter4));
  nand2 gate1672(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1673(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1674(.a(G1096), .O(gate460inter7));
  inv1  gate1675(.a(G1192), .O(gate460inter8));
  nand2 gate1676(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1677(.a(s_161), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1678(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1679(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1680(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1093(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1094(.a(gate462inter0), .b(s_78), .O(gate462inter1));
  and2  gate1095(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1096(.a(s_78), .O(gate462inter3));
  inv1  gate1097(.a(s_79), .O(gate462inter4));
  nand2 gate1098(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1099(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1100(.a(G1099), .O(gate462inter7));
  inv1  gate1101(.a(G1195), .O(gate462inter8));
  nand2 gate1102(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1103(.a(s_79), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1104(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1105(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1106(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1695(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1696(.a(gate465inter0), .b(s_164), .O(gate465inter1));
  and2  gate1697(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1698(.a(s_164), .O(gate465inter3));
  inv1  gate1699(.a(s_165), .O(gate465inter4));
  nand2 gate1700(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1701(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1702(.a(G24), .O(gate465inter7));
  inv1  gate1703(.a(G1201), .O(gate465inter8));
  nand2 gate1704(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1705(.a(s_165), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1706(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1707(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1708(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1527(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1528(.a(gate471inter0), .b(s_140), .O(gate471inter1));
  and2  gate1529(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1530(.a(s_140), .O(gate471inter3));
  inv1  gate1531(.a(s_141), .O(gate471inter4));
  nand2 gate1532(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1533(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1534(.a(G27), .O(gate471inter7));
  inv1  gate1535(.a(G1210), .O(gate471inter8));
  nand2 gate1536(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1537(.a(s_141), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1538(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1539(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1540(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate729(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate730(.a(gate477inter0), .b(s_26), .O(gate477inter1));
  and2  gate731(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate732(.a(s_26), .O(gate477inter3));
  inv1  gate733(.a(s_27), .O(gate477inter4));
  nand2 gate734(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate735(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate736(.a(G30), .O(gate477inter7));
  inv1  gate737(.a(G1219), .O(gate477inter8));
  nand2 gate738(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate739(.a(s_27), .b(gate477inter3), .O(gate477inter10));
  nor2  gate740(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate741(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate742(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate547(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate548(.a(gate478inter0), .b(s_0), .O(gate478inter1));
  and2  gate549(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate550(.a(s_0), .O(gate478inter3));
  inv1  gate551(.a(s_1), .O(gate478inter4));
  nand2 gate552(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate553(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate554(.a(G1123), .O(gate478inter7));
  inv1  gate555(.a(G1219), .O(gate478inter8));
  nand2 gate556(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate557(.a(s_1), .b(gate478inter3), .O(gate478inter10));
  nor2  gate558(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate559(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate560(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1485(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1486(.a(gate485inter0), .b(s_134), .O(gate485inter1));
  and2  gate1487(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1488(.a(s_134), .O(gate485inter3));
  inv1  gate1489(.a(s_135), .O(gate485inter4));
  nand2 gate1490(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1491(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1492(.a(G1232), .O(gate485inter7));
  inv1  gate1493(.a(G1233), .O(gate485inter8));
  nand2 gate1494(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1495(.a(s_135), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1496(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1497(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1498(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate827(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate828(.a(gate490inter0), .b(s_40), .O(gate490inter1));
  and2  gate829(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate830(.a(s_40), .O(gate490inter3));
  inv1  gate831(.a(s_41), .O(gate490inter4));
  nand2 gate832(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate833(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate834(.a(G1242), .O(gate490inter7));
  inv1  gate835(.a(G1243), .O(gate490inter8));
  nand2 gate836(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate837(.a(s_41), .b(gate490inter3), .O(gate490inter10));
  nor2  gate838(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate839(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate840(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1471(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1472(.a(gate492inter0), .b(s_132), .O(gate492inter1));
  and2  gate1473(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1474(.a(s_132), .O(gate492inter3));
  inv1  gate1475(.a(s_133), .O(gate492inter4));
  nand2 gate1476(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1477(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1478(.a(G1246), .O(gate492inter7));
  inv1  gate1479(.a(G1247), .O(gate492inter8));
  nand2 gate1480(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1481(.a(s_133), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1482(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1483(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1484(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate967(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate968(.a(gate499inter0), .b(s_60), .O(gate499inter1));
  and2  gate969(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate970(.a(s_60), .O(gate499inter3));
  inv1  gate971(.a(s_61), .O(gate499inter4));
  nand2 gate972(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate973(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate974(.a(G1260), .O(gate499inter7));
  inv1  gate975(.a(G1261), .O(gate499inter8));
  nand2 gate976(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate977(.a(s_61), .b(gate499inter3), .O(gate499inter10));
  nor2  gate978(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate979(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate980(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2017(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2018(.a(gate500inter0), .b(s_210), .O(gate500inter1));
  and2  gate2019(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2020(.a(s_210), .O(gate500inter3));
  inv1  gate2021(.a(s_211), .O(gate500inter4));
  nand2 gate2022(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2023(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2024(.a(G1262), .O(gate500inter7));
  inv1  gate2025(.a(G1263), .O(gate500inter8));
  nand2 gate2026(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2027(.a(s_211), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2028(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2029(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2030(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1681(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1682(.a(gate508inter0), .b(s_162), .O(gate508inter1));
  and2  gate1683(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1684(.a(s_162), .O(gate508inter3));
  inv1  gate1685(.a(s_163), .O(gate508inter4));
  nand2 gate1686(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1687(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1688(.a(G1278), .O(gate508inter7));
  inv1  gate1689(.a(G1279), .O(gate508inter8));
  nand2 gate1690(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1691(.a(s_163), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1692(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1693(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1694(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate673(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate674(.a(gate512inter0), .b(s_18), .O(gate512inter1));
  and2  gate675(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate676(.a(s_18), .O(gate512inter3));
  inv1  gate677(.a(s_19), .O(gate512inter4));
  nand2 gate678(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate679(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate680(.a(G1286), .O(gate512inter7));
  inv1  gate681(.a(G1287), .O(gate512inter8));
  nand2 gate682(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate683(.a(s_19), .b(gate512inter3), .O(gate512inter10));
  nor2  gate684(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate685(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate686(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1303(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1304(.a(gate514inter0), .b(s_108), .O(gate514inter1));
  and2  gate1305(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1306(.a(s_108), .O(gate514inter3));
  inv1  gate1307(.a(s_109), .O(gate514inter4));
  nand2 gate1308(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1309(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1310(.a(G1290), .O(gate514inter7));
  inv1  gate1311(.a(G1291), .O(gate514inter8));
  nand2 gate1312(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1313(.a(s_109), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1314(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1315(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1316(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule