module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );

  xor2  gate357(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate358(.a(gate21inter0), .b(s_28), .O(gate21inter1));
  and2  gate359(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate360(.a(s_28), .O(gate21inter3));
  inv1  gate361(.a(s_29), .O(gate21inter4));
  nand2 gate362(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate363(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate364(.a(N14), .O(gate21inter7));
  inv1  gate365(.a(N119), .O(gate21inter8));
  nand2 gate366(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate367(.a(s_29), .b(gate21inter3), .O(gate21inter10));
  nor2  gate368(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate369(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate370(.a(gate21inter12), .b(gate21inter1), .O(N158));

  xor2  gate287(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate288(.a(gate22inter0), .b(s_18), .O(gate22inter1));
  and2  gate289(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate290(.a(s_18), .O(gate22inter3));
  inv1  gate291(.a(s_19), .O(gate22inter4));
  nand2 gate292(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate293(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate294(.a(N122), .O(gate22inter7));
  inv1  gate295(.a(N17), .O(gate22inter8));
  nand2 gate296(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate297(.a(s_19), .b(gate22inter3), .O(gate22inter10));
  nor2  gate298(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate299(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate300(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate301(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate302(.a(gate27inter0), .b(s_20), .O(gate27inter1));
  and2  gate303(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate304(.a(s_20), .O(gate27inter3));
  inv1  gate305(.a(s_21), .O(gate27inter4));
  nand2 gate306(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate307(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate308(.a(N142), .O(gate27inter7));
  inv1  gate309(.a(N82), .O(gate27inter8));
  nand2 gate310(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate311(.a(s_21), .b(gate27inter3), .O(gate27inter10));
  nor2  gate312(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate313(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate314(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate315(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate316(.a(gate29inter0), .b(s_22), .O(gate29inter1));
  and2  gate317(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate318(.a(s_22), .O(gate29inter3));
  inv1  gate319(.a(s_23), .O(gate29inter4));
  nand2 gate320(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate321(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate322(.a(N150), .O(gate29inter7));
  inv1  gate323(.a(N108), .O(gate29inter8));
  nand2 gate324(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate325(.a(s_23), .b(gate29inter3), .O(gate29inter10));
  nor2  gate326(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate327(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate328(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );

  xor2  gate329(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate330(.a(gate42inter0), .b(s_24), .O(gate42inter1));
  and2  gate331(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate332(.a(s_24), .O(gate42inter3));
  inv1  gate333(.a(s_25), .O(gate42inter4));
  nand2 gate334(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate335(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate336(.a(N99), .O(gate42inter7));
  inv1  gate337(.a(N147), .O(gate42inter8));
  nand2 gate338(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate339(.a(s_25), .b(gate42inter3), .O(gate42inter10));
  nor2  gate340(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate341(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate342(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );

  xor2  gate385(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate386(.a(gate51inter0), .b(s_32), .O(gate51inter1));
  and2  gate387(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate388(.a(s_32), .O(gate51inter3));
  inv1  gate389(.a(s_33), .O(gate51inter4));
  nand2 gate390(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate391(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate392(.a(N203), .O(gate51inter7));
  inv1  gate393(.a(N159), .O(gate51inter8));
  nand2 gate394(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate395(.a(s_33), .b(gate51inter3), .O(gate51inter10));
  nor2  gate396(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate397(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate398(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );

  xor2  gate217(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate218(.a(gate55inter0), .b(s_8), .O(gate55inter1));
  and2  gate219(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate220(.a(s_8), .O(gate55inter3));
  inv1  gate221(.a(s_9), .O(gate55inter4));
  nand2 gate222(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate223(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate224(.a(N203), .O(gate55inter7));
  inv1  gate225(.a(N171), .O(gate55inter8));
  nand2 gate226(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate227(.a(s_9), .b(gate55inter3), .O(gate55inter10));
  nor2  gate228(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate229(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate230(.a(gate55inter12), .b(gate55inter1), .O(N239));
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate231(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate232(.a(gate59inter0), .b(s_10), .O(gate59inter1));
  and2  gate233(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate234(.a(s_10), .O(gate59inter3));
  inv1  gate235(.a(s_11), .O(gate59inter4));
  nand2 gate236(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate237(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate238(.a(N203), .O(gate59inter7));
  inv1  gate239(.a(N177), .O(gate59inter8));
  nand2 gate240(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate241(.a(s_11), .b(gate59inter3), .O(gate59inter10));
  nor2  gate242(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate243(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate244(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );

  xor2  gate399(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate400(.a(gate64inter0), .b(s_34), .O(gate64inter1));
  and2  gate401(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate402(.a(s_34), .O(gate64inter3));
  inv1  gate403(.a(s_35), .O(gate64inter4));
  nand2 gate404(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate405(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate406(.a(N213), .O(gate64inter7));
  inv1  gate407(.a(N63), .O(gate64inter8));
  nand2 gate408(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate409(.a(s_35), .b(gate64inter3), .O(gate64inter10));
  nor2  gate410(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate411(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate412(.a(gate64inter12), .b(gate64inter1), .O(N256));

  xor2  gate245(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate246(.a(gate65inter0), .b(s_12), .O(gate65inter1));
  and2  gate247(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate248(.a(s_12), .O(gate65inter3));
  inv1  gate249(.a(s_13), .O(gate65inter4));
  nand2 gate250(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate251(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate252(.a(N213), .O(gate65inter7));
  inv1  gate253(.a(N76), .O(gate65inter8));
  nand2 gate254(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate255(.a(s_13), .b(gate65inter3), .O(gate65inter10));
  nor2  gate256(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate257(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate258(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate343(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate344(.a(gate75inter0), .b(s_26), .O(gate75inter1));
  and2  gate345(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate346(.a(s_26), .O(gate75inter3));
  inv1  gate347(.a(s_27), .O(gate75inter4));
  nand2 gate348(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate349(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate350(.a(N243), .O(gate75inter7));
  inv1  gate351(.a(N193), .O(gate75inter8));
  nand2 gate352(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate353(.a(s_27), .b(gate75inter3), .O(gate75inter10));
  nor2  gate354(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate355(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate356(.a(gate75inter12), .b(gate75inter1), .O(N279));

  xor2  gate427(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate428(.a(gate76inter0), .b(s_38), .O(gate76inter1));
  and2  gate429(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate430(.a(s_38), .O(gate76inter3));
  inv1  gate431(.a(s_39), .O(gate76inter4));
  nand2 gate432(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate433(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate434(.a(N247), .O(gate76inter7));
  inv1  gate435(.a(N195), .O(gate76inter8));
  nand2 gate436(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate437(.a(s_39), .b(gate76inter3), .O(gate76inter10));
  nor2  gate438(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate439(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate440(.a(gate76inter12), .b(gate76inter1), .O(N282));

  xor2  gate371(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate372(.a(gate77inter0), .b(s_30), .O(gate77inter1));
  and2  gate373(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate374(.a(s_30), .O(gate77inter3));
  inv1  gate375(.a(s_31), .O(gate77inter4));
  nand2 gate376(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate377(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate378(.a(N251), .O(gate77inter7));
  inv1  gate379(.a(N197), .O(gate77inter8));
  nand2 gate380(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate381(.a(s_31), .b(gate77inter3), .O(gate77inter10));
  nor2  gate382(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate383(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate384(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );

  xor2  gate259(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate260(.a(gate100inter0), .b(s_14), .O(gate100inter1));
  and2  gate261(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate262(.a(s_14), .O(gate100inter3));
  inv1  gate263(.a(s_15), .O(gate100inter4));
  nand2 gate264(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate265(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate266(.a(N309), .O(gate100inter7));
  inv1  gate267(.a(N264), .O(gate100inter8));
  nand2 gate268(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate269(.a(s_15), .b(gate100inter3), .O(gate100inter10));
  nor2  gate270(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate271(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate272(.a(gate100inter12), .b(gate100inter1), .O(N331));

  xor2  gate413(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate414(.a(gate101inter0), .b(s_36), .O(gate101inter1));
  and2  gate415(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate416(.a(s_36), .O(gate101inter3));
  inv1  gate417(.a(s_37), .O(gate101inter4));
  nand2 gate418(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate419(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate420(.a(N309), .O(gate101inter7));
  inv1  gate421(.a(N267), .O(gate101inter8));
  nand2 gate422(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate423(.a(s_37), .b(gate101inter3), .O(gate101inter10));
  nor2  gate424(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate425(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate426(.a(gate101inter12), .b(gate101inter1), .O(N332));
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate441(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate442(.a(gate103inter0), .b(s_40), .O(gate103inter1));
  and2  gate443(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate444(.a(s_40), .O(gate103inter3));
  inv1  gate445(.a(s_41), .O(gate103inter4));
  nand2 gate446(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate447(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate448(.a(N8), .O(gate103inter7));
  inv1  gate449(.a(N319), .O(gate103inter8));
  nand2 gate450(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate451(.a(s_41), .b(gate103inter3), .O(gate103inter10));
  nor2  gate452(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate453(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate454(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );

  xor2  gate189(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate190(.a(gate107inter0), .b(s_4), .O(gate107inter1));
  and2  gate191(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate192(.a(s_4), .O(gate107inter3));
  inv1  gate193(.a(s_5), .O(gate107inter4));
  nand2 gate194(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate195(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate196(.a(N319), .O(gate107inter7));
  inv1  gate197(.a(N34), .O(gate107inter8));
  nand2 gate198(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate199(.a(s_5), .b(gate107inter3), .O(gate107inter10));
  nor2  gate200(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate201(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate202(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate161(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate162(.a(gate113inter0), .b(s_0), .O(gate113inter1));
  and2  gate163(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate164(.a(s_0), .O(gate113inter3));
  inv1  gate165(.a(s_1), .O(gate113inter4));
  nand2 gate166(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate167(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate168(.a(N319), .O(gate113inter7));
  inv1  gate169(.a(N73), .O(gate113inter8));
  nand2 gate170(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate171(.a(s_1), .b(gate113inter3), .O(gate113inter10));
  nor2  gate172(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate173(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate174(.a(gate113inter12), .b(gate113inter1), .O(N344));

  xor2  gate273(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate274(.a(gate114inter0), .b(s_16), .O(gate114inter1));
  and2  gate275(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate276(.a(s_16), .O(gate114inter3));
  inv1  gate277(.a(s_17), .O(gate114inter4));
  nand2 gate278(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate279(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate280(.a(N319), .O(gate114inter7));
  inv1  gate281(.a(N86), .O(gate114inter8));
  nand2 gate282(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate283(.a(s_17), .b(gate114inter3), .O(gate114inter10));
  nor2  gate284(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate285(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate286(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate203(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate204(.a(gate135inter0), .b(s_6), .O(gate135inter1));
  and2  gate205(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate206(.a(s_6), .O(gate135inter3));
  inv1  gate207(.a(s_7), .O(gate135inter4));
  nand2 gate208(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate209(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate210(.a(N360), .O(gate135inter7));
  inv1  gate211(.a(N92), .O(gate135inter8));
  nand2 gate212(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate213(.a(s_7), .b(gate135inter3), .O(gate135inter10));
  nor2  gate214(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate215(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate216(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );

  xor2  gate175(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate176(.a(gate137inter0), .b(s_2), .O(gate137inter1));
  and2  gate177(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate178(.a(s_2), .O(gate137inter3));
  inv1  gate179(.a(s_3), .O(gate137inter4));
  nand2 gate180(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate181(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate182(.a(N360), .O(gate137inter7));
  inv1  gate183(.a(N115), .O(gate137inter8));
  nand2 gate184(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate185(.a(s_3), .b(gate137inter3), .O(gate137inter10));
  nor2  gate186(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate187(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate188(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule