module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate371(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate372(.a(gate3inter0), .b(s_24), .O(gate3inter1));
  and2  gate373(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate374(.a(s_24), .O(gate3inter3));
  inv1  gate375(.a(s_25), .O(gate3inter4));
  nand2 gate376(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate377(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate378(.a(N17), .O(gate3inter7));
  inv1  gate379(.a(N21), .O(gate3inter8));
  nand2 gate380(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate381(.a(s_25), .b(gate3inter3), .O(gate3inter10));
  nor2  gate382(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate383(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate384(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );

  xor2  gate385(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate386(.a(gate5inter0), .b(s_26), .O(gate5inter1));
  and2  gate387(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate388(.a(s_26), .O(gate5inter3));
  inv1  gate389(.a(s_27), .O(gate5inter4));
  nand2 gate390(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate391(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate392(.a(N33), .O(gate5inter7));
  inv1  gate393(.a(N37), .O(gate5inter8));
  nand2 gate394(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate395(.a(s_27), .b(gate5inter3), .O(gate5inter10));
  nor2  gate396(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate397(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate398(.a(gate5inter12), .b(gate5inter1), .O(N254));

  xor2  gate539(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate540(.a(gate6inter0), .b(s_48), .O(gate6inter1));
  and2  gate541(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate542(.a(s_48), .O(gate6inter3));
  inv1  gate543(.a(s_49), .O(gate6inter4));
  nand2 gate544(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate545(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate546(.a(N41), .O(gate6inter7));
  inv1  gate547(.a(N45), .O(gate6inter8));
  nand2 gate548(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate549(.a(s_49), .b(gate6inter3), .O(gate6inter10));
  nor2  gate550(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate551(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate552(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );

  xor2  gate413(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate414(.a(gate9inter0), .b(s_30), .O(gate9inter1));
  and2  gate415(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate416(.a(s_30), .O(gate9inter3));
  inv1  gate417(.a(s_31), .O(gate9inter4));
  nand2 gate418(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate419(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate420(.a(N65), .O(gate9inter7));
  inv1  gate421(.a(N69), .O(gate9inter8));
  nand2 gate422(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate423(.a(s_31), .b(gate9inter3), .O(gate9inter10));
  nor2  gate424(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate425(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate426(.a(gate9inter12), .b(gate9inter1), .O(N258));
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );

  xor2  gate287(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate288(.a(gate16inter0), .b(s_12), .O(gate16inter1));
  and2  gate289(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate290(.a(s_12), .O(gate16inter3));
  inv1  gate291(.a(s_13), .O(gate16inter4));
  nand2 gate292(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate293(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate294(.a(N121), .O(gate16inter7));
  inv1  gate295(.a(N125), .O(gate16inter8));
  nand2 gate296(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate297(.a(s_13), .b(gate16inter3), .O(gate16inter10));
  nor2  gate298(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate299(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate300(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );

  xor2  gate483(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate484(.a(gate29inter0), .b(s_40), .O(gate29inter1));
  and2  gate485(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate486(.a(s_40), .O(gate29inter3));
  inv1  gate487(.a(s_41), .O(gate29inter4));
  nand2 gate488(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate489(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate490(.a(N9), .O(gate29inter7));
  inv1  gate491(.a(N25), .O(gate29inter8));
  nand2 gate492(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate493(.a(s_41), .b(gate29inter3), .O(gate29inter10));
  nor2  gate494(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate495(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate496(.a(gate29inter12), .b(gate29inter1), .O(N278));

  xor2  gate553(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate554(.a(gate30inter0), .b(s_50), .O(gate30inter1));
  and2  gate555(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate556(.a(s_50), .O(gate30inter3));
  inv1  gate557(.a(s_51), .O(gate30inter4));
  nand2 gate558(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate559(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate560(.a(N41), .O(gate30inter7));
  inv1  gate561(.a(N57), .O(gate30inter8));
  nand2 gate562(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate563(.a(s_51), .b(gate30inter3), .O(gate30inter10));
  nor2  gate564(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate565(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate566(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );

  xor2  gate357(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate358(.a(gate33inter0), .b(s_22), .O(gate33inter1));
  and2  gate359(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate360(.a(s_22), .O(gate33inter3));
  inv1  gate361(.a(s_23), .O(gate33inter4));
  nand2 gate362(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate363(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate364(.a(N65), .O(gate33inter7));
  inv1  gate365(.a(N81), .O(gate33inter8));
  nand2 gate366(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate367(.a(s_23), .b(gate33inter3), .O(gate33inter10));
  nor2  gate368(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate369(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate370(.a(gate33inter12), .b(gate33inter1), .O(N282));
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );

  xor2  gate651(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate652(.a(gate38inter0), .b(s_64), .O(gate38inter1));
  and2  gate653(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate654(.a(s_64), .O(gate38inter3));
  inv1  gate655(.a(s_65), .O(gate38inter4));
  nand2 gate656(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate657(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate658(.a(N105), .O(gate38inter7));
  inv1  gate659(.a(N121), .O(gate38inter8));
  nand2 gate660(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate661(.a(s_65), .b(gate38inter3), .O(gate38inter10));
  nor2  gate662(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate663(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate664(.a(gate38inter12), .b(gate38inter1), .O(N287));
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );

  xor2  gate511(.a(N251), .b(N250), .O(gate41inter0));
  nand2 gate512(.a(gate41inter0), .b(s_44), .O(gate41inter1));
  and2  gate513(.a(N251), .b(N250), .O(gate41inter2));
  inv1  gate514(.a(s_44), .O(gate41inter3));
  inv1  gate515(.a(s_45), .O(gate41inter4));
  nand2 gate516(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate517(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate518(.a(N250), .O(gate41inter7));
  inv1  gate519(.a(N251), .O(gate41inter8));
  nand2 gate520(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate521(.a(s_45), .b(gate41inter3), .O(gate41inter10));
  nor2  gate522(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate523(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate524(.a(gate41inter12), .b(gate41inter1), .O(N290));
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );

  xor2  gate301(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate302(.a(gate45inter0), .b(s_14), .O(gate45inter1));
  and2  gate303(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate304(.a(s_14), .O(gate45inter3));
  inv1  gate305(.a(s_15), .O(gate45inter4));
  nand2 gate306(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate307(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate308(.a(N258), .O(gate45inter7));
  inv1  gate309(.a(N259), .O(gate45inter8));
  nand2 gate310(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate311(.a(s_15), .b(gate45inter3), .O(gate45inter10));
  nor2  gate312(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate313(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate314(.a(gate45inter12), .b(gate45inter1), .O(N302));

  xor2  gate497(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate498(.a(gate46inter0), .b(s_42), .O(gate46inter1));
  and2  gate499(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate500(.a(s_42), .O(gate46inter3));
  inv1  gate501(.a(s_43), .O(gate46inter4));
  nand2 gate502(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate503(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate504(.a(N260), .O(gate46inter7));
  inv1  gate505(.a(N261), .O(gate46inter8));
  nand2 gate506(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate507(.a(s_43), .b(gate46inter3), .O(gate46inter10));
  nor2  gate508(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate509(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate510(.a(gate46inter12), .b(gate46inter1), .O(N305));
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate203(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate204(.a(gate50inter0), .b(s_0), .O(gate50inter1));
  and2  gate205(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate206(.a(s_0), .O(gate50inter3));
  inv1  gate207(.a(s_1), .O(gate50inter4));
  nand2 gate208(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate209(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate210(.a(N276), .O(gate50inter7));
  inv1  gate211(.a(N277), .O(gate50inter8));
  nand2 gate212(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate213(.a(s_1), .b(gate50inter3), .O(gate50inter10));
  nor2  gate214(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate215(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate216(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate245(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate246(.a(gate55inter0), .b(s_6), .O(gate55inter1));
  and2  gate247(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate248(.a(s_6), .O(gate55inter3));
  inv1  gate249(.a(s_7), .O(gate55inter4));
  nand2 gate250(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate251(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate252(.a(N286), .O(gate55inter7));
  inv1  gate253(.a(N287), .O(gate55inter8));
  nand2 gate254(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate255(.a(s_7), .b(gate55inter3), .O(gate55inter10));
  nor2  gate256(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate257(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate258(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );

  xor2  gate679(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate680(.a(gate58inter0), .b(s_68), .O(gate58inter1));
  and2  gate681(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate682(.a(s_68), .O(gate58inter3));
  inv1  gate683(.a(s_69), .O(gate58inter4));
  nand2 gate684(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate685(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate686(.a(N296), .O(gate58inter7));
  inv1  gate687(.a(N299), .O(gate58inter8));
  nand2 gate688(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate689(.a(s_69), .b(gate58inter3), .O(gate58inter10));
  nor2  gate690(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate691(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate692(.a(gate58inter12), .b(gate58inter1), .O(N339));
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate525(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate526(.a(gate65inter0), .b(s_46), .O(gate65inter1));
  and2  gate527(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate528(.a(s_46), .O(gate65inter3));
  inv1  gate529(.a(s_47), .O(gate65inter4));
  nand2 gate530(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate531(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate532(.a(N266), .O(gate65inter7));
  inv1  gate533(.a(N342), .O(gate65inter8));
  nand2 gate534(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate535(.a(s_47), .b(gate65inter3), .O(gate65inter10));
  nor2  gate536(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate537(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate538(.a(gate65inter12), .b(gate65inter1), .O(N346));

  xor2  gate623(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate624(.a(gate66inter0), .b(s_60), .O(gate66inter1));
  and2  gate625(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate626(.a(s_60), .O(gate66inter3));
  inv1  gate627(.a(s_61), .O(gate66inter4));
  nand2 gate628(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate629(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate630(.a(N267), .O(gate66inter7));
  inv1  gate631(.a(N343), .O(gate66inter8));
  nand2 gate632(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate633(.a(s_61), .b(gate66inter3), .O(gate66inter10));
  nor2  gate634(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate635(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate636(.a(gate66inter12), .b(gate66inter1), .O(N347));
xor2 gate67( .a(N268), .b(N344), .O(N348) );

  xor2  gate469(.a(N345), .b(N269), .O(gate68inter0));
  nand2 gate470(.a(gate68inter0), .b(s_38), .O(gate68inter1));
  and2  gate471(.a(N345), .b(N269), .O(gate68inter2));
  inv1  gate472(.a(s_38), .O(gate68inter3));
  inv1  gate473(.a(s_39), .O(gate68inter4));
  nand2 gate474(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate475(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate476(.a(N269), .O(gate68inter7));
  inv1  gate477(.a(N345), .O(gate68inter8));
  nand2 gate478(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate479(.a(s_39), .b(gate68inter3), .O(gate68inter10));
  nor2  gate480(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate481(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate482(.a(gate68inter12), .b(gate68inter1), .O(N349));
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );

  xor2  gate693(.a(N340), .b(N272), .O(gate71inter0));
  nand2 gate694(.a(gate71inter0), .b(s_70), .O(gate71inter1));
  and2  gate695(.a(N340), .b(N272), .O(gate71inter2));
  inv1  gate696(.a(s_70), .O(gate71inter3));
  inv1  gate697(.a(s_71), .O(gate71inter4));
  nand2 gate698(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate699(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate700(.a(N272), .O(gate71inter7));
  inv1  gate701(.a(N340), .O(gate71inter8));
  nand2 gate702(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate703(.a(s_71), .b(gate71inter3), .O(gate71inter10));
  nor2  gate704(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate705(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate706(.a(gate71inter12), .b(gate71inter1), .O(N352));

  xor2  gate315(.a(N341), .b(N273), .O(gate72inter0));
  nand2 gate316(.a(gate72inter0), .b(s_16), .O(gate72inter1));
  and2  gate317(.a(N341), .b(N273), .O(gate72inter2));
  inv1  gate318(.a(s_16), .O(gate72inter3));
  inv1  gate319(.a(s_17), .O(gate72inter4));
  nand2 gate320(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate321(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate322(.a(N273), .O(gate72inter7));
  inv1  gate323(.a(N341), .O(gate72inter8));
  nand2 gate324(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate325(.a(s_17), .b(gate72inter3), .O(gate72inter10));
  nor2  gate326(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate327(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate328(.a(gate72inter12), .b(gate72inter1), .O(N353));
xor2 gate73( .a(N314), .b(N346), .O(N354) );

  xor2  gate455(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate456(.a(gate74inter0), .b(s_36), .O(gate74inter1));
  and2  gate457(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate458(.a(s_36), .O(gate74inter3));
  inv1  gate459(.a(s_37), .O(gate74inter4));
  nand2 gate460(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate461(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate462(.a(N315), .O(gate74inter7));
  inv1  gate463(.a(N347), .O(gate74inter8));
  nand2 gate464(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate465(.a(s_37), .b(gate74inter3), .O(gate74inter10));
  nor2  gate466(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate467(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate468(.a(gate74inter12), .b(gate74inter1), .O(N367));

  xor2  gate329(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate330(.a(gate75inter0), .b(s_18), .O(gate75inter1));
  and2  gate331(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate332(.a(s_18), .O(gate75inter3));
  inv1  gate333(.a(s_19), .O(gate75inter4));
  nand2 gate334(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate335(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate336(.a(N316), .O(gate75inter7));
  inv1  gate337(.a(N348), .O(gate75inter8));
  nand2 gate338(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate339(.a(s_19), .b(gate75inter3), .O(gate75inter10));
  nor2  gate340(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate341(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate342(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );

  xor2  gate441(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate442(.a(gate77inter0), .b(s_34), .O(gate77inter1));
  and2  gate443(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate444(.a(s_34), .O(gate77inter3));
  inv1  gate445(.a(s_35), .O(gate77inter4));
  nand2 gate446(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate447(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate448(.a(N318), .O(gate77inter7));
  inv1  gate449(.a(N350), .O(gate77inter8));
  nand2 gate450(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate451(.a(s_35), .b(gate77inter3), .O(gate77inter10));
  nor2  gate452(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate453(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate454(.a(gate77inter12), .b(gate77inter1), .O(N406));

  xor2  gate581(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate582(.a(gate78inter0), .b(s_54), .O(gate78inter1));
  and2  gate583(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate584(.a(s_54), .O(gate78inter3));
  inv1  gate585(.a(s_55), .O(gate78inter4));
  nand2 gate586(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate587(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate588(.a(N319), .O(gate78inter7));
  inv1  gate589(.a(N351), .O(gate78inter8));
  nand2 gate590(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate591(.a(s_55), .b(gate78inter3), .O(gate78inter10));
  nor2  gate592(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate593(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate594(.a(gate78inter12), .b(gate78inter1), .O(N419));

  xor2  gate637(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate638(.a(gate79inter0), .b(s_62), .O(gate79inter1));
  and2  gate639(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate640(.a(s_62), .O(gate79inter3));
  inv1  gate641(.a(s_63), .O(gate79inter4));
  nand2 gate642(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate643(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate644(.a(N320), .O(gate79inter7));
  inv1  gate645(.a(N352), .O(gate79inter8));
  nand2 gate646(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate647(.a(s_63), .b(gate79inter3), .O(gate79inter10));
  nor2  gate648(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate649(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate650(.a(gate79inter12), .b(gate79inter1), .O(N432));

  xor2  gate399(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate400(.a(gate80inter0), .b(s_28), .O(gate80inter1));
  and2  gate401(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate402(.a(s_28), .O(gate80inter3));
  inv1  gate403(.a(s_29), .O(gate80inter4));
  nand2 gate404(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate405(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate406(.a(N321), .O(gate80inter7));
  inv1  gate407(.a(N353), .O(gate80inter8));
  nand2 gate408(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate409(.a(s_29), .b(gate80inter3), .O(gate80inter10));
  nor2  gate410(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate411(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate412(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );

  xor2  gate595(.a(N692), .b(N1), .O(gate171inter0));
  nand2 gate596(.a(gate171inter0), .b(s_56), .O(gate171inter1));
  and2  gate597(.a(N692), .b(N1), .O(gate171inter2));
  inv1  gate598(.a(s_56), .O(gate171inter3));
  inv1  gate599(.a(s_57), .O(gate171inter4));
  nand2 gate600(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate601(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate602(.a(N1), .O(gate171inter7));
  inv1  gate603(.a(N692), .O(gate171inter8));
  nand2 gate604(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate605(.a(s_57), .b(gate171inter3), .O(gate171inter10));
  nor2  gate606(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate607(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate608(.a(gate171inter12), .b(gate171inter1), .O(N724));
xor2 gate172( .a(N5), .b(N693), .O(N725) );

  xor2  gate427(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate428(.a(gate173inter0), .b(s_32), .O(gate173inter1));
  and2  gate429(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate430(.a(s_32), .O(gate173inter3));
  inv1  gate431(.a(s_33), .O(gate173inter4));
  nand2 gate432(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate433(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate434(.a(N9), .O(gate173inter7));
  inv1  gate435(.a(N694), .O(gate173inter8));
  nand2 gate436(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate437(.a(s_33), .b(gate173inter3), .O(gate173inter10));
  nor2  gate438(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate439(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate440(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );

  xor2  gate273(.a(N696), .b(N17), .O(gate175inter0));
  nand2 gate274(.a(gate175inter0), .b(s_10), .O(gate175inter1));
  and2  gate275(.a(N696), .b(N17), .O(gate175inter2));
  inv1  gate276(.a(s_10), .O(gate175inter3));
  inv1  gate277(.a(s_11), .O(gate175inter4));
  nand2 gate278(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate279(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate280(.a(N17), .O(gate175inter7));
  inv1  gate281(.a(N696), .O(gate175inter8));
  nand2 gate282(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate283(.a(s_11), .b(gate175inter3), .O(gate175inter10));
  nor2  gate284(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate285(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate286(.a(gate175inter12), .b(gate175inter1), .O(N728));
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );

  xor2  gate259(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate260(.a(gate178inter0), .b(s_8), .O(gate178inter1));
  and2  gate261(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate262(.a(s_8), .O(gate178inter3));
  inv1  gate263(.a(s_9), .O(gate178inter4));
  nand2 gate264(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate265(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate266(.a(N29), .O(gate178inter7));
  inv1  gate267(.a(N699), .O(gate178inter8));
  nand2 gate268(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate269(.a(s_9), .b(gate178inter3), .O(gate178inter10));
  nor2  gate270(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate271(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate272(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate217(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate218(.a(gate186inter0), .b(s_2), .O(gate186inter1));
  and2  gate219(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate220(.a(s_2), .O(gate186inter3));
  inv1  gate221(.a(s_3), .O(gate186inter4));
  nand2 gate222(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate223(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate224(.a(N61), .O(gate186inter7));
  inv1  gate225(.a(N707), .O(gate186inter8));
  nand2 gate226(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate227(.a(s_3), .b(gate186inter3), .O(gate186inter10));
  nor2  gate228(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate229(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate230(.a(gate186inter12), .b(gate186inter1), .O(N739));
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );

  xor2  gate665(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate666(.a(gate191inter0), .b(s_66), .O(gate191inter1));
  and2  gate667(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate668(.a(s_66), .O(gate191inter3));
  inv1  gate669(.a(s_67), .O(gate191inter4));
  nand2 gate670(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate671(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate672(.a(N81), .O(gate191inter7));
  inv1  gate673(.a(N712), .O(gate191inter8));
  nand2 gate674(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate675(.a(s_67), .b(gate191inter3), .O(gate191inter10));
  nor2  gate676(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate677(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate678(.a(gate191inter12), .b(gate191inter1), .O(N744));
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );

  xor2  gate231(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate232(.a(gate194inter0), .b(s_4), .O(gate194inter1));
  and2  gate233(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate234(.a(s_4), .O(gate194inter3));
  inv1  gate235(.a(s_5), .O(gate194inter4));
  nand2 gate236(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate237(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate238(.a(N93), .O(gate194inter7));
  inv1  gate239(.a(N715), .O(gate194inter8));
  nand2 gate240(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate241(.a(s_5), .b(gate194inter3), .O(gate194inter10));
  nor2  gate242(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate243(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate244(.a(gate194inter12), .b(gate194inter1), .O(N747));

  xor2  gate343(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate344(.a(gate195inter0), .b(s_20), .O(gate195inter1));
  and2  gate345(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate346(.a(s_20), .O(gate195inter3));
  inv1  gate347(.a(s_21), .O(gate195inter4));
  nand2 gate348(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate349(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate350(.a(N97), .O(gate195inter7));
  inv1  gate351(.a(N716), .O(gate195inter8));
  nand2 gate352(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate353(.a(s_21), .b(gate195inter3), .O(gate195inter10));
  nor2  gate354(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate355(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate356(.a(gate195inter12), .b(gate195inter1), .O(N748));
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );

  xor2  gate567(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate568(.a(gate199inter0), .b(s_52), .O(gate199inter1));
  and2  gate569(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate570(.a(s_52), .O(gate199inter3));
  inv1  gate571(.a(s_53), .O(gate199inter4));
  nand2 gate572(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate573(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate574(.a(N113), .O(gate199inter7));
  inv1  gate575(.a(N720), .O(gate199inter8));
  nand2 gate576(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate577(.a(s_53), .b(gate199inter3), .O(gate199inter10));
  nor2  gate578(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate579(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate580(.a(gate199inter12), .b(gate199inter1), .O(N752));
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate609(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate610(.a(gate201inter0), .b(s_58), .O(gate201inter1));
  and2  gate611(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate612(.a(s_58), .O(gate201inter3));
  inv1  gate613(.a(s_59), .O(gate201inter4));
  nand2 gate614(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate615(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate616(.a(N121), .O(gate201inter7));
  inv1  gate617(.a(N722), .O(gate201inter8));
  nand2 gate618(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate619(.a(s_59), .b(gate201inter3), .O(gate201inter10));
  nor2  gate620(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate621(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate622(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule