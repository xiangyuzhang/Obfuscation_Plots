module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1597(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1598(.a(gate13inter0), .b(s_150), .O(gate13inter1));
  and2  gate1599(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1600(.a(s_150), .O(gate13inter3));
  inv1  gate1601(.a(s_151), .O(gate13inter4));
  nand2 gate1602(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1603(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1604(.a(G9), .O(gate13inter7));
  inv1  gate1605(.a(G10), .O(gate13inter8));
  nand2 gate1606(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1607(.a(s_151), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1608(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1609(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1610(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate561(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate562(.a(gate18inter0), .b(s_2), .O(gate18inter1));
  and2  gate563(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate564(.a(s_2), .O(gate18inter3));
  inv1  gate565(.a(s_3), .O(gate18inter4));
  nand2 gate566(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate567(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate568(.a(G19), .O(gate18inter7));
  inv1  gate569(.a(G20), .O(gate18inter8));
  nand2 gate570(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate571(.a(s_3), .b(gate18inter3), .O(gate18inter10));
  nor2  gate572(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate573(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate574(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate701(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate702(.a(gate22inter0), .b(s_22), .O(gate22inter1));
  and2  gate703(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate704(.a(s_22), .O(gate22inter3));
  inv1  gate705(.a(s_23), .O(gate22inter4));
  nand2 gate706(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate707(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate708(.a(G27), .O(gate22inter7));
  inv1  gate709(.a(G28), .O(gate22inter8));
  nand2 gate710(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate711(.a(s_23), .b(gate22inter3), .O(gate22inter10));
  nor2  gate712(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate713(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate714(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate981(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate982(.a(gate25inter0), .b(s_62), .O(gate25inter1));
  and2  gate983(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate984(.a(s_62), .O(gate25inter3));
  inv1  gate985(.a(s_63), .O(gate25inter4));
  nand2 gate986(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate987(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate988(.a(G1), .O(gate25inter7));
  inv1  gate989(.a(G5), .O(gate25inter8));
  nand2 gate990(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate991(.a(s_63), .b(gate25inter3), .O(gate25inter10));
  nor2  gate992(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate993(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate994(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1611(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1612(.a(gate29inter0), .b(s_152), .O(gate29inter1));
  and2  gate1613(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1614(.a(s_152), .O(gate29inter3));
  inv1  gate1615(.a(s_153), .O(gate29inter4));
  nand2 gate1616(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1617(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1618(.a(G3), .O(gate29inter7));
  inv1  gate1619(.a(G7), .O(gate29inter8));
  nand2 gate1620(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1621(.a(s_153), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1622(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1623(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1624(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate855(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate856(.a(gate36inter0), .b(s_44), .O(gate36inter1));
  and2  gate857(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate858(.a(s_44), .O(gate36inter3));
  inv1  gate859(.a(s_45), .O(gate36inter4));
  nand2 gate860(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate861(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate862(.a(G26), .O(gate36inter7));
  inv1  gate863(.a(G30), .O(gate36inter8));
  nand2 gate864(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate865(.a(s_45), .b(gate36inter3), .O(gate36inter10));
  nor2  gate866(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate867(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate868(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate841(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate842(.a(gate38inter0), .b(s_42), .O(gate38inter1));
  and2  gate843(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate844(.a(s_42), .O(gate38inter3));
  inv1  gate845(.a(s_43), .O(gate38inter4));
  nand2 gate846(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate847(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate848(.a(G27), .O(gate38inter7));
  inv1  gate849(.a(G31), .O(gate38inter8));
  nand2 gate850(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate851(.a(s_43), .b(gate38inter3), .O(gate38inter10));
  nor2  gate852(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate853(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate854(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1653(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1654(.a(gate39inter0), .b(s_158), .O(gate39inter1));
  and2  gate1655(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1656(.a(s_158), .O(gate39inter3));
  inv1  gate1657(.a(s_159), .O(gate39inter4));
  nand2 gate1658(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1659(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1660(.a(G20), .O(gate39inter7));
  inv1  gate1661(.a(G24), .O(gate39inter8));
  nand2 gate1662(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1663(.a(s_159), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1664(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1665(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1666(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1667(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1668(.a(gate40inter0), .b(s_160), .O(gate40inter1));
  and2  gate1669(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1670(.a(s_160), .O(gate40inter3));
  inv1  gate1671(.a(s_161), .O(gate40inter4));
  nand2 gate1672(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1673(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1674(.a(G28), .O(gate40inter7));
  inv1  gate1675(.a(G32), .O(gate40inter8));
  nand2 gate1676(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1677(.a(s_161), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1678(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1679(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1680(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1275(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1276(.a(gate44inter0), .b(s_104), .O(gate44inter1));
  and2  gate1277(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1278(.a(s_104), .O(gate44inter3));
  inv1  gate1279(.a(s_105), .O(gate44inter4));
  nand2 gate1280(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1281(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1282(.a(G4), .O(gate44inter7));
  inv1  gate1283(.a(G269), .O(gate44inter8));
  nand2 gate1284(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1285(.a(s_105), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1286(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1287(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1288(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1569(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1570(.a(gate54inter0), .b(s_146), .O(gate54inter1));
  and2  gate1571(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1572(.a(s_146), .O(gate54inter3));
  inv1  gate1573(.a(s_147), .O(gate54inter4));
  nand2 gate1574(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1575(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1576(.a(G14), .O(gate54inter7));
  inv1  gate1577(.a(G284), .O(gate54inter8));
  nand2 gate1578(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1579(.a(s_147), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1580(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1581(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1582(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1541(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1542(.a(gate55inter0), .b(s_142), .O(gate55inter1));
  and2  gate1543(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1544(.a(s_142), .O(gate55inter3));
  inv1  gate1545(.a(s_143), .O(gate55inter4));
  nand2 gate1546(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1547(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1548(.a(G15), .O(gate55inter7));
  inv1  gate1549(.a(G287), .O(gate55inter8));
  nand2 gate1550(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1551(.a(s_143), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1552(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1553(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1554(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1415(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1416(.a(gate57inter0), .b(s_124), .O(gate57inter1));
  and2  gate1417(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1418(.a(s_124), .O(gate57inter3));
  inv1  gate1419(.a(s_125), .O(gate57inter4));
  nand2 gate1420(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1421(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1422(.a(G17), .O(gate57inter7));
  inv1  gate1423(.a(G290), .O(gate57inter8));
  nand2 gate1424(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1425(.a(s_125), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1426(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1427(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1428(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate757(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate758(.a(gate58inter0), .b(s_30), .O(gate58inter1));
  and2  gate759(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate760(.a(s_30), .O(gate58inter3));
  inv1  gate761(.a(s_31), .O(gate58inter4));
  nand2 gate762(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate763(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate764(.a(G18), .O(gate58inter7));
  inv1  gate765(.a(G290), .O(gate58inter8));
  nand2 gate766(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate767(.a(s_31), .b(gate58inter3), .O(gate58inter10));
  nor2  gate768(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate769(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate770(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate897(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate898(.a(gate60inter0), .b(s_50), .O(gate60inter1));
  and2  gate899(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate900(.a(s_50), .O(gate60inter3));
  inv1  gate901(.a(s_51), .O(gate60inter4));
  nand2 gate902(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate903(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate904(.a(G20), .O(gate60inter7));
  inv1  gate905(.a(G293), .O(gate60inter8));
  nand2 gate906(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate907(.a(s_51), .b(gate60inter3), .O(gate60inter10));
  nor2  gate908(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate909(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate910(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate617(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate618(.a(gate69inter0), .b(s_10), .O(gate69inter1));
  and2  gate619(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate620(.a(s_10), .O(gate69inter3));
  inv1  gate621(.a(s_11), .O(gate69inter4));
  nand2 gate622(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate623(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate624(.a(G29), .O(gate69inter7));
  inv1  gate625(.a(G308), .O(gate69inter8));
  nand2 gate626(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate627(.a(s_11), .b(gate69inter3), .O(gate69inter10));
  nor2  gate628(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate629(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate630(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1107(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1108(.a(gate70inter0), .b(s_80), .O(gate70inter1));
  and2  gate1109(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1110(.a(s_80), .O(gate70inter3));
  inv1  gate1111(.a(s_81), .O(gate70inter4));
  nand2 gate1112(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1113(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1114(.a(G30), .O(gate70inter7));
  inv1  gate1115(.a(G308), .O(gate70inter8));
  nand2 gate1116(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1117(.a(s_81), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1118(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1119(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1120(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1247(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1248(.a(gate72inter0), .b(s_100), .O(gate72inter1));
  and2  gate1249(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1250(.a(s_100), .O(gate72inter3));
  inv1  gate1251(.a(s_101), .O(gate72inter4));
  nand2 gate1252(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1253(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1254(.a(G32), .O(gate72inter7));
  inv1  gate1255(.a(G311), .O(gate72inter8));
  nand2 gate1256(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1257(.a(s_101), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1258(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1259(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1260(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate967(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate968(.a(gate80inter0), .b(s_60), .O(gate80inter1));
  and2  gate969(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate970(.a(s_60), .O(gate80inter3));
  inv1  gate971(.a(s_61), .O(gate80inter4));
  nand2 gate972(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate973(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate974(.a(G14), .O(gate80inter7));
  inv1  gate975(.a(G323), .O(gate80inter8));
  nand2 gate976(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate977(.a(s_61), .b(gate80inter3), .O(gate80inter10));
  nor2  gate978(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate979(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate980(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate575(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate576(.a(gate81inter0), .b(s_4), .O(gate81inter1));
  and2  gate577(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate578(.a(s_4), .O(gate81inter3));
  inv1  gate579(.a(s_5), .O(gate81inter4));
  nand2 gate580(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate581(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate582(.a(G3), .O(gate81inter7));
  inv1  gate583(.a(G326), .O(gate81inter8));
  nand2 gate584(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate585(.a(s_5), .b(gate81inter3), .O(gate81inter10));
  nor2  gate586(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate587(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate588(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1527(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1528(.a(gate86inter0), .b(s_140), .O(gate86inter1));
  and2  gate1529(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1530(.a(s_140), .O(gate86inter3));
  inv1  gate1531(.a(s_141), .O(gate86inter4));
  nand2 gate1532(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1533(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1534(.a(G8), .O(gate86inter7));
  inv1  gate1535(.a(G332), .O(gate86inter8));
  nand2 gate1536(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1537(.a(s_141), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1538(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1539(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1540(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate743(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate744(.a(gate101inter0), .b(s_28), .O(gate101inter1));
  and2  gate745(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate746(.a(s_28), .O(gate101inter3));
  inv1  gate747(.a(s_29), .O(gate101inter4));
  nand2 gate748(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate749(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate750(.a(G20), .O(gate101inter7));
  inv1  gate751(.a(G356), .O(gate101inter8));
  nand2 gate752(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate753(.a(s_29), .b(gate101inter3), .O(gate101inter10));
  nor2  gate754(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate755(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate756(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate925(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate926(.a(gate105inter0), .b(s_54), .O(gate105inter1));
  and2  gate927(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate928(.a(s_54), .O(gate105inter3));
  inv1  gate929(.a(s_55), .O(gate105inter4));
  nand2 gate930(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate931(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate932(.a(G362), .O(gate105inter7));
  inv1  gate933(.a(G363), .O(gate105inter8));
  nand2 gate934(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate935(.a(s_55), .b(gate105inter3), .O(gate105inter10));
  nor2  gate936(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate937(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate938(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1261(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1262(.a(gate110inter0), .b(s_102), .O(gate110inter1));
  and2  gate1263(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1264(.a(s_102), .O(gate110inter3));
  inv1  gate1265(.a(s_103), .O(gate110inter4));
  nand2 gate1266(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1267(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1268(.a(G372), .O(gate110inter7));
  inv1  gate1269(.a(G373), .O(gate110inter8));
  nand2 gate1270(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1271(.a(s_103), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1272(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1273(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1274(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1429(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1430(.a(gate114inter0), .b(s_126), .O(gate114inter1));
  and2  gate1431(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1432(.a(s_126), .O(gate114inter3));
  inv1  gate1433(.a(s_127), .O(gate114inter4));
  nand2 gate1434(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1435(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1436(.a(G380), .O(gate114inter7));
  inv1  gate1437(.a(G381), .O(gate114inter8));
  nand2 gate1438(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1439(.a(s_127), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1440(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1441(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1442(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate673(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate674(.a(gate121inter0), .b(s_18), .O(gate121inter1));
  and2  gate675(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate676(.a(s_18), .O(gate121inter3));
  inv1  gate677(.a(s_19), .O(gate121inter4));
  nand2 gate678(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate679(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate680(.a(G394), .O(gate121inter7));
  inv1  gate681(.a(G395), .O(gate121inter8));
  nand2 gate682(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate683(.a(s_19), .b(gate121inter3), .O(gate121inter10));
  nor2  gate684(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate685(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate686(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1513(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1514(.a(gate126inter0), .b(s_138), .O(gate126inter1));
  and2  gate1515(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1516(.a(s_138), .O(gate126inter3));
  inv1  gate1517(.a(s_139), .O(gate126inter4));
  nand2 gate1518(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1519(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1520(.a(G404), .O(gate126inter7));
  inv1  gate1521(.a(G405), .O(gate126inter8));
  nand2 gate1522(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1523(.a(s_139), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1524(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1525(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1526(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate883(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate884(.a(gate129inter0), .b(s_48), .O(gate129inter1));
  and2  gate885(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate886(.a(s_48), .O(gate129inter3));
  inv1  gate887(.a(s_49), .O(gate129inter4));
  nand2 gate888(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate889(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate890(.a(G410), .O(gate129inter7));
  inv1  gate891(.a(G411), .O(gate129inter8));
  nand2 gate892(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate893(.a(s_49), .b(gate129inter3), .O(gate129inter10));
  nor2  gate894(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate895(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate896(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1289(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1290(.a(gate131inter0), .b(s_106), .O(gate131inter1));
  and2  gate1291(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1292(.a(s_106), .O(gate131inter3));
  inv1  gate1293(.a(s_107), .O(gate131inter4));
  nand2 gate1294(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1295(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1296(.a(G414), .O(gate131inter7));
  inv1  gate1297(.a(G415), .O(gate131inter8));
  nand2 gate1298(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1299(.a(s_107), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1300(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1301(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1302(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1709(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1710(.a(gate134inter0), .b(s_166), .O(gate134inter1));
  and2  gate1711(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1712(.a(s_166), .O(gate134inter3));
  inv1  gate1713(.a(s_167), .O(gate134inter4));
  nand2 gate1714(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1715(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1716(.a(G420), .O(gate134inter7));
  inv1  gate1717(.a(G421), .O(gate134inter8));
  nand2 gate1718(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1719(.a(s_167), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1720(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1721(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1722(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1401(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1402(.a(gate142inter0), .b(s_122), .O(gate142inter1));
  and2  gate1403(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1404(.a(s_122), .O(gate142inter3));
  inv1  gate1405(.a(s_123), .O(gate142inter4));
  nand2 gate1406(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1407(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1408(.a(G456), .O(gate142inter7));
  inv1  gate1409(.a(G459), .O(gate142inter8));
  nand2 gate1410(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1411(.a(s_123), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1412(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1413(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1414(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1149(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1150(.a(gate169inter0), .b(s_86), .O(gate169inter1));
  and2  gate1151(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1152(.a(s_86), .O(gate169inter3));
  inv1  gate1153(.a(s_87), .O(gate169inter4));
  nand2 gate1154(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1155(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1156(.a(G474), .O(gate169inter7));
  inv1  gate1157(.a(G546), .O(gate169inter8));
  nand2 gate1158(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1159(.a(s_87), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1160(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1161(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1162(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1205(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1206(.a(gate170inter0), .b(s_94), .O(gate170inter1));
  and2  gate1207(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1208(.a(s_94), .O(gate170inter3));
  inv1  gate1209(.a(s_95), .O(gate170inter4));
  nand2 gate1210(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1211(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1212(.a(G477), .O(gate170inter7));
  inv1  gate1213(.a(G546), .O(gate170inter8));
  nand2 gate1214(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1215(.a(s_95), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1216(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1217(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1218(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1163(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1164(.a(gate174inter0), .b(s_88), .O(gate174inter1));
  and2  gate1165(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1166(.a(s_88), .O(gate174inter3));
  inv1  gate1167(.a(s_89), .O(gate174inter4));
  nand2 gate1168(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1169(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1170(.a(G489), .O(gate174inter7));
  inv1  gate1171(.a(G552), .O(gate174inter8));
  nand2 gate1172(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1173(.a(s_89), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1174(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1175(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1176(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1499(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1500(.a(gate177inter0), .b(s_136), .O(gate177inter1));
  and2  gate1501(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1502(.a(s_136), .O(gate177inter3));
  inv1  gate1503(.a(s_137), .O(gate177inter4));
  nand2 gate1504(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1505(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1506(.a(G498), .O(gate177inter7));
  inv1  gate1507(.a(G558), .O(gate177inter8));
  nand2 gate1508(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1509(.a(s_137), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1510(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1511(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1512(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1331(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1332(.a(gate182inter0), .b(s_112), .O(gate182inter1));
  and2  gate1333(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1334(.a(s_112), .O(gate182inter3));
  inv1  gate1335(.a(s_113), .O(gate182inter4));
  nand2 gate1336(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1337(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1338(.a(G513), .O(gate182inter7));
  inv1  gate1339(.a(G564), .O(gate182inter8));
  nand2 gate1340(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1341(.a(s_113), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1342(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1343(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1344(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1485(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1486(.a(gate185inter0), .b(s_134), .O(gate185inter1));
  and2  gate1487(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1488(.a(s_134), .O(gate185inter3));
  inv1  gate1489(.a(s_135), .O(gate185inter4));
  nand2 gate1490(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1491(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1492(.a(G570), .O(gate185inter7));
  inv1  gate1493(.a(G571), .O(gate185inter8));
  nand2 gate1494(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1495(.a(s_135), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1496(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1497(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1498(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1387(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1388(.a(gate186inter0), .b(s_120), .O(gate186inter1));
  and2  gate1389(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1390(.a(s_120), .O(gate186inter3));
  inv1  gate1391(.a(s_121), .O(gate186inter4));
  nand2 gate1392(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1393(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1394(.a(G572), .O(gate186inter7));
  inv1  gate1395(.a(G573), .O(gate186inter8));
  nand2 gate1396(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1397(.a(s_121), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1398(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1399(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1400(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1093(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1094(.a(gate190inter0), .b(s_78), .O(gate190inter1));
  and2  gate1095(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1096(.a(s_78), .O(gate190inter3));
  inv1  gate1097(.a(s_79), .O(gate190inter4));
  nand2 gate1098(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1099(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1100(.a(G580), .O(gate190inter7));
  inv1  gate1101(.a(G581), .O(gate190inter8));
  nand2 gate1102(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1103(.a(s_79), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1104(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1105(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1106(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1345(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1346(.a(gate193inter0), .b(s_114), .O(gate193inter1));
  and2  gate1347(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1348(.a(s_114), .O(gate193inter3));
  inv1  gate1349(.a(s_115), .O(gate193inter4));
  nand2 gate1350(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1351(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1352(.a(G586), .O(gate193inter7));
  inv1  gate1353(.a(G587), .O(gate193inter8));
  nand2 gate1354(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1355(.a(s_115), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1356(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1357(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1358(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate729(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate730(.a(gate194inter0), .b(s_26), .O(gate194inter1));
  and2  gate731(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate732(.a(s_26), .O(gate194inter3));
  inv1  gate733(.a(s_27), .O(gate194inter4));
  nand2 gate734(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate735(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate736(.a(G588), .O(gate194inter7));
  inv1  gate737(.a(G589), .O(gate194inter8));
  nand2 gate738(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate739(.a(s_27), .b(gate194inter3), .O(gate194inter10));
  nor2  gate740(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate741(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate742(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1135(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1136(.a(gate195inter0), .b(s_84), .O(gate195inter1));
  and2  gate1137(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1138(.a(s_84), .O(gate195inter3));
  inv1  gate1139(.a(s_85), .O(gate195inter4));
  nand2 gate1140(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1141(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1142(.a(G590), .O(gate195inter7));
  inv1  gate1143(.a(G591), .O(gate195inter8));
  nand2 gate1144(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1145(.a(s_85), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1146(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1147(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1148(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1051(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1052(.a(gate196inter0), .b(s_72), .O(gate196inter1));
  and2  gate1053(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1054(.a(s_72), .O(gate196inter3));
  inv1  gate1055(.a(s_73), .O(gate196inter4));
  nand2 gate1056(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1057(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1058(.a(G592), .O(gate196inter7));
  inv1  gate1059(.a(G593), .O(gate196inter8));
  nand2 gate1060(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1061(.a(s_73), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1062(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1063(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1064(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate827(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate828(.a(gate202inter0), .b(s_40), .O(gate202inter1));
  and2  gate829(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate830(.a(s_40), .O(gate202inter3));
  inv1  gate831(.a(s_41), .O(gate202inter4));
  nand2 gate832(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate833(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate834(.a(G612), .O(gate202inter7));
  inv1  gate835(.a(G617), .O(gate202inter8));
  nand2 gate836(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate837(.a(s_41), .b(gate202inter3), .O(gate202inter10));
  nor2  gate838(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate839(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate840(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate547(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate548(.a(gate212inter0), .b(s_0), .O(gate212inter1));
  and2  gate549(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate550(.a(s_0), .O(gate212inter3));
  inv1  gate551(.a(s_1), .O(gate212inter4));
  nand2 gate552(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate553(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate554(.a(G617), .O(gate212inter7));
  inv1  gate555(.a(G669), .O(gate212inter8));
  nand2 gate556(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate557(.a(s_1), .b(gate212inter3), .O(gate212inter10));
  nor2  gate558(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate559(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate560(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1121(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1122(.a(gate216inter0), .b(s_82), .O(gate216inter1));
  and2  gate1123(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1124(.a(s_82), .O(gate216inter3));
  inv1  gate1125(.a(s_83), .O(gate216inter4));
  nand2 gate1126(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1127(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1128(.a(G617), .O(gate216inter7));
  inv1  gate1129(.a(G675), .O(gate216inter8));
  nand2 gate1130(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1131(.a(s_83), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1132(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1133(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1134(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate869(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate870(.a(gate234inter0), .b(s_46), .O(gate234inter1));
  and2  gate871(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate872(.a(s_46), .O(gate234inter3));
  inv1  gate873(.a(s_47), .O(gate234inter4));
  nand2 gate874(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate875(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate876(.a(G245), .O(gate234inter7));
  inv1  gate877(.a(G721), .O(gate234inter8));
  nand2 gate878(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate879(.a(s_47), .b(gate234inter3), .O(gate234inter10));
  nor2  gate880(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate881(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate882(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1723(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1724(.a(gate237inter0), .b(s_168), .O(gate237inter1));
  and2  gate1725(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1726(.a(s_168), .O(gate237inter3));
  inv1  gate1727(.a(s_169), .O(gate237inter4));
  nand2 gate1728(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1729(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1730(.a(G254), .O(gate237inter7));
  inv1  gate1731(.a(G706), .O(gate237inter8));
  nand2 gate1732(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1733(.a(s_169), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1734(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1735(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1736(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1639(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1640(.a(gate242inter0), .b(s_156), .O(gate242inter1));
  and2  gate1641(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1642(.a(s_156), .O(gate242inter3));
  inv1  gate1643(.a(s_157), .O(gate242inter4));
  nand2 gate1644(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1645(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1646(.a(G718), .O(gate242inter7));
  inv1  gate1647(.a(G730), .O(gate242inter8));
  nand2 gate1648(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1649(.a(s_157), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1650(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1651(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1652(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate939(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate940(.a(gate250inter0), .b(s_56), .O(gate250inter1));
  and2  gate941(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate942(.a(s_56), .O(gate250inter3));
  inv1  gate943(.a(s_57), .O(gate250inter4));
  nand2 gate944(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate945(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate946(.a(G706), .O(gate250inter7));
  inv1  gate947(.a(G742), .O(gate250inter8));
  nand2 gate948(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate949(.a(s_57), .b(gate250inter3), .O(gate250inter10));
  nor2  gate950(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate951(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate952(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate995(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate996(.a(gate252inter0), .b(s_64), .O(gate252inter1));
  and2  gate997(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate998(.a(s_64), .O(gate252inter3));
  inv1  gate999(.a(s_65), .O(gate252inter4));
  nand2 gate1000(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1001(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1002(.a(G709), .O(gate252inter7));
  inv1  gate1003(.a(G745), .O(gate252inter8));
  nand2 gate1004(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1005(.a(s_65), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1006(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1007(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1008(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1625(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1626(.a(gate256inter0), .b(s_154), .O(gate256inter1));
  and2  gate1627(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1628(.a(s_154), .O(gate256inter3));
  inv1  gate1629(.a(s_155), .O(gate256inter4));
  nand2 gate1630(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1631(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1632(.a(G715), .O(gate256inter7));
  inv1  gate1633(.a(G751), .O(gate256inter8));
  nand2 gate1634(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1635(.a(s_155), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1636(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1637(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1638(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate911(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate912(.a(gate257inter0), .b(s_52), .O(gate257inter1));
  and2  gate913(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate914(.a(s_52), .O(gate257inter3));
  inv1  gate915(.a(s_53), .O(gate257inter4));
  nand2 gate916(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate917(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate918(.a(G754), .O(gate257inter7));
  inv1  gate919(.a(G755), .O(gate257inter8));
  nand2 gate920(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate921(.a(s_53), .b(gate257inter3), .O(gate257inter10));
  nor2  gate922(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate923(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate924(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate813(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate814(.a(gate268inter0), .b(s_38), .O(gate268inter1));
  and2  gate815(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate816(.a(s_38), .O(gate268inter3));
  inv1  gate817(.a(s_39), .O(gate268inter4));
  nand2 gate818(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate819(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate820(.a(G651), .O(gate268inter7));
  inv1  gate821(.a(G779), .O(gate268inter8));
  nand2 gate822(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate823(.a(s_39), .b(gate268inter3), .O(gate268inter10));
  nor2  gate824(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate825(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate826(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1065(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1066(.a(gate276inter0), .b(s_74), .O(gate276inter1));
  and2  gate1067(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1068(.a(s_74), .O(gate276inter3));
  inv1  gate1069(.a(s_75), .O(gate276inter4));
  nand2 gate1070(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1071(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1072(.a(G773), .O(gate276inter7));
  inv1  gate1073(.a(G797), .O(gate276inter8));
  nand2 gate1074(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1075(.a(s_75), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1076(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1077(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1078(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate589(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate590(.a(gate387inter0), .b(s_6), .O(gate387inter1));
  and2  gate591(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate592(.a(s_6), .O(gate387inter3));
  inv1  gate593(.a(s_7), .O(gate387inter4));
  nand2 gate594(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate595(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate596(.a(G1), .O(gate387inter7));
  inv1  gate597(.a(G1036), .O(gate387inter8));
  nand2 gate598(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate599(.a(s_7), .b(gate387inter3), .O(gate387inter10));
  nor2  gate600(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate601(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate602(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1023(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1024(.a(gate388inter0), .b(s_68), .O(gate388inter1));
  and2  gate1025(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1026(.a(s_68), .O(gate388inter3));
  inv1  gate1027(.a(s_69), .O(gate388inter4));
  nand2 gate1028(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1029(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1030(.a(G2), .O(gate388inter7));
  inv1  gate1031(.a(G1039), .O(gate388inter8));
  nand2 gate1032(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1033(.a(s_69), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1034(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1035(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1036(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate603(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate604(.a(gate390inter0), .b(s_8), .O(gate390inter1));
  and2  gate605(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate606(.a(s_8), .O(gate390inter3));
  inv1  gate607(.a(s_9), .O(gate390inter4));
  nand2 gate608(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate609(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate610(.a(G4), .O(gate390inter7));
  inv1  gate611(.a(G1045), .O(gate390inter8));
  nand2 gate612(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate613(.a(s_9), .b(gate390inter3), .O(gate390inter10));
  nor2  gate614(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate615(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate616(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1009(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1010(.a(gate398inter0), .b(s_66), .O(gate398inter1));
  and2  gate1011(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1012(.a(s_66), .O(gate398inter3));
  inv1  gate1013(.a(s_67), .O(gate398inter4));
  nand2 gate1014(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1015(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1016(.a(G12), .O(gate398inter7));
  inv1  gate1017(.a(G1069), .O(gate398inter8));
  nand2 gate1018(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1019(.a(s_67), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1020(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1021(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1022(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1079(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1080(.a(gate399inter0), .b(s_76), .O(gate399inter1));
  and2  gate1081(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1082(.a(s_76), .O(gate399inter3));
  inv1  gate1083(.a(s_77), .O(gate399inter4));
  nand2 gate1084(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1085(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1086(.a(G13), .O(gate399inter7));
  inv1  gate1087(.a(G1072), .O(gate399inter8));
  nand2 gate1088(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1089(.a(s_77), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1090(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1091(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1092(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1555(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1556(.a(gate400inter0), .b(s_144), .O(gate400inter1));
  and2  gate1557(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1558(.a(s_144), .O(gate400inter3));
  inv1  gate1559(.a(s_145), .O(gate400inter4));
  nand2 gate1560(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1561(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1562(.a(G14), .O(gate400inter7));
  inv1  gate1563(.a(G1075), .O(gate400inter8));
  nand2 gate1564(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1565(.a(s_145), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1566(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1567(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1568(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1303(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1304(.a(gate401inter0), .b(s_108), .O(gate401inter1));
  and2  gate1305(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1306(.a(s_108), .O(gate401inter3));
  inv1  gate1307(.a(s_109), .O(gate401inter4));
  nand2 gate1308(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1309(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1310(.a(G15), .O(gate401inter7));
  inv1  gate1311(.a(G1078), .O(gate401inter8));
  nand2 gate1312(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1313(.a(s_109), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1314(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1315(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1316(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate645(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate646(.a(gate406inter0), .b(s_14), .O(gate406inter1));
  and2  gate647(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate648(.a(s_14), .O(gate406inter3));
  inv1  gate649(.a(s_15), .O(gate406inter4));
  nand2 gate650(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate651(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate652(.a(G20), .O(gate406inter7));
  inv1  gate653(.a(G1093), .O(gate406inter8));
  nand2 gate654(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate655(.a(s_15), .b(gate406inter3), .O(gate406inter10));
  nor2  gate656(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate657(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate658(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate687(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate688(.a(gate409inter0), .b(s_20), .O(gate409inter1));
  and2  gate689(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate690(.a(s_20), .O(gate409inter3));
  inv1  gate691(.a(s_21), .O(gate409inter4));
  nand2 gate692(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate693(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate694(.a(G23), .O(gate409inter7));
  inv1  gate695(.a(G1102), .O(gate409inter8));
  nand2 gate696(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate697(.a(s_21), .b(gate409inter3), .O(gate409inter10));
  nor2  gate698(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate699(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate700(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1583(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1584(.a(gate412inter0), .b(s_148), .O(gate412inter1));
  and2  gate1585(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1586(.a(s_148), .O(gate412inter3));
  inv1  gate1587(.a(s_149), .O(gate412inter4));
  nand2 gate1588(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1589(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1590(.a(G26), .O(gate412inter7));
  inv1  gate1591(.a(G1111), .O(gate412inter8));
  nand2 gate1592(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1593(.a(s_149), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1594(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1595(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1596(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1373(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1374(.a(gate417inter0), .b(s_118), .O(gate417inter1));
  and2  gate1375(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1376(.a(s_118), .O(gate417inter3));
  inv1  gate1377(.a(s_119), .O(gate417inter4));
  nand2 gate1378(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1379(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1380(.a(G31), .O(gate417inter7));
  inv1  gate1381(.a(G1126), .O(gate417inter8));
  nand2 gate1382(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1383(.a(s_119), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1384(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1385(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1386(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1737(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1738(.a(gate418inter0), .b(s_170), .O(gate418inter1));
  and2  gate1739(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1740(.a(s_170), .O(gate418inter3));
  inv1  gate1741(.a(s_171), .O(gate418inter4));
  nand2 gate1742(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1743(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1744(.a(G32), .O(gate418inter7));
  inv1  gate1745(.a(G1129), .O(gate418inter8));
  nand2 gate1746(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1747(.a(s_171), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1748(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1749(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1750(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1191(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1192(.a(gate427inter0), .b(s_92), .O(gate427inter1));
  and2  gate1193(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1194(.a(s_92), .O(gate427inter3));
  inv1  gate1195(.a(s_93), .O(gate427inter4));
  nand2 gate1196(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1197(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1198(.a(G5), .O(gate427inter7));
  inv1  gate1199(.a(G1144), .O(gate427inter8));
  nand2 gate1200(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1201(.a(s_93), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1202(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1203(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1204(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1681(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1682(.a(gate429inter0), .b(s_162), .O(gate429inter1));
  and2  gate1683(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1684(.a(s_162), .O(gate429inter3));
  inv1  gate1685(.a(s_163), .O(gate429inter4));
  nand2 gate1686(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1687(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1688(.a(G6), .O(gate429inter7));
  inv1  gate1689(.a(G1147), .O(gate429inter8));
  nand2 gate1690(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1691(.a(s_163), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1692(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1693(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1694(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate659(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate660(.a(gate441inter0), .b(s_16), .O(gate441inter1));
  and2  gate661(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate662(.a(s_16), .O(gate441inter3));
  inv1  gate663(.a(s_17), .O(gate441inter4));
  nand2 gate664(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate665(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate666(.a(G12), .O(gate441inter7));
  inv1  gate667(.a(G1165), .O(gate441inter8));
  nand2 gate668(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate669(.a(s_17), .b(gate441inter3), .O(gate441inter10));
  nor2  gate670(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate671(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate672(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1695(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1696(.a(gate444inter0), .b(s_164), .O(gate444inter1));
  and2  gate1697(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1698(.a(s_164), .O(gate444inter3));
  inv1  gate1699(.a(s_165), .O(gate444inter4));
  nand2 gate1700(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1701(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1702(.a(G1072), .O(gate444inter7));
  inv1  gate1703(.a(G1168), .O(gate444inter8));
  nand2 gate1704(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1705(.a(s_165), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1706(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1707(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1708(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1443(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1444(.a(gate447inter0), .b(s_128), .O(gate447inter1));
  and2  gate1445(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1446(.a(s_128), .O(gate447inter3));
  inv1  gate1447(.a(s_129), .O(gate447inter4));
  nand2 gate1448(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1449(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1450(.a(G15), .O(gate447inter7));
  inv1  gate1451(.a(G1174), .O(gate447inter8));
  nand2 gate1452(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1453(.a(s_129), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1454(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1455(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1456(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate953(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate954(.a(gate450inter0), .b(s_58), .O(gate450inter1));
  and2  gate955(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate956(.a(s_58), .O(gate450inter3));
  inv1  gate957(.a(s_59), .O(gate450inter4));
  nand2 gate958(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate959(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate960(.a(G1081), .O(gate450inter7));
  inv1  gate961(.a(G1177), .O(gate450inter8));
  nand2 gate962(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate963(.a(s_59), .b(gate450inter3), .O(gate450inter10));
  nor2  gate964(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate965(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate966(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1471(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1472(.a(gate452inter0), .b(s_132), .O(gate452inter1));
  and2  gate1473(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1474(.a(s_132), .O(gate452inter3));
  inv1  gate1475(.a(s_133), .O(gate452inter4));
  nand2 gate1476(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1477(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1478(.a(G1084), .O(gate452inter7));
  inv1  gate1479(.a(G1180), .O(gate452inter8));
  nand2 gate1480(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1481(.a(s_133), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1482(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1483(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1484(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1317(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1318(.a(gate454inter0), .b(s_110), .O(gate454inter1));
  and2  gate1319(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1320(.a(s_110), .O(gate454inter3));
  inv1  gate1321(.a(s_111), .O(gate454inter4));
  nand2 gate1322(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1323(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1324(.a(G1087), .O(gate454inter7));
  inv1  gate1325(.a(G1183), .O(gate454inter8));
  nand2 gate1326(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1327(.a(s_111), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1328(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1329(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1330(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1457(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1458(.a(gate455inter0), .b(s_130), .O(gate455inter1));
  and2  gate1459(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1460(.a(s_130), .O(gate455inter3));
  inv1  gate1461(.a(s_131), .O(gate455inter4));
  nand2 gate1462(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1463(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1464(.a(G19), .O(gate455inter7));
  inv1  gate1465(.a(G1186), .O(gate455inter8));
  nand2 gate1466(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1467(.a(s_131), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1468(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1469(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1470(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1233(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1234(.a(gate462inter0), .b(s_98), .O(gate462inter1));
  and2  gate1235(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1236(.a(s_98), .O(gate462inter3));
  inv1  gate1237(.a(s_99), .O(gate462inter4));
  nand2 gate1238(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1239(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1240(.a(G1099), .O(gate462inter7));
  inv1  gate1241(.a(G1195), .O(gate462inter8));
  nand2 gate1242(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1243(.a(s_99), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1244(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1245(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1246(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate785(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate786(.a(gate466inter0), .b(s_34), .O(gate466inter1));
  and2  gate787(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate788(.a(s_34), .O(gate466inter3));
  inv1  gate789(.a(s_35), .O(gate466inter4));
  nand2 gate790(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate791(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate792(.a(G1105), .O(gate466inter7));
  inv1  gate793(.a(G1201), .O(gate466inter8));
  nand2 gate794(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate795(.a(s_35), .b(gate466inter3), .O(gate466inter10));
  nor2  gate796(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate797(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate798(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1037(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1038(.a(gate470inter0), .b(s_70), .O(gate470inter1));
  and2  gate1039(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1040(.a(s_70), .O(gate470inter3));
  inv1  gate1041(.a(s_71), .O(gate470inter4));
  nand2 gate1042(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1043(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1044(.a(G1111), .O(gate470inter7));
  inv1  gate1045(.a(G1207), .O(gate470inter8));
  nand2 gate1046(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1047(.a(s_71), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1048(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1049(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1050(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate715(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate716(.a(gate471inter0), .b(s_24), .O(gate471inter1));
  and2  gate717(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate718(.a(s_24), .O(gate471inter3));
  inv1  gate719(.a(s_25), .O(gate471inter4));
  nand2 gate720(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate721(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate722(.a(G27), .O(gate471inter7));
  inv1  gate723(.a(G1210), .O(gate471inter8));
  nand2 gate724(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate725(.a(s_25), .b(gate471inter3), .O(gate471inter10));
  nor2  gate726(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate727(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate728(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate631(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate632(.a(gate477inter0), .b(s_12), .O(gate477inter1));
  and2  gate633(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate634(.a(s_12), .O(gate477inter3));
  inv1  gate635(.a(s_13), .O(gate477inter4));
  nand2 gate636(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate637(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate638(.a(G30), .O(gate477inter7));
  inv1  gate639(.a(G1219), .O(gate477inter8));
  nand2 gate640(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate641(.a(s_13), .b(gate477inter3), .O(gate477inter10));
  nor2  gate642(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate643(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate644(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1177(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1178(.a(gate481inter0), .b(s_90), .O(gate481inter1));
  and2  gate1179(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1180(.a(s_90), .O(gate481inter3));
  inv1  gate1181(.a(s_91), .O(gate481inter4));
  nand2 gate1182(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1183(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1184(.a(G32), .O(gate481inter7));
  inv1  gate1185(.a(G1225), .O(gate481inter8));
  nand2 gate1186(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1187(.a(s_91), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1188(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1189(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1190(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1359(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1360(.a(gate484inter0), .b(s_116), .O(gate484inter1));
  and2  gate1361(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1362(.a(s_116), .O(gate484inter3));
  inv1  gate1363(.a(s_117), .O(gate484inter4));
  nand2 gate1364(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1365(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1366(.a(G1230), .O(gate484inter7));
  inv1  gate1367(.a(G1231), .O(gate484inter8));
  nand2 gate1368(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1369(.a(s_117), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1370(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1371(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1372(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate799(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate800(.a(gate485inter0), .b(s_36), .O(gate485inter1));
  and2  gate801(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate802(.a(s_36), .O(gate485inter3));
  inv1  gate803(.a(s_37), .O(gate485inter4));
  nand2 gate804(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate805(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate806(.a(G1232), .O(gate485inter7));
  inv1  gate807(.a(G1233), .O(gate485inter8));
  nand2 gate808(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate809(.a(s_37), .b(gate485inter3), .O(gate485inter10));
  nor2  gate810(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate811(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate812(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1219(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1220(.a(gate491inter0), .b(s_96), .O(gate491inter1));
  and2  gate1221(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1222(.a(s_96), .O(gate491inter3));
  inv1  gate1223(.a(s_97), .O(gate491inter4));
  nand2 gate1224(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1225(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1226(.a(G1244), .O(gate491inter7));
  inv1  gate1227(.a(G1245), .O(gate491inter8));
  nand2 gate1228(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1229(.a(s_97), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1230(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1231(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1232(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate771(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate772(.a(gate507inter0), .b(s_32), .O(gate507inter1));
  and2  gate773(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate774(.a(s_32), .O(gate507inter3));
  inv1  gate775(.a(s_33), .O(gate507inter4));
  nand2 gate776(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate777(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate778(.a(G1276), .O(gate507inter7));
  inv1  gate779(.a(G1277), .O(gate507inter8));
  nand2 gate780(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate781(.a(s_33), .b(gate507inter3), .O(gate507inter10));
  nor2  gate782(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate783(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate784(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule