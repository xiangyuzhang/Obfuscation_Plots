module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2367(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2368(.a(gate15inter0), .b(s_260), .O(gate15inter1));
  and2  gate2369(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2370(.a(s_260), .O(gate15inter3));
  inv1  gate2371(.a(s_261), .O(gate15inter4));
  nand2 gate2372(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2373(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2374(.a(G13), .O(gate15inter7));
  inv1  gate2375(.a(G14), .O(gate15inter8));
  nand2 gate2376(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2377(.a(s_261), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2378(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2379(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2380(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1415(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1416(.a(gate19inter0), .b(s_124), .O(gate19inter1));
  and2  gate1417(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1418(.a(s_124), .O(gate19inter3));
  inv1  gate1419(.a(s_125), .O(gate19inter4));
  nand2 gate1420(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1421(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1422(.a(G21), .O(gate19inter7));
  inv1  gate1423(.a(G22), .O(gate19inter8));
  nand2 gate1424(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1425(.a(s_125), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1426(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1427(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1428(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1975(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1976(.a(gate21inter0), .b(s_204), .O(gate21inter1));
  and2  gate1977(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1978(.a(s_204), .O(gate21inter3));
  inv1  gate1979(.a(s_205), .O(gate21inter4));
  nand2 gate1980(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1981(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1982(.a(G25), .O(gate21inter7));
  inv1  gate1983(.a(G26), .O(gate21inter8));
  nand2 gate1984(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1985(.a(s_205), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1986(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1987(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1988(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2227(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2228(.a(gate23inter0), .b(s_240), .O(gate23inter1));
  and2  gate2229(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2230(.a(s_240), .O(gate23inter3));
  inv1  gate2231(.a(s_241), .O(gate23inter4));
  nand2 gate2232(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2233(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2234(.a(G29), .O(gate23inter7));
  inv1  gate2235(.a(G30), .O(gate23inter8));
  nand2 gate2236(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2237(.a(s_241), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2238(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2239(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2240(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate869(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate870(.a(gate24inter0), .b(s_46), .O(gate24inter1));
  and2  gate871(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate872(.a(s_46), .O(gate24inter3));
  inv1  gate873(.a(s_47), .O(gate24inter4));
  nand2 gate874(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate875(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate876(.a(G31), .O(gate24inter7));
  inv1  gate877(.a(G32), .O(gate24inter8));
  nand2 gate878(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate879(.a(s_47), .b(gate24inter3), .O(gate24inter10));
  nor2  gate880(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate881(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate882(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate2647(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2648(.a(gate25inter0), .b(s_300), .O(gate25inter1));
  and2  gate2649(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2650(.a(s_300), .O(gate25inter3));
  inv1  gate2651(.a(s_301), .O(gate25inter4));
  nand2 gate2652(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2653(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2654(.a(G1), .O(gate25inter7));
  inv1  gate2655(.a(G5), .O(gate25inter8));
  nand2 gate2656(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2657(.a(s_301), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2658(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2659(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2660(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1709(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1710(.a(gate26inter0), .b(s_166), .O(gate26inter1));
  and2  gate1711(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1712(.a(s_166), .O(gate26inter3));
  inv1  gate1713(.a(s_167), .O(gate26inter4));
  nand2 gate1714(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1715(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1716(.a(G9), .O(gate26inter7));
  inv1  gate1717(.a(G13), .O(gate26inter8));
  nand2 gate1718(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1719(.a(s_167), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1720(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1721(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1722(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2997(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2998(.a(gate28inter0), .b(s_350), .O(gate28inter1));
  and2  gate2999(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate3000(.a(s_350), .O(gate28inter3));
  inv1  gate3001(.a(s_351), .O(gate28inter4));
  nand2 gate3002(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate3003(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate3004(.a(G10), .O(gate28inter7));
  inv1  gate3005(.a(G14), .O(gate28inter8));
  nand2 gate3006(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate3007(.a(s_351), .b(gate28inter3), .O(gate28inter10));
  nor2  gate3008(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate3009(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate3010(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate911(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate912(.a(gate33inter0), .b(s_52), .O(gate33inter1));
  and2  gate913(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate914(.a(s_52), .O(gate33inter3));
  inv1  gate915(.a(s_53), .O(gate33inter4));
  nand2 gate916(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate917(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate918(.a(G17), .O(gate33inter7));
  inv1  gate919(.a(G21), .O(gate33inter8));
  nand2 gate920(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate921(.a(s_53), .b(gate33inter3), .O(gate33inter10));
  nor2  gate922(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate923(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate924(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2115(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2116(.a(gate34inter0), .b(s_224), .O(gate34inter1));
  and2  gate2117(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2118(.a(s_224), .O(gate34inter3));
  inv1  gate2119(.a(s_225), .O(gate34inter4));
  nand2 gate2120(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2121(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2122(.a(G25), .O(gate34inter7));
  inv1  gate2123(.a(G29), .O(gate34inter8));
  nand2 gate2124(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2125(.a(s_225), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2126(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2127(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2128(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate659(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate660(.a(gate35inter0), .b(s_16), .O(gate35inter1));
  and2  gate661(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate662(.a(s_16), .O(gate35inter3));
  inv1  gate663(.a(s_17), .O(gate35inter4));
  nand2 gate664(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate665(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate666(.a(G18), .O(gate35inter7));
  inv1  gate667(.a(G22), .O(gate35inter8));
  nand2 gate668(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate669(.a(s_17), .b(gate35inter3), .O(gate35inter10));
  nor2  gate670(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate671(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate672(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1723(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1724(.a(gate38inter0), .b(s_168), .O(gate38inter1));
  and2  gate1725(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1726(.a(s_168), .O(gate38inter3));
  inv1  gate1727(.a(s_169), .O(gate38inter4));
  nand2 gate1728(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1729(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1730(.a(G27), .O(gate38inter7));
  inv1  gate1731(.a(G31), .O(gate38inter8));
  nand2 gate1732(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1733(.a(s_169), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1734(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1735(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1736(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1149(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1150(.a(gate40inter0), .b(s_86), .O(gate40inter1));
  and2  gate1151(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1152(.a(s_86), .O(gate40inter3));
  inv1  gate1153(.a(s_87), .O(gate40inter4));
  nand2 gate1154(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1155(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1156(.a(G28), .O(gate40inter7));
  inv1  gate1157(.a(G32), .O(gate40inter8));
  nand2 gate1158(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1159(.a(s_87), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1160(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1161(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1162(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2493(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2494(.a(gate41inter0), .b(s_278), .O(gate41inter1));
  and2  gate2495(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2496(.a(s_278), .O(gate41inter3));
  inv1  gate2497(.a(s_279), .O(gate41inter4));
  nand2 gate2498(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2499(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2500(.a(G1), .O(gate41inter7));
  inv1  gate2501(.a(G266), .O(gate41inter8));
  nand2 gate2502(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2503(.a(s_279), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2504(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2505(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2506(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2031(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2032(.a(gate46inter0), .b(s_212), .O(gate46inter1));
  and2  gate2033(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2034(.a(s_212), .O(gate46inter3));
  inv1  gate2035(.a(s_213), .O(gate46inter4));
  nand2 gate2036(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2037(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2038(.a(G6), .O(gate46inter7));
  inv1  gate2039(.a(G272), .O(gate46inter8));
  nand2 gate2040(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2041(.a(s_213), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2042(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2043(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2044(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2759(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2760(.a(gate49inter0), .b(s_316), .O(gate49inter1));
  and2  gate2761(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2762(.a(s_316), .O(gate49inter3));
  inv1  gate2763(.a(s_317), .O(gate49inter4));
  nand2 gate2764(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2765(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2766(.a(G9), .O(gate49inter7));
  inv1  gate2767(.a(G278), .O(gate49inter8));
  nand2 gate2768(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2769(.a(s_317), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2770(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2771(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2772(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1219(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1220(.a(gate50inter0), .b(s_96), .O(gate50inter1));
  and2  gate1221(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1222(.a(s_96), .O(gate50inter3));
  inv1  gate1223(.a(s_97), .O(gate50inter4));
  nand2 gate1224(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1225(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1226(.a(G10), .O(gate50inter7));
  inv1  gate1227(.a(G278), .O(gate50inter8));
  nand2 gate1228(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1229(.a(s_97), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1230(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1231(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1232(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2269(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2270(.a(gate51inter0), .b(s_246), .O(gate51inter1));
  and2  gate2271(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2272(.a(s_246), .O(gate51inter3));
  inv1  gate2273(.a(s_247), .O(gate51inter4));
  nand2 gate2274(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2275(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2276(.a(G11), .O(gate51inter7));
  inv1  gate2277(.a(G281), .O(gate51inter8));
  nand2 gate2278(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2279(.a(s_247), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2280(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2281(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2282(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1079(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1080(.a(gate55inter0), .b(s_76), .O(gate55inter1));
  and2  gate1081(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1082(.a(s_76), .O(gate55inter3));
  inv1  gate1083(.a(s_77), .O(gate55inter4));
  nand2 gate1084(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1085(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1086(.a(G15), .O(gate55inter7));
  inv1  gate1087(.a(G287), .O(gate55inter8));
  nand2 gate1088(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1089(.a(s_77), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1090(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1091(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1092(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate953(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate954(.a(gate58inter0), .b(s_58), .O(gate58inter1));
  and2  gate955(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate956(.a(s_58), .O(gate58inter3));
  inv1  gate957(.a(s_59), .O(gate58inter4));
  nand2 gate958(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate959(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate960(.a(G18), .O(gate58inter7));
  inv1  gate961(.a(G290), .O(gate58inter8));
  nand2 gate962(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate963(.a(s_59), .b(gate58inter3), .O(gate58inter10));
  nor2  gate964(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate965(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate966(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2507(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2508(.a(gate62inter0), .b(s_280), .O(gate62inter1));
  and2  gate2509(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2510(.a(s_280), .O(gate62inter3));
  inv1  gate2511(.a(s_281), .O(gate62inter4));
  nand2 gate2512(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2513(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2514(.a(G22), .O(gate62inter7));
  inv1  gate2515(.a(G296), .O(gate62inter8));
  nand2 gate2516(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2517(.a(s_281), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2518(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2519(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2520(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate925(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate926(.a(gate64inter0), .b(s_54), .O(gate64inter1));
  and2  gate927(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate928(.a(s_54), .O(gate64inter3));
  inv1  gate929(.a(s_55), .O(gate64inter4));
  nand2 gate930(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate931(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate932(.a(G24), .O(gate64inter7));
  inv1  gate933(.a(G299), .O(gate64inter8));
  nand2 gate934(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate935(.a(s_55), .b(gate64inter3), .O(gate64inter10));
  nor2  gate936(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate937(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate938(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate2857(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2858(.a(gate65inter0), .b(s_330), .O(gate65inter1));
  and2  gate2859(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2860(.a(s_330), .O(gate65inter3));
  inv1  gate2861(.a(s_331), .O(gate65inter4));
  nand2 gate2862(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2863(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2864(.a(G25), .O(gate65inter7));
  inv1  gate2865(.a(G302), .O(gate65inter8));
  nand2 gate2866(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2867(.a(s_331), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2868(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2869(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2870(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1569(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1570(.a(gate66inter0), .b(s_146), .O(gate66inter1));
  and2  gate1571(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1572(.a(s_146), .O(gate66inter3));
  inv1  gate1573(.a(s_147), .O(gate66inter4));
  nand2 gate1574(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1575(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1576(.a(G26), .O(gate66inter7));
  inv1  gate1577(.a(G302), .O(gate66inter8));
  nand2 gate1578(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1579(.a(s_147), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1580(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1581(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1582(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1905(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1906(.a(gate67inter0), .b(s_194), .O(gate67inter1));
  and2  gate1907(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1908(.a(s_194), .O(gate67inter3));
  inv1  gate1909(.a(s_195), .O(gate67inter4));
  nand2 gate1910(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1911(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1912(.a(G27), .O(gate67inter7));
  inv1  gate1913(.a(G305), .O(gate67inter8));
  nand2 gate1914(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1915(.a(s_195), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1916(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1917(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1918(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate2409(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2410(.a(gate68inter0), .b(s_266), .O(gate68inter1));
  and2  gate2411(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2412(.a(s_266), .O(gate68inter3));
  inv1  gate2413(.a(s_267), .O(gate68inter4));
  nand2 gate2414(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2415(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2416(.a(G28), .O(gate68inter7));
  inv1  gate2417(.a(G305), .O(gate68inter8));
  nand2 gate2418(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2419(.a(s_267), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2420(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2421(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2422(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2087(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2088(.a(gate72inter0), .b(s_220), .O(gate72inter1));
  and2  gate2089(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2090(.a(s_220), .O(gate72inter3));
  inv1  gate2091(.a(s_221), .O(gate72inter4));
  nand2 gate2092(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2093(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2094(.a(G32), .O(gate72inter7));
  inv1  gate2095(.a(G311), .O(gate72inter8));
  nand2 gate2096(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2097(.a(s_221), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2098(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2099(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2100(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1317(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1318(.a(gate73inter0), .b(s_110), .O(gate73inter1));
  and2  gate1319(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1320(.a(s_110), .O(gate73inter3));
  inv1  gate1321(.a(s_111), .O(gate73inter4));
  nand2 gate1322(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1323(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1324(.a(G1), .O(gate73inter7));
  inv1  gate1325(.a(G314), .O(gate73inter8));
  nand2 gate1326(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1327(.a(s_111), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1328(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1329(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1330(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2003(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2004(.a(gate74inter0), .b(s_208), .O(gate74inter1));
  and2  gate2005(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2006(.a(s_208), .O(gate74inter3));
  inv1  gate2007(.a(s_209), .O(gate74inter4));
  nand2 gate2008(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2009(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2010(.a(G5), .O(gate74inter7));
  inv1  gate2011(.a(G314), .O(gate74inter8));
  nand2 gate2012(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2013(.a(s_209), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2014(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2015(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2016(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2871(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2872(.a(gate77inter0), .b(s_332), .O(gate77inter1));
  and2  gate2873(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2874(.a(s_332), .O(gate77inter3));
  inv1  gate2875(.a(s_333), .O(gate77inter4));
  nand2 gate2876(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2877(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2878(.a(G2), .O(gate77inter7));
  inv1  gate2879(.a(G320), .O(gate77inter8));
  nand2 gate2880(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2881(.a(s_333), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2882(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2883(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2884(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2605(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2606(.a(gate90inter0), .b(s_294), .O(gate90inter1));
  and2  gate2607(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2608(.a(s_294), .O(gate90inter3));
  inv1  gate2609(.a(s_295), .O(gate90inter4));
  nand2 gate2610(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2611(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2612(.a(G21), .O(gate90inter7));
  inv1  gate2613(.a(G338), .O(gate90inter8));
  nand2 gate2614(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2615(.a(s_295), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2616(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2617(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2618(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate701(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate702(.a(gate92inter0), .b(s_22), .O(gate92inter1));
  and2  gate703(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate704(.a(s_22), .O(gate92inter3));
  inv1  gate705(.a(s_23), .O(gate92inter4));
  nand2 gate706(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate707(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate708(.a(G29), .O(gate92inter7));
  inv1  gate709(.a(G341), .O(gate92inter8));
  nand2 gate710(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate711(.a(s_23), .b(gate92inter3), .O(gate92inter10));
  nor2  gate712(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate713(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate714(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1401(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1402(.a(gate93inter0), .b(s_122), .O(gate93inter1));
  and2  gate1403(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1404(.a(s_122), .O(gate93inter3));
  inv1  gate1405(.a(s_123), .O(gate93inter4));
  nand2 gate1406(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1407(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1408(.a(G18), .O(gate93inter7));
  inv1  gate1409(.a(G344), .O(gate93inter8));
  nand2 gate1410(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1411(.a(s_123), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1412(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1413(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1414(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate2255(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2256(.a(gate94inter0), .b(s_244), .O(gate94inter1));
  and2  gate2257(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2258(.a(s_244), .O(gate94inter3));
  inv1  gate2259(.a(s_245), .O(gate94inter4));
  nand2 gate2260(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2261(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2262(.a(G22), .O(gate94inter7));
  inv1  gate2263(.a(G344), .O(gate94inter8));
  nand2 gate2264(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2265(.a(s_245), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2266(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2267(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2268(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1499(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1500(.a(gate96inter0), .b(s_136), .O(gate96inter1));
  and2  gate1501(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1502(.a(s_136), .O(gate96inter3));
  inv1  gate1503(.a(s_137), .O(gate96inter4));
  nand2 gate1504(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1505(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1506(.a(G30), .O(gate96inter7));
  inv1  gate1507(.a(G347), .O(gate96inter8));
  nand2 gate1508(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1509(.a(s_137), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1510(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1511(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1512(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1835(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1836(.a(gate97inter0), .b(s_184), .O(gate97inter1));
  and2  gate1837(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1838(.a(s_184), .O(gate97inter3));
  inv1  gate1839(.a(s_185), .O(gate97inter4));
  nand2 gate1840(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1841(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1842(.a(G19), .O(gate97inter7));
  inv1  gate1843(.a(G350), .O(gate97inter8));
  nand2 gate1844(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1845(.a(s_185), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1846(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1847(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1848(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1023(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1024(.a(gate98inter0), .b(s_68), .O(gate98inter1));
  and2  gate1025(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1026(.a(s_68), .O(gate98inter3));
  inv1  gate1027(.a(s_69), .O(gate98inter4));
  nand2 gate1028(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1029(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1030(.a(G23), .O(gate98inter7));
  inv1  gate1031(.a(G350), .O(gate98inter8));
  nand2 gate1032(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1033(.a(s_69), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1034(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1035(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1036(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1639(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1640(.a(gate102inter0), .b(s_156), .O(gate102inter1));
  and2  gate1641(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1642(.a(s_156), .O(gate102inter3));
  inv1  gate1643(.a(s_157), .O(gate102inter4));
  nand2 gate1644(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1645(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1646(.a(G24), .O(gate102inter7));
  inv1  gate1647(.a(G356), .O(gate102inter8));
  nand2 gate1648(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1649(.a(s_157), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1650(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1651(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1652(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1107(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1108(.a(gate103inter0), .b(s_80), .O(gate103inter1));
  and2  gate1109(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1110(.a(s_80), .O(gate103inter3));
  inv1  gate1111(.a(s_81), .O(gate103inter4));
  nand2 gate1112(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1113(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1114(.a(G28), .O(gate103inter7));
  inv1  gate1115(.a(G359), .O(gate103inter8));
  nand2 gate1116(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1117(.a(s_81), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1118(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1119(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1120(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1667(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1668(.a(gate104inter0), .b(s_160), .O(gate104inter1));
  and2  gate1669(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1670(.a(s_160), .O(gate104inter3));
  inv1  gate1671(.a(s_161), .O(gate104inter4));
  nand2 gate1672(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1673(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1674(.a(G32), .O(gate104inter7));
  inv1  gate1675(.a(G359), .O(gate104inter8));
  nand2 gate1676(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1677(.a(s_161), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1678(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1679(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1680(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2577(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2578(.a(gate106inter0), .b(s_290), .O(gate106inter1));
  and2  gate2579(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2580(.a(s_290), .O(gate106inter3));
  inv1  gate2581(.a(s_291), .O(gate106inter4));
  nand2 gate2582(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2583(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2584(.a(G364), .O(gate106inter7));
  inv1  gate2585(.a(G365), .O(gate106inter8));
  nand2 gate2586(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2587(.a(s_291), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2588(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2589(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2590(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate2731(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2732(.a(gate109inter0), .b(s_312), .O(gate109inter1));
  and2  gate2733(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2734(.a(s_312), .O(gate109inter3));
  inv1  gate2735(.a(s_313), .O(gate109inter4));
  nand2 gate2736(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2737(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2738(.a(G370), .O(gate109inter7));
  inv1  gate2739(.a(G371), .O(gate109inter8));
  nand2 gate2740(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2741(.a(s_313), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2742(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2743(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2744(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1303(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1304(.a(gate110inter0), .b(s_108), .O(gate110inter1));
  and2  gate1305(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1306(.a(s_108), .O(gate110inter3));
  inv1  gate1307(.a(s_109), .O(gate110inter4));
  nand2 gate1308(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1309(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1310(.a(G372), .O(gate110inter7));
  inv1  gate1311(.a(G373), .O(gate110inter8));
  nand2 gate1312(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1313(.a(s_109), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1314(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1315(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1316(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1261(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1262(.a(gate111inter0), .b(s_102), .O(gate111inter1));
  and2  gate1263(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1264(.a(s_102), .O(gate111inter3));
  inv1  gate1265(.a(s_103), .O(gate111inter4));
  nand2 gate1266(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1267(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1268(.a(G374), .O(gate111inter7));
  inv1  gate1269(.a(G375), .O(gate111inter8));
  nand2 gate1270(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1271(.a(s_103), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1272(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1273(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1274(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2199(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2200(.a(gate112inter0), .b(s_236), .O(gate112inter1));
  and2  gate2201(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2202(.a(s_236), .O(gate112inter3));
  inv1  gate2203(.a(s_237), .O(gate112inter4));
  nand2 gate2204(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2205(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2206(.a(G376), .O(gate112inter7));
  inv1  gate2207(.a(G377), .O(gate112inter8));
  nand2 gate2208(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2209(.a(s_237), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2210(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2211(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2212(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate995(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate996(.a(gate113inter0), .b(s_64), .O(gate113inter1));
  and2  gate997(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate998(.a(s_64), .O(gate113inter3));
  inv1  gate999(.a(s_65), .O(gate113inter4));
  nand2 gate1000(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1001(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1002(.a(G378), .O(gate113inter7));
  inv1  gate1003(.a(G379), .O(gate113inter8));
  nand2 gate1004(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1005(.a(s_65), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1006(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1007(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1008(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate2017(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2018(.a(gate114inter0), .b(s_210), .O(gate114inter1));
  and2  gate2019(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2020(.a(s_210), .O(gate114inter3));
  inv1  gate2021(.a(s_211), .O(gate114inter4));
  nand2 gate2022(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2023(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2024(.a(G380), .O(gate114inter7));
  inv1  gate2025(.a(G381), .O(gate114inter8));
  nand2 gate2026(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2027(.a(s_211), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2028(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2029(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2030(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2437(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2438(.a(gate116inter0), .b(s_270), .O(gate116inter1));
  and2  gate2439(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2440(.a(s_270), .O(gate116inter3));
  inv1  gate2441(.a(s_271), .O(gate116inter4));
  nand2 gate2442(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2443(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2444(.a(G384), .O(gate116inter7));
  inv1  gate2445(.a(G385), .O(gate116inter8));
  nand2 gate2446(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2447(.a(s_271), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2448(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2449(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2450(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate729(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate730(.a(gate119inter0), .b(s_26), .O(gate119inter1));
  and2  gate731(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate732(.a(s_26), .O(gate119inter3));
  inv1  gate733(.a(s_27), .O(gate119inter4));
  nand2 gate734(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate735(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate736(.a(G390), .O(gate119inter7));
  inv1  gate737(.a(G391), .O(gate119inter8));
  nand2 gate738(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate739(.a(s_27), .b(gate119inter3), .O(gate119inter10));
  nor2  gate740(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate741(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate742(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2591(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2592(.a(gate124inter0), .b(s_292), .O(gate124inter1));
  and2  gate2593(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2594(.a(s_292), .O(gate124inter3));
  inv1  gate2595(.a(s_293), .O(gate124inter4));
  nand2 gate2596(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2597(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2598(.a(G400), .O(gate124inter7));
  inv1  gate2599(.a(G401), .O(gate124inter8));
  nand2 gate2600(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2601(.a(s_293), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2602(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2603(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2604(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2535(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2536(.a(gate127inter0), .b(s_284), .O(gate127inter1));
  and2  gate2537(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2538(.a(s_284), .O(gate127inter3));
  inv1  gate2539(.a(s_285), .O(gate127inter4));
  nand2 gate2540(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2541(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2542(.a(G406), .O(gate127inter7));
  inv1  gate2543(.a(G407), .O(gate127inter8));
  nand2 gate2544(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2545(.a(s_285), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2546(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2547(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2548(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1527(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1528(.a(gate131inter0), .b(s_140), .O(gate131inter1));
  and2  gate1529(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1530(.a(s_140), .O(gate131inter3));
  inv1  gate1531(.a(s_141), .O(gate131inter4));
  nand2 gate1532(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1533(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1534(.a(G414), .O(gate131inter7));
  inv1  gate1535(.a(G415), .O(gate131inter8));
  nand2 gate1536(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1537(.a(s_141), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1538(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1539(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1540(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate827(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate828(.a(gate132inter0), .b(s_40), .O(gate132inter1));
  and2  gate829(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate830(.a(s_40), .O(gate132inter3));
  inv1  gate831(.a(s_41), .O(gate132inter4));
  nand2 gate832(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate833(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate834(.a(G416), .O(gate132inter7));
  inv1  gate835(.a(G417), .O(gate132inter8));
  nand2 gate836(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate837(.a(s_41), .b(gate132inter3), .O(gate132inter10));
  nor2  gate838(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate839(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate840(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate855(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate856(.a(gate135inter0), .b(s_44), .O(gate135inter1));
  and2  gate857(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate858(.a(s_44), .O(gate135inter3));
  inv1  gate859(.a(s_45), .O(gate135inter4));
  nand2 gate860(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate861(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate862(.a(G422), .O(gate135inter7));
  inv1  gate863(.a(G423), .O(gate135inter8));
  nand2 gate864(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate865(.a(s_45), .b(gate135inter3), .O(gate135inter10));
  nor2  gate866(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate867(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate868(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2353(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2354(.a(gate137inter0), .b(s_258), .O(gate137inter1));
  and2  gate2355(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2356(.a(s_258), .O(gate137inter3));
  inv1  gate2357(.a(s_259), .O(gate137inter4));
  nand2 gate2358(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2359(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2360(.a(G426), .O(gate137inter7));
  inv1  gate2361(.a(G429), .O(gate137inter8));
  nand2 gate2362(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2363(.a(s_259), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2364(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2365(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2366(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2745(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2746(.a(gate141inter0), .b(s_314), .O(gate141inter1));
  and2  gate2747(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2748(.a(s_314), .O(gate141inter3));
  inv1  gate2749(.a(s_315), .O(gate141inter4));
  nand2 gate2750(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2751(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2752(.a(G450), .O(gate141inter7));
  inv1  gate2753(.a(G453), .O(gate141inter8));
  nand2 gate2754(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2755(.a(s_315), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2756(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2757(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2758(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate3053(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate3054(.a(gate143inter0), .b(s_358), .O(gate143inter1));
  and2  gate3055(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate3056(.a(s_358), .O(gate143inter3));
  inv1  gate3057(.a(s_359), .O(gate143inter4));
  nand2 gate3058(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate3059(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate3060(.a(G462), .O(gate143inter7));
  inv1  gate3061(.a(G465), .O(gate143inter8));
  nand2 gate3062(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate3063(.a(s_359), .b(gate143inter3), .O(gate143inter10));
  nor2  gate3064(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate3065(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate3066(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate3039(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate3040(.a(gate148inter0), .b(s_356), .O(gate148inter1));
  and2  gate3041(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate3042(.a(s_356), .O(gate148inter3));
  inv1  gate3043(.a(s_357), .O(gate148inter4));
  nand2 gate3044(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate3045(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate3046(.a(G492), .O(gate148inter7));
  inv1  gate3047(.a(G495), .O(gate148inter8));
  nand2 gate3048(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate3049(.a(s_357), .b(gate148inter3), .O(gate148inter10));
  nor2  gate3050(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate3051(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate3052(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1513(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1514(.a(gate151inter0), .b(s_138), .O(gate151inter1));
  and2  gate1515(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1516(.a(s_138), .O(gate151inter3));
  inv1  gate1517(.a(s_139), .O(gate151inter4));
  nand2 gate1518(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1519(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1520(.a(G510), .O(gate151inter7));
  inv1  gate1521(.a(G513), .O(gate151inter8));
  nand2 gate1522(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1523(.a(s_139), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1524(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1525(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1526(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2661(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2662(.a(gate152inter0), .b(s_302), .O(gate152inter1));
  and2  gate2663(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2664(.a(s_302), .O(gate152inter3));
  inv1  gate2665(.a(s_303), .O(gate152inter4));
  nand2 gate2666(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2667(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2668(.a(G516), .O(gate152inter7));
  inv1  gate2669(.a(G519), .O(gate152inter8));
  nand2 gate2670(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2671(.a(s_303), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2672(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2673(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2674(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate575(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate576(.a(gate154inter0), .b(s_4), .O(gate154inter1));
  and2  gate577(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate578(.a(s_4), .O(gate154inter3));
  inv1  gate579(.a(s_5), .O(gate154inter4));
  nand2 gate580(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate581(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate582(.a(G429), .O(gate154inter7));
  inv1  gate583(.a(G522), .O(gate154inter8));
  nand2 gate584(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate585(.a(s_5), .b(gate154inter3), .O(gate154inter10));
  nor2  gate586(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate587(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate588(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1611(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1612(.a(gate155inter0), .b(s_152), .O(gate155inter1));
  and2  gate1613(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1614(.a(s_152), .O(gate155inter3));
  inv1  gate1615(.a(s_153), .O(gate155inter4));
  nand2 gate1616(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1617(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1618(.a(G432), .O(gate155inter7));
  inv1  gate1619(.a(G525), .O(gate155inter8));
  nand2 gate1620(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1621(.a(s_153), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1622(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1623(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1624(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1247(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1248(.a(gate156inter0), .b(s_100), .O(gate156inter1));
  and2  gate1249(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1250(.a(s_100), .O(gate156inter3));
  inv1  gate1251(.a(s_101), .O(gate156inter4));
  nand2 gate1252(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1253(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1254(.a(G435), .O(gate156inter7));
  inv1  gate1255(.a(G525), .O(gate156inter8));
  nand2 gate1256(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1257(.a(s_101), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1258(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1259(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1260(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2213(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2214(.a(gate157inter0), .b(s_238), .O(gate157inter1));
  and2  gate2215(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2216(.a(s_238), .O(gate157inter3));
  inv1  gate2217(.a(s_239), .O(gate157inter4));
  nand2 gate2218(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2219(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2220(.a(G438), .O(gate157inter7));
  inv1  gate2221(.a(G528), .O(gate157inter8));
  nand2 gate2222(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2223(.a(s_239), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2224(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2225(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2226(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate645(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate646(.a(gate158inter0), .b(s_14), .O(gate158inter1));
  and2  gate647(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate648(.a(s_14), .O(gate158inter3));
  inv1  gate649(.a(s_15), .O(gate158inter4));
  nand2 gate650(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate651(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate652(.a(G441), .O(gate158inter7));
  inv1  gate653(.a(G528), .O(gate158inter8));
  nand2 gate654(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate655(.a(s_15), .b(gate158inter3), .O(gate158inter10));
  nor2  gate656(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate657(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate658(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1373(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1374(.a(gate160inter0), .b(s_118), .O(gate160inter1));
  and2  gate1375(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1376(.a(s_118), .O(gate160inter3));
  inv1  gate1377(.a(s_119), .O(gate160inter4));
  nand2 gate1378(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1379(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1380(.a(G447), .O(gate160inter7));
  inv1  gate1381(.a(G531), .O(gate160inter8));
  nand2 gate1382(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1383(.a(s_119), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1384(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1385(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1386(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1051(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1052(.a(gate161inter0), .b(s_72), .O(gate161inter1));
  and2  gate1053(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1054(.a(s_72), .O(gate161inter3));
  inv1  gate1055(.a(s_73), .O(gate161inter4));
  nand2 gate1056(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1057(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1058(.a(G450), .O(gate161inter7));
  inv1  gate1059(.a(G534), .O(gate161inter8));
  nand2 gate1060(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1061(.a(s_73), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1062(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1063(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1064(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2941(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2942(.a(gate164inter0), .b(s_342), .O(gate164inter1));
  and2  gate2943(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2944(.a(s_342), .O(gate164inter3));
  inv1  gate2945(.a(s_343), .O(gate164inter4));
  nand2 gate2946(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2947(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2948(.a(G459), .O(gate164inter7));
  inv1  gate2949(.a(G537), .O(gate164inter8));
  nand2 gate2950(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2951(.a(s_343), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2952(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2953(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2954(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2927(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2928(.a(gate172inter0), .b(s_340), .O(gate172inter1));
  and2  gate2929(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2930(.a(s_340), .O(gate172inter3));
  inv1  gate2931(.a(s_341), .O(gate172inter4));
  nand2 gate2932(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2933(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2934(.a(G483), .O(gate172inter7));
  inv1  gate2935(.a(G549), .O(gate172inter8));
  nand2 gate2936(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2937(.a(s_341), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2938(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2939(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2940(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1653(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1654(.a(gate175inter0), .b(s_158), .O(gate175inter1));
  and2  gate1655(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1656(.a(s_158), .O(gate175inter3));
  inv1  gate1657(.a(s_159), .O(gate175inter4));
  nand2 gate1658(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1659(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1660(.a(G492), .O(gate175inter7));
  inv1  gate1661(.a(G555), .O(gate175inter8));
  nand2 gate1662(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1663(.a(s_159), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1664(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1665(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1666(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1289(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1290(.a(gate176inter0), .b(s_106), .O(gate176inter1));
  and2  gate1291(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1292(.a(s_106), .O(gate176inter3));
  inv1  gate1293(.a(s_107), .O(gate176inter4));
  nand2 gate1294(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1295(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1296(.a(G495), .O(gate176inter7));
  inv1  gate1297(.a(G555), .O(gate176inter8));
  nand2 gate1298(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1299(.a(s_107), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1300(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1301(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1302(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1457(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1458(.a(gate180inter0), .b(s_130), .O(gate180inter1));
  and2  gate1459(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1460(.a(s_130), .O(gate180inter3));
  inv1  gate1461(.a(s_131), .O(gate180inter4));
  nand2 gate1462(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1463(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1464(.a(G507), .O(gate180inter7));
  inv1  gate1465(.a(G561), .O(gate180inter8));
  nand2 gate1466(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1467(.a(s_131), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1468(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1469(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1470(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1863(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1864(.a(gate185inter0), .b(s_188), .O(gate185inter1));
  and2  gate1865(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1866(.a(s_188), .O(gate185inter3));
  inv1  gate1867(.a(s_189), .O(gate185inter4));
  nand2 gate1868(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1869(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1870(.a(G570), .O(gate185inter7));
  inv1  gate1871(.a(G571), .O(gate185inter8));
  nand2 gate1872(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1873(.a(s_189), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1874(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1875(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1876(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate897(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate898(.a(gate186inter0), .b(s_50), .O(gate186inter1));
  and2  gate899(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate900(.a(s_50), .O(gate186inter3));
  inv1  gate901(.a(s_51), .O(gate186inter4));
  nand2 gate902(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate903(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate904(.a(G572), .O(gate186inter7));
  inv1  gate905(.a(G573), .O(gate186inter8));
  nand2 gate906(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate907(.a(s_51), .b(gate186inter3), .O(gate186inter10));
  nor2  gate908(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate909(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate910(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate743(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate744(.a(gate188inter0), .b(s_28), .O(gate188inter1));
  and2  gate745(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate746(.a(s_28), .O(gate188inter3));
  inv1  gate747(.a(s_29), .O(gate188inter4));
  nand2 gate748(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate749(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate750(.a(G576), .O(gate188inter7));
  inv1  gate751(.a(G577), .O(gate188inter8));
  nand2 gate752(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate753(.a(s_29), .b(gate188inter3), .O(gate188inter10));
  nor2  gate754(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate755(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate756(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2451(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2452(.a(gate190inter0), .b(s_272), .O(gate190inter1));
  and2  gate2453(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2454(.a(s_272), .O(gate190inter3));
  inv1  gate2455(.a(s_273), .O(gate190inter4));
  nand2 gate2456(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2457(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2458(.a(G580), .O(gate190inter7));
  inv1  gate2459(.a(G581), .O(gate190inter8));
  nand2 gate2460(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2461(.a(s_273), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2462(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2463(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2464(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2689(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2690(.a(gate191inter0), .b(s_306), .O(gate191inter1));
  and2  gate2691(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2692(.a(s_306), .O(gate191inter3));
  inv1  gate2693(.a(s_307), .O(gate191inter4));
  nand2 gate2694(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2695(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2696(.a(G582), .O(gate191inter7));
  inv1  gate2697(.a(G583), .O(gate191inter8));
  nand2 gate2698(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2699(.a(s_307), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2700(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2701(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2702(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate3011(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate3012(.a(gate192inter0), .b(s_352), .O(gate192inter1));
  and2  gate3013(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate3014(.a(s_352), .O(gate192inter3));
  inv1  gate3015(.a(s_353), .O(gate192inter4));
  nand2 gate3016(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate3017(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate3018(.a(G584), .O(gate192inter7));
  inv1  gate3019(.a(G585), .O(gate192inter8));
  nand2 gate3020(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate3021(.a(s_353), .b(gate192inter3), .O(gate192inter10));
  nor2  gate3022(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate3023(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate3024(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1093(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1094(.a(gate194inter0), .b(s_78), .O(gate194inter1));
  and2  gate1095(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1096(.a(s_78), .O(gate194inter3));
  inv1  gate1097(.a(s_79), .O(gate194inter4));
  nand2 gate1098(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1099(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1100(.a(G588), .O(gate194inter7));
  inv1  gate1101(.a(G589), .O(gate194inter8));
  nand2 gate1102(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1103(.a(s_79), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1104(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1105(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1106(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2955(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2956(.a(gate197inter0), .b(s_344), .O(gate197inter1));
  and2  gate2957(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2958(.a(s_344), .O(gate197inter3));
  inv1  gate2959(.a(s_345), .O(gate197inter4));
  nand2 gate2960(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2961(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2962(.a(G594), .O(gate197inter7));
  inv1  gate2963(.a(G595), .O(gate197inter8));
  nand2 gate2964(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2965(.a(s_345), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2966(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2967(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2968(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1961(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1962(.a(gate198inter0), .b(s_202), .O(gate198inter1));
  and2  gate1963(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1964(.a(s_202), .O(gate198inter3));
  inv1  gate1965(.a(s_203), .O(gate198inter4));
  nand2 gate1966(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1967(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1968(.a(G596), .O(gate198inter7));
  inv1  gate1969(.a(G597), .O(gate198inter8));
  nand2 gate1970(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1971(.a(s_203), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1972(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1973(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1974(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1163(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1164(.a(gate207inter0), .b(s_88), .O(gate207inter1));
  and2  gate1165(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1166(.a(s_88), .O(gate207inter3));
  inv1  gate1167(.a(s_89), .O(gate207inter4));
  nand2 gate1168(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1169(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1170(.a(G622), .O(gate207inter7));
  inv1  gate1171(.a(G632), .O(gate207inter8));
  nand2 gate1172(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1173(.a(s_89), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1174(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1175(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1176(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2717(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2718(.a(gate208inter0), .b(s_310), .O(gate208inter1));
  and2  gate2719(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2720(.a(s_310), .O(gate208inter3));
  inv1  gate2721(.a(s_311), .O(gate208inter4));
  nand2 gate2722(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2723(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2724(.a(G627), .O(gate208inter7));
  inv1  gate2725(.a(G637), .O(gate208inter8));
  nand2 gate2726(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2727(.a(s_311), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2728(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2729(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2730(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2549(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2550(.a(gate209inter0), .b(s_286), .O(gate209inter1));
  and2  gate2551(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2552(.a(s_286), .O(gate209inter3));
  inv1  gate2553(.a(s_287), .O(gate209inter4));
  nand2 gate2554(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2555(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2556(.a(G602), .O(gate209inter7));
  inv1  gate2557(.a(G666), .O(gate209inter8));
  nand2 gate2558(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2559(.a(s_287), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2560(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2561(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2562(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate3025(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate3026(.a(gate214inter0), .b(s_354), .O(gate214inter1));
  and2  gate3027(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate3028(.a(s_354), .O(gate214inter3));
  inv1  gate3029(.a(s_355), .O(gate214inter4));
  nand2 gate3030(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate3031(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate3032(.a(G612), .O(gate214inter7));
  inv1  gate3033(.a(G672), .O(gate214inter8));
  nand2 gate3034(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate3035(.a(s_355), .b(gate214inter3), .O(gate214inter10));
  nor2  gate3036(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate3037(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate3038(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1065(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1066(.a(gate215inter0), .b(s_74), .O(gate215inter1));
  and2  gate1067(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1068(.a(s_74), .O(gate215inter3));
  inv1  gate1069(.a(s_75), .O(gate215inter4));
  nand2 gate1070(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1071(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1072(.a(G607), .O(gate215inter7));
  inv1  gate1073(.a(G675), .O(gate215inter8));
  nand2 gate1074(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1075(.a(s_75), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1076(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1077(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1078(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2381(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2382(.a(gate217inter0), .b(s_262), .O(gate217inter1));
  and2  gate2383(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2384(.a(s_262), .O(gate217inter3));
  inv1  gate2385(.a(s_263), .O(gate217inter4));
  nand2 gate2386(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2387(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2388(.a(G622), .O(gate217inter7));
  inv1  gate2389(.a(G678), .O(gate217inter8));
  nand2 gate2390(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2391(.a(s_263), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2392(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2393(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2394(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate757(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate758(.a(gate222inter0), .b(s_30), .O(gate222inter1));
  and2  gate759(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate760(.a(s_30), .O(gate222inter3));
  inv1  gate761(.a(s_31), .O(gate222inter4));
  nand2 gate762(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate763(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate764(.a(G632), .O(gate222inter7));
  inv1  gate765(.a(G684), .O(gate222inter8));
  nand2 gate766(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate767(.a(s_31), .b(gate222inter3), .O(gate222inter10));
  nor2  gate768(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate769(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate770(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1765(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1766(.a(gate225inter0), .b(s_174), .O(gate225inter1));
  and2  gate1767(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1768(.a(s_174), .O(gate225inter3));
  inv1  gate1769(.a(s_175), .O(gate225inter4));
  nand2 gate1770(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1771(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1772(.a(G690), .O(gate225inter7));
  inv1  gate1773(.a(G691), .O(gate225inter8));
  nand2 gate1774(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1775(.a(s_175), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1776(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1777(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1778(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate2101(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate2102(.a(gate226inter0), .b(s_222), .O(gate226inter1));
  and2  gate2103(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate2104(.a(s_222), .O(gate226inter3));
  inv1  gate2105(.a(s_223), .O(gate226inter4));
  nand2 gate2106(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate2107(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate2108(.a(G692), .O(gate226inter7));
  inv1  gate2109(.a(G693), .O(gate226inter8));
  nand2 gate2110(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate2111(.a(s_223), .b(gate226inter3), .O(gate226inter10));
  nor2  gate2112(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate2113(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate2114(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1891(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1892(.a(gate228inter0), .b(s_192), .O(gate228inter1));
  and2  gate1893(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1894(.a(s_192), .O(gate228inter3));
  inv1  gate1895(.a(s_193), .O(gate228inter4));
  nand2 gate1896(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1897(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1898(.a(G696), .O(gate228inter7));
  inv1  gate1899(.a(G697), .O(gate228inter8));
  nand2 gate1900(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1901(.a(s_193), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1902(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1903(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1904(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1821(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1822(.a(gate230inter0), .b(s_182), .O(gate230inter1));
  and2  gate1823(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1824(.a(s_182), .O(gate230inter3));
  inv1  gate1825(.a(s_183), .O(gate230inter4));
  nand2 gate1826(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1827(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1828(.a(G700), .O(gate230inter7));
  inv1  gate1829(.a(G701), .O(gate230inter8));
  nand2 gate1830(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1831(.a(s_183), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1832(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1833(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1834(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2185(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2186(.a(gate231inter0), .b(s_234), .O(gate231inter1));
  and2  gate2187(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2188(.a(s_234), .O(gate231inter3));
  inv1  gate2189(.a(s_235), .O(gate231inter4));
  nand2 gate2190(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2191(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2192(.a(G702), .O(gate231inter7));
  inv1  gate2193(.a(G703), .O(gate231inter8));
  nand2 gate2194(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2195(.a(s_235), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2196(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2197(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2198(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate631(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate632(.a(gate235inter0), .b(s_12), .O(gate235inter1));
  and2  gate633(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate634(.a(s_12), .O(gate235inter3));
  inv1  gate635(.a(s_13), .O(gate235inter4));
  nand2 gate636(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate637(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate638(.a(G248), .O(gate235inter7));
  inv1  gate639(.a(G724), .O(gate235inter8));
  nand2 gate640(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate641(.a(s_13), .b(gate235inter3), .O(gate235inter10));
  nor2  gate642(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate643(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate644(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate841(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate842(.a(gate237inter0), .b(s_42), .O(gate237inter1));
  and2  gate843(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate844(.a(s_42), .O(gate237inter3));
  inv1  gate845(.a(s_43), .O(gate237inter4));
  nand2 gate846(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate847(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate848(.a(G254), .O(gate237inter7));
  inv1  gate849(.a(G706), .O(gate237inter8));
  nand2 gate850(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate851(.a(s_43), .b(gate237inter3), .O(gate237inter10));
  nor2  gate852(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate853(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate854(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1443(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1444(.a(gate240inter0), .b(s_128), .O(gate240inter1));
  and2  gate1445(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1446(.a(s_128), .O(gate240inter3));
  inv1  gate1447(.a(s_129), .O(gate240inter4));
  nand2 gate1448(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1449(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1450(.a(G263), .O(gate240inter7));
  inv1  gate1451(.a(G715), .O(gate240inter8));
  nand2 gate1452(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1453(.a(s_129), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1454(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1455(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1456(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate2325(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2326(.a(gate241inter0), .b(s_254), .O(gate241inter1));
  and2  gate2327(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2328(.a(s_254), .O(gate241inter3));
  inv1  gate2329(.a(s_255), .O(gate241inter4));
  nand2 gate2330(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2331(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2332(.a(G242), .O(gate241inter7));
  inv1  gate2333(.a(G730), .O(gate241inter8));
  nand2 gate2334(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2335(.a(s_255), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2336(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2337(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2338(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate603(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate604(.a(gate243inter0), .b(s_8), .O(gate243inter1));
  and2  gate605(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate606(.a(s_8), .O(gate243inter3));
  inv1  gate607(.a(s_9), .O(gate243inter4));
  nand2 gate608(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate609(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate610(.a(G245), .O(gate243inter7));
  inv1  gate611(.a(G733), .O(gate243inter8));
  nand2 gate612(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate613(.a(s_9), .b(gate243inter3), .O(gate243inter10));
  nor2  gate614(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate615(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate616(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate2479(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2480(.a(gate244inter0), .b(s_276), .O(gate244inter1));
  and2  gate2481(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2482(.a(s_276), .O(gate244inter3));
  inv1  gate2483(.a(s_277), .O(gate244inter4));
  nand2 gate2484(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2485(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2486(.a(G721), .O(gate244inter7));
  inv1  gate2487(.a(G733), .O(gate244inter8));
  nand2 gate2488(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2489(.a(s_277), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2490(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2491(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2492(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate799(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate800(.a(gate245inter0), .b(s_36), .O(gate245inter1));
  and2  gate801(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate802(.a(s_36), .O(gate245inter3));
  inv1  gate803(.a(s_37), .O(gate245inter4));
  nand2 gate804(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate805(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate806(.a(G248), .O(gate245inter7));
  inv1  gate807(.a(G736), .O(gate245inter8));
  nand2 gate808(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate809(.a(s_37), .b(gate245inter3), .O(gate245inter10));
  nor2  gate810(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate811(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate812(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2787(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2788(.a(gate246inter0), .b(s_320), .O(gate246inter1));
  and2  gate2789(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2790(.a(s_320), .O(gate246inter3));
  inv1  gate2791(.a(s_321), .O(gate246inter4));
  nand2 gate2792(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2793(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2794(.a(G724), .O(gate246inter7));
  inv1  gate2795(.a(G736), .O(gate246inter8));
  nand2 gate2796(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2797(.a(s_321), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2798(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2799(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2800(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2171(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2172(.a(gate248inter0), .b(s_232), .O(gate248inter1));
  and2  gate2173(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2174(.a(s_232), .O(gate248inter3));
  inv1  gate2175(.a(s_233), .O(gate248inter4));
  nand2 gate2176(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2177(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2178(.a(G727), .O(gate248inter7));
  inv1  gate2179(.a(G739), .O(gate248inter8));
  nand2 gate2180(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2181(.a(s_233), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2182(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2183(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2184(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2521(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2522(.a(gate249inter0), .b(s_282), .O(gate249inter1));
  and2  gate2523(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2524(.a(s_282), .O(gate249inter3));
  inv1  gate2525(.a(s_283), .O(gate249inter4));
  nand2 gate2526(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2527(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2528(.a(G254), .O(gate249inter7));
  inv1  gate2529(.a(G742), .O(gate249inter8));
  nand2 gate2530(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2531(.a(s_283), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2532(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2533(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2534(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2885(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2886(.a(gate251inter0), .b(s_334), .O(gate251inter1));
  and2  gate2887(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2888(.a(s_334), .O(gate251inter3));
  inv1  gate2889(.a(s_335), .O(gate251inter4));
  nand2 gate2890(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2891(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2892(.a(G257), .O(gate251inter7));
  inv1  gate2893(.a(G745), .O(gate251inter8));
  nand2 gate2894(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2895(.a(s_335), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2896(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2897(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2898(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2339(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2340(.a(gate253inter0), .b(s_256), .O(gate253inter1));
  and2  gate2341(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2342(.a(s_256), .O(gate253inter3));
  inv1  gate2343(.a(s_257), .O(gate253inter4));
  nand2 gate2344(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2345(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2346(.a(G260), .O(gate253inter7));
  inv1  gate2347(.a(G748), .O(gate253inter8));
  nand2 gate2348(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2349(.a(s_257), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2350(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2351(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2352(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1037(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1038(.a(gate255inter0), .b(s_70), .O(gate255inter1));
  and2  gate1039(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1040(.a(s_70), .O(gate255inter3));
  inv1  gate1041(.a(s_71), .O(gate255inter4));
  nand2 gate1042(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1043(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1044(.a(G263), .O(gate255inter7));
  inv1  gate1045(.a(G751), .O(gate255inter8));
  nand2 gate1046(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1047(.a(s_71), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1048(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1049(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1050(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2773(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2774(.a(gate257inter0), .b(s_318), .O(gate257inter1));
  and2  gate2775(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2776(.a(s_318), .O(gate257inter3));
  inv1  gate2777(.a(s_319), .O(gate257inter4));
  nand2 gate2778(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2779(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2780(.a(G754), .O(gate257inter7));
  inv1  gate2781(.a(G755), .O(gate257inter8));
  nand2 gate2782(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2783(.a(s_319), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2784(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2785(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2786(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1233(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1234(.a(gate259inter0), .b(s_98), .O(gate259inter1));
  and2  gate1235(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1236(.a(s_98), .O(gate259inter3));
  inv1  gate1237(.a(s_99), .O(gate259inter4));
  nand2 gate1238(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1239(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1240(.a(G758), .O(gate259inter7));
  inv1  gate1241(.a(G759), .O(gate259inter8));
  nand2 gate1242(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1243(.a(s_99), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1244(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1245(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1246(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1849(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1850(.a(gate261inter0), .b(s_186), .O(gate261inter1));
  and2  gate1851(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1852(.a(s_186), .O(gate261inter3));
  inv1  gate1853(.a(s_187), .O(gate261inter4));
  nand2 gate1854(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1855(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1856(.a(G762), .O(gate261inter7));
  inv1  gate1857(.a(G763), .O(gate261inter8));
  nand2 gate1858(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1859(.a(s_187), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1860(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1861(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1862(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2913(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2914(.a(gate263inter0), .b(s_338), .O(gate263inter1));
  and2  gate2915(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2916(.a(s_338), .O(gate263inter3));
  inv1  gate2917(.a(s_339), .O(gate263inter4));
  nand2 gate2918(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2919(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2920(.a(G766), .O(gate263inter7));
  inv1  gate2921(.a(G767), .O(gate263inter8));
  nand2 gate2922(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2923(.a(s_339), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2924(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2925(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2926(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1737(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1738(.a(gate267inter0), .b(s_170), .O(gate267inter1));
  and2  gate1739(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1740(.a(s_170), .O(gate267inter3));
  inv1  gate1741(.a(s_171), .O(gate267inter4));
  nand2 gate1742(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1743(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1744(.a(G648), .O(gate267inter7));
  inv1  gate1745(.a(G776), .O(gate267inter8));
  nand2 gate1746(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1747(.a(s_171), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1748(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1749(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1750(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2283(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2284(.a(gate268inter0), .b(s_248), .O(gate268inter1));
  and2  gate2285(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2286(.a(s_248), .O(gate268inter3));
  inv1  gate2287(.a(s_249), .O(gate268inter4));
  nand2 gate2288(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2289(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2290(.a(G651), .O(gate268inter7));
  inv1  gate2291(.a(G779), .O(gate268inter8));
  nand2 gate2292(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2293(.a(s_249), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2294(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2295(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2296(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate939(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate940(.a(gate272inter0), .b(s_56), .O(gate272inter1));
  and2  gate941(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate942(.a(s_56), .O(gate272inter3));
  inv1  gate943(.a(s_57), .O(gate272inter4));
  nand2 gate944(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate945(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate946(.a(G663), .O(gate272inter7));
  inv1  gate947(.a(G791), .O(gate272inter8));
  nand2 gate948(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate949(.a(s_57), .b(gate272inter3), .O(gate272inter10));
  nor2  gate950(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate951(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate952(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2675(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2676(.a(gate275inter0), .b(s_304), .O(gate275inter1));
  and2  gate2677(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2678(.a(s_304), .O(gate275inter3));
  inv1  gate2679(.a(s_305), .O(gate275inter4));
  nand2 gate2680(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2681(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2682(.a(G645), .O(gate275inter7));
  inv1  gate2683(.a(G797), .O(gate275inter8));
  nand2 gate2684(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2685(.a(s_305), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2686(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2687(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2688(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1779(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1780(.a(gate277inter0), .b(s_176), .O(gate277inter1));
  and2  gate1781(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1782(.a(s_176), .O(gate277inter3));
  inv1  gate1783(.a(s_177), .O(gate277inter4));
  nand2 gate1784(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1785(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1786(.a(G648), .O(gate277inter7));
  inv1  gate1787(.a(G800), .O(gate277inter8));
  nand2 gate1788(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1789(.a(s_177), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1790(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1791(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1792(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate617(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate618(.a(gate280inter0), .b(s_10), .O(gate280inter1));
  and2  gate619(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate620(.a(s_10), .O(gate280inter3));
  inv1  gate621(.a(s_11), .O(gate280inter4));
  nand2 gate622(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate623(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate624(.a(G779), .O(gate280inter7));
  inv1  gate625(.a(G803), .O(gate280inter8));
  nand2 gate626(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate627(.a(s_11), .b(gate280inter3), .O(gate280inter10));
  nor2  gate628(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate629(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate630(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1625(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1626(.a(gate282inter0), .b(s_154), .O(gate282inter1));
  and2  gate1627(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1628(.a(s_154), .O(gate282inter3));
  inv1  gate1629(.a(s_155), .O(gate282inter4));
  nand2 gate1630(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1631(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1632(.a(G782), .O(gate282inter7));
  inv1  gate1633(.a(G806), .O(gate282inter8));
  nand2 gate1634(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1635(.a(s_155), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1636(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1637(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1638(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate771(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate772(.a(gate284inter0), .b(s_32), .O(gate284inter1));
  and2  gate773(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate774(.a(s_32), .O(gate284inter3));
  inv1  gate775(.a(s_33), .O(gate284inter4));
  nand2 gate776(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate777(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate778(.a(G785), .O(gate284inter7));
  inv1  gate779(.a(G809), .O(gate284inter8));
  nand2 gate780(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate781(.a(s_33), .b(gate284inter3), .O(gate284inter10));
  nor2  gate782(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate783(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate784(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate813(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate814(.a(gate285inter0), .b(s_38), .O(gate285inter1));
  and2  gate815(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate816(.a(s_38), .O(gate285inter3));
  inv1  gate817(.a(s_39), .O(gate285inter4));
  nand2 gate818(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate819(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate820(.a(G660), .O(gate285inter7));
  inv1  gate821(.a(G812), .O(gate285inter8));
  nand2 gate822(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate823(.a(s_39), .b(gate285inter3), .O(gate285inter10));
  nor2  gate824(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate825(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate826(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1919(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1920(.a(gate287inter0), .b(s_196), .O(gate287inter1));
  and2  gate1921(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1922(.a(s_196), .O(gate287inter3));
  inv1  gate1923(.a(s_197), .O(gate287inter4));
  nand2 gate1924(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1925(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1926(.a(G663), .O(gate287inter7));
  inv1  gate1927(.a(G815), .O(gate287inter8));
  nand2 gate1928(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1929(.a(s_197), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1930(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1931(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1932(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate589(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate590(.a(gate288inter0), .b(s_6), .O(gate288inter1));
  and2  gate591(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate592(.a(s_6), .O(gate288inter3));
  inv1  gate593(.a(s_7), .O(gate288inter4));
  nand2 gate594(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate595(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate596(.a(G791), .O(gate288inter7));
  inv1  gate597(.a(G815), .O(gate288inter8));
  nand2 gate598(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate599(.a(s_7), .b(gate288inter3), .O(gate288inter10));
  nor2  gate600(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate601(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate602(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1485(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1486(.a(gate289inter0), .b(s_134), .O(gate289inter1));
  and2  gate1487(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1488(.a(s_134), .O(gate289inter3));
  inv1  gate1489(.a(s_135), .O(gate289inter4));
  nand2 gate1490(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1491(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1492(.a(G818), .O(gate289inter7));
  inv1  gate1493(.a(G819), .O(gate289inter8));
  nand2 gate1494(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1495(.a(s_135), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1496(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1497(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1498(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2801(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2802(.a(gate291inter0), .b(s_322), .O(gate291inter1));
  and2  gate2803(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2804(.a(s_322), .O(gate291inter3));
  inv1  gate2805(.a(s_323), .O(gate291inter4));
  nand2 gate2806(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2807(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2808(.a(G822), .O(gate291inter7));
  inv1  gate2809(.a(G823), .O(gate291inter8));
  nand2 gate2810(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2811(.a(s_323), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2812(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2813(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2814(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1681(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1682(.a(gate292inter0), .b(s_162), .O(gate292inter1));
  and2  gate1683(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1684(.a(s_162), .O(gate292inter3));
  inv1  gate1685(.a(s_163), .O(gate292inter4));
  nand2 gate1686(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1687(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1688(.a(G824), .O(gate292inter7));
  inv1  gate1689(.a(G825), .O(gate292inter8));
  nand2 gate1690(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1691(.a(s_163), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1692(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1693(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1694(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1191(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1192(.a(gate294inter0), .b(s_92), .O(gate294inter1));
  and2  gate1193(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1194(.a(s_92), .O(gate294inter3));
  inv1  gate1195(.a(s_93), .O(gate294inter4));
  nand2 gate1196(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1197(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1198(.a(G832), .O(gate294inter7));
  inv1  gate1199(.a(G833), .O(gate294inter8));
  nand2 gate1200(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1201(.a(s_93), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1202(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1203(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1204(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2619(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2620(.a(gate389inter0), .b(s_296), .O(gate389inter1));
  and2  gate2621(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2622(.a(s_296), .O(gate389inter3));
  inv1  gate2623(.a(s_297), .O(gate389inter4));
  nand2 gate2624(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2625(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2626(.a(G3), .O(gate389inter7));
  inv1  gate2627(.a(G1042), .O(gate389inter8));
  nand2 gate2628(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2629(.a(s_297), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2630(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2631(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2632(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate561(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate562(.a(gate390inter0), .b(s_2), .O(gate390inter1));
  and2  gate563(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate564(.a(s_2), .O(gate390inter3));
  inv1  gate565(.a(s_3), .O(gate390inter4));
  nand2 gate566(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate567(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate568(.a(G4), .O(gate390inter7));
  inv1  gate569(.a(G1045), .O(gate390inter8));
  nand2 gate570(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate571(.a(s_3), .b(gate390inter3), .O(gate390inter10));
  nor2  gate572(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate573(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate574(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1359(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1360(.a(gate393inter0), .b(s_116), .O(gate393inter1));
  and2  gate1361(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1362(.a(s_116), .O(gate393inter3));
  inv1  gate1363(.a(s_117), .O(gate393inter4));
  nand2 gate1364(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1365(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1366(.a(G7), .O(gate393inter7));
  inv1  gate1367(.a(G1054), .O(gate393inter8));
  nand2 gate1368(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1369(.a(s_117), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1370(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1371(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1372(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1541(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1542(.a(gate395inter0), .b(s_142), .O(gate395inter1));
  and2  gate1543(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1544(.a(s_142), .O(gate395inter3));
  inv1  gate1545(.a(s_143), .O(gate395inter4));
  nand2 gate1546(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1547(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1548(.a(G9), .O(gate395inter7));
  inv1  gate1549(.a(G1060), .O(gate395inter8));
  nand2 gate1550(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1551(.a(s_143), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1552(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1553(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1554(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2815(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2816(.a(gate396inter0), .b(s_324), .O(gate396inter1));
  and2  gate2817(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2818(.a(s_324), .O(gate396inter3));
  inv1  gate2819(.a(s_325), .O(gate396inter4));
  nand2 gate2820(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2821(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2822(.a(G10), .O(gate396inter7));
  inv1  gate2823(.a(G1063), .O(gate396inter8));
  nand2 gate2824(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2825(.a(s_325), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2826(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2827(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2828(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2129(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2130(.a(gate400inter0), .b(s_226), .O(gate400inter1));
  and2  gate2131(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2132(.a(s_226), .O(gate400inter3));
  inv1  gate2133(.a(s_227), .O(gate400inter4));
  nand2 gate2134(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2135(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2136(.a(G14), .O(gate400inter7));
  inv1  gate2137(.a(G1075), .O(gate400inter8));
  nand2 gate2138(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2139(.a(s_227), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2140(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2141(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2142(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2563(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2564(.a(gate401inter0), .b(s_288), .O(gate401inter1));
  and2  gate2565(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2566(.a(s_288), .O(gate401inter3));
  inv1  gate2567(.a(s_289), .O(gate401inter4));
  nand2 gate2568(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2569(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2570(.a(G15), .O(gate401inter7));
  inv1  gate2571(.a(G1078), .O(gate401inter8));
  nand2 gate2572(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2573(.a(s_289), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2574(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2575(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2576(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1947(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1948(.a(gate404inter0), .b(s_200), .O(gate404inter1));
  and2  gate1949(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1950(.a(s_200), .O(gate404inter3));
  inv1  gate1951(.a(s_201), .O(gate404inter4));
  nand2 gate1952(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1953(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1954(.a(G18), .O(gate404inter7));
  inv1  gate1955(.a(G1087), .O(gate404inter8));
  nand2 gate1956(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1957(.a(s_201), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1958(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1959(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1960(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2633(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2634(.a(gate406inter0), .b(s_298), .O(gate406inter1));
  and2  gate2635(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2636(.a(s_298), .O(gate406inter3));
  inv1  gate2637(.a(s_299), .O(gate406inter4));
  nand2 gate2638(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2639(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2640(.a(G20), .O(gate406inter7));
  inv1  gate2641(.a(G1093), .O(gate406inter8));
  nand2 gate2642(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2643(.a(s_299), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2644(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2645(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2646(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1205(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1206(.a(gate408inter0), .b(s_94), .O(gate408inter1));
  and2  gate1207(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1208(.a(s_94), .O(gate408inter3));
  inv1  gate1209(.a(s_95), .O(gate408inter4));
  nand2 gate1210(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1211(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1212(.a(G22), .O(gate408inter7));
  inv1  gate1213(.a(G1099), .O(gate408inter8));
  nand2 gate1214(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1215(.a(s_95), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1216(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1217(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1218(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate2157(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2158(.a(gate409inter0), .b(s_230), .O(gate409inter1));
  and2  gate2159(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2160(.a(s_230), .O(gate409inter3));
  inv1  gate2161(.a(s_231), .O(gate409inter4));
  nand2 gate2162(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2163(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2164(.a(G23), .O(gate409inter7));
  inv1  gate2165(.a(G1102), .O(gate409inter8));
  nand2 gate2166(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2167(.a(s_231), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2168(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2169(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2170(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1275(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1276(.a(gate410inter0), .b(s_104), .O(gate410inter1));
  and2  gate1277(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1278(.a(s_104), .O(gate410inter3));
  inv1  gate1279(.a(s_105), .O(gate410inter4));
  nand2 gate1280(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1281(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1282(.a(G24), .O(gate410inter7));
  inv1  gate1283(.a(G1105), .O(gate410inter8));
  nand2 gate1284(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1285(.a(s_105), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1286(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1287(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1288(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate2423(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2424(.a(gate411inter0), .b(s_268), .O(gate411inter1));
  and2  gate2425(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2426(.a(s_268), .O(gate411inter3));
  inv1  gate2427(.a(s_269), .O(gate411inter4));
  nand2 gate2428(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2429(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2430(.a(G25), .O(gate411inter7));
  inv1  gate2431(.a(G1108), .O(gate411inter8));
  nand2 gate2432(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2433(.a(s_269), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2434(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2435(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2436(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1807(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1808(.a(gate412inter0), .b(s_180), .O(gate412inter1));
  and2  gate1809(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1810(.a(s_180), .O(gate412inter3));
  inv1  gate1811(.a(s_181), .O(gate412inter4));
  nand2 gate1812(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1813(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1814(.a(G26), .O(gate412inter7));
  inv1  gate1815(.a(G1111), .O(gate412inter8));
  nand2 gate1816(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1817(.a(s_181), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1818(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1819(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1820(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1793(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1794(.a(gate413inter0), .b(s_178), .O(gate413inter1));
  and2  gate1795(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1796(.a(s_178), .O(gate413inter3));
  inv1  gate1797(.a(s_179), .O(gate413inter4));
  nand2 gate1798(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1799(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1800(.a(G27), .O(gate413inter7));
  inv1  gate1801(.a(G1114), .O(gate413inter8));
  nand2 gate1802(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1803(.a(s_179), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1804(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1805(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1806(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2983(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2984(.a(gate418inter0), .b(s_348), .O(gate418inter1));
  and2  gate2985(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2986(.a(s_348), .O(gate418inter3));
  inv1  gate2987(.a(s_349), .O(gate418inter4));
  nand2 gate2988(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2989(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2990(.a(G32), .O(gate418inter7));
  inv1  gate2991(.a(G1129), .O(gate418inter8));
  nand2 gate2992(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2993(.a(s_349), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2994(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2995(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2996(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate981(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate982(.a(gate419inter0), .b(s_62), .O(gate419inter1));
  and2  gate983(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate984(.a(s_62), .O(gate419inter3));
  inv1  gate985(.a(s_63), .O(gate419inter4));
  nand2 gate986(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate987(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate988(.a(G1), .O(gate419inter7));
  inv1  gate989(.a(G1132), .O(gate419inter8));
  nand2 gate990(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate991(.a(s_63), .b(gate419inter3), .O(gate419inter10));
  nor2  gate992(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate993(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate994(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1177(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1178(.a(gate420inter0), .b(s_90), .O(gate420inter1));
  and2  gate1179(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1180(.a(s_90), .O(gate420inter3));
  inv1  gate1181(.a(s_91), .O(gate420inter4));
  nand2 gate1182(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1183(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1184(.a(G1036), .O(gate420inter7));
  inv1  gate1185(.a(G1132), .O(gate420inter8));
  nand2 gate1186(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1187(.a(s_91), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1188(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1189(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1190(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2703(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2704(.a(gate421inter0), .b(s_308), .O(gate421inter1));
  and2  gate2705(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2706(.a(s_308), .O(gate421inter3));
  inv1  gate2707(.a(s_309), .O(gate421inter4));
  nand2 gate2708(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2709(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2710(.a(G2), .O(gate421inter7));
  inv1  gate2711(.a(G1135), .O(gate421inter8));
  nand2 gate2712(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2713(.a(s_309), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2714(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2715(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2716(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1583(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1584(.a(gate423inter0), .b(s_148), .O(gate423inter1));
  and2  gate1585(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1586(.a(s_148), .O(gate423inter3));
  inv1  gate1587(.a(s_149), .O(gate423inter4));
  nand2 gate1588(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1589(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1590(.a(G3), .O(gate423inter7));
  inv1  gate1591(.a(G1138), .O(gate423inter8));
  nand2 gate1592(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1593(.a(s_149), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1594(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1595(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1596(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2241(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2242(.a(gate428inter0), .b(s_242), .O(gate428inter1));
  and2  gate2243(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2244(.a(s_242), .O(gate428inter3));
  inv1  gate2245(.a(s_243), .O(gate428inter4));
  nand2 gate2246(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2247(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2248(.a(G1048), .O(gate428inter7));
  inv1  gate2249(.a(G1144), .O(gate428inter8));
  nand2 gate2250(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2251(.a(s_243), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2252(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2253(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2254(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate547(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate548(.a(gate431inter0), .b(s_0), .O(gate431inter1));
  and2  gate549(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate550(.a(s_0), .O(gate431inter3));
  inv1  gate551(.a(s_1), .O(gate431inter4));
  nand2 gate552(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate553(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate554(.a(G7), .O(gate431inter7));
  inv1  gate555(.a(G1150), .O(gate431inter8));
  nand2 gate556(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate557(.a(s_1), .b(gate431inter3), .O(gate431inter10));
  nor2  gate558(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate559(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate560(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate883(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate884(.a(gate432inter0), .b(s_48), .O(gate432inter1));
  and2  gate885(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate886(.a(s_48), .O(gate432inter3));
  inv1  gate887(.a(s_49), .O(gate432inter4));
  nand2 gate888(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate889(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate890(.a(G1054), .O(gate432inter7));
  inv1  gate891(.a(G1150), .O(gate432inter8));
  nand2 gate892(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate893(.a(s_49), .b(gate432inter3), .O(gate432inter10));
  nor2  gate894(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate895(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate896(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1877(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1878(.a(gate435inter0), .b(s_190), .O(gate435inter1));
  and2  gate1879(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1880(.a(s_190), .O(gate435inter3));
  inv1  gate1881(.a(s_191), .O(gate435inter4));
  nand2 gate1882(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1883(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1884(.a(G9), .O(gate435inter7));
  inv1  gate1885(.a(G1156), .O(gate435inter8));
  nand2 gate1886(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1887(.a(s_191), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1888(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1889(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1890(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate2143(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2144(.a(gate439inter0), .b(s_228), .O(gate439inter1));
  and2  gate2145(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2146(.a(s_228), .O(gate439inter3));
  inv1  gate2147(.a(s_229), .O(gate439inter4));
  nand2 gate2148(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2149(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2150(.a(G11), .O(gate439inter7));
  inv1  gate2151(.a(G1162), .O(gate439inter8));
  nand2 gate2152(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2153(.a(s_229), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2154(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2155(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2156(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1695(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1696(.a(gate440inter0), .b(s_164), .O(gate440inter1));
  and2  gate1697(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1698(.a(s_164), .O(gate440inter3));
  inv1  gate1699(.a(s_165), .O(gate440inter4));
  nand2 gate1700(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1701(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1702(.a(G1066), .O(gate440inter7));
  inv1  gate1703(.a(G1162), .O(gate440inter8));
  nand2 gate1704(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1705(.a(s_165), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1706(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1707(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1708(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate967(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate968(.a(gate442inter0), .b(s_60), .O(gate442inter1));
  and2  gate969(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate970(.a(s_60), .O(gate442inter3));
  inv1  gate971(.a(s_61), .O(gate442inter4));
  nand2 gate972(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate973(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate974(.a(G1069), .O(gate442inter7));
  inv1  gate975(.a(G1165), .O(gate442inter8));
  nand2 gate976(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate977(.a(s_61), .b(gate442inter3), .O(gate442inter10));
  nor2  gate978(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate979(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate980(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2297(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2298(.a(gate445inter0), .b(s_250), .O(gate445inter1));
  and2  gate2299(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2300(.a(s_250), .O(gate445inter3));
  inv1  gate2301(.a(s_251), .O(gate445inter4));
  nand2 gate2302(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2303(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2304(.a(G14), .O(gate445inter7));
  inv1  gate2305(.a(G1171), .O(gate445inter8));
  nand2 gate2306(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2307(.a(s_251), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2308(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2309(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2310(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1555(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1556(.a(gate446inter0), .b(s_144), .O(gate446inter1));
  and2  gate1557(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1558(.a(s_144), .O(gate446inter3));
  inv1  gate1559(.a(s_145), .O(gate446inter4));
  nand2 gate1560(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1561(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1562(.a(G1075), .O(gate446inter7));
  inv1  gate1563(.a(G1171), .O(gate446inter8));
  nand2 gate1564(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1565(.a(s_145), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1566(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1567(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1568(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2395(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2396(.a(gate447inter0), .b(s_264), .O(gate447inter1));
  and2  gate2397(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2398(.a(s_264), .O(gate447inter3));
  inv1  gate2399(.a(s_265), .O(gate447inter4));
  nand2 gate2400(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2401(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2402(.a(G15), .O(gate447inter7));
  inv1  gate2403(.a(G1174), .O(gate447inter8));
  nand2 gate2404(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2405(.a(s_265), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2406(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2407(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2408(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2969(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2970(.a(gate448inter0), .b(s_346), .O(gate448inter1));
  and2  gate2971(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2972(.a(s_346), .O(gate448inter3));
  inv1  gate2973(.a(s_347), .O(gate448inter4));
  nand2 gate2974(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2975(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2976(.a(G1078), .O(gate448inter7));
  inv1  gate2977(.a(G1174), .O(gate448inter8));
  nand2 gate2978(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2979(.a(s_347), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2980(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2981(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2982(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate785(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate786(.a(gate450inter0), .b(s_34), .O(gate450inter1));
  and2  gate787(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate788(.a(s_34), .O(gate450inter3));
  inv1  gate789(.a(s_35), .O(gate450inter4));
  nand2 gate790(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate791(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate792(.a(G1081), .O(gate450inter7));
  inv1  gate793(.a(G1177), .O(gate450inter8));
  nand2 gate794(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate795(.a(s_35), .b(gate450inter3), .O(gate450inter10));
  nor2  gate796(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate797(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate798(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1121(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1122(.a(gate451inter0), .b(s_82), .O(gate451inter1));
  and2  gate1123(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1124(.a(s_82), .O(gate451inter3));
  inv1  gate1125(.a(s_83), .O(gate451inter4));
  nand2 gate1126(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1127(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1128(.a(G17), .O(gate451inter7));
  inv1  gate1129(.a(G1180), .O(gate451inter8));
  nand2 gate1130(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1131(.a(s_83), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1132(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1133(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1134(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate2465(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2466(.a(gate452inter0), .b(s_274), .O(gate452inter1));
  and2  gate2467(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2468(.a(s_274), .O(gate452inter3));
  inv1  gate2469(.a(s_275), .O(gate452inter4));
  nand2 gate2470(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2471(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2472(.a(G1084), .O(gate452inter7));
  inv1  gate2473(.a(G1180), .O(gate452inter8));
  nand2 gate2474(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2475(.a(s_275), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2476(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2477(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2478(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1751(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1752(.a(gate454inter0), .b(s_172), .O(gate454inter1));
  and2  gate1753(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1754(.a(s_172), .O(gate454inter3));
  inv1  gate1755(.a(s_173), .O(gate454inter4));
  nand2 gate1756(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1757(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1758(.a(G1087), .O(gate454inter7));
  inv1  gate1759(.a(G1183), .O(gate454inter8));
  nand2 gate1760(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1761(.a(s_173), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1762(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1763(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1764(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate3067(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate3068(.a(gate455inter0), .b(s_360), .O(gate455inter1));
  and2  gate3069(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate3070(.a(s_360), .O(gate455inter3));
  inv1  gate3071(.a(s_361), .O(gate455inter4));
  nand2 gate3072(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate3073(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate3074(.a(G19), .O(gate455inter7));
  inv1  gate3075(.a(G1186), .O(gate455inter8));
  nand2 gate3076(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate3077(.a(s_361), .b(gate455inter3), .O(gate455inter10));
  nor2  gate3078(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate3079(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate3080(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1009(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1010(.a(gate458inter0), .b(s_66), .O(gate458inter1));
  and2  gate1011(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1012(.a(s_66), .O(gate458inter3));
  inv1  gate1013(.a(s_67), .O(gate458inter4));
  nand2 gate1014(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1015(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1016(.a(G1093), .O(gate458inter7));
  inv1  gate1017(.a(G1189), .O(gate458inter8));
  nand2 gate1018(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1019(.a(s_67), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1020(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1021(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1022(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate2311(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2312(.a(gate459inter0), .b(s_252), .O(gate459inter1));
  and2  gate2313(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2314(.a(s_252), .O(gate459inter3));
  inv1  gate2315(.a(s_253), .O(gate459inter4));
  nand2 gate2316(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2317(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2318(.a(G21), .O(gate459inter7));
  inv1  gate2319(.a(G1192), .O(gate459inter8));
  nand2 gate2320(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2321(.a(s_253), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2322(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2323(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2324(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2829(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2830(.a(gate461inter0), .b(s_326), .O(gate461inter1));
  and2  gate2831(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2832(.a(s_326), .O(gate461inter3));
  inv1  gate2833(.a(s_327), .O(gate461inter4));
  nand2 gate2834(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2835(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2836(.a(G22), .O(gate461inter7));
  inv1  gate2837(.a(G1195), .O(gate461inter8));
  nand2 gate2838(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2839(.a(s_327), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2840(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2841(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2842(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1387(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1388(.a(gate463inter0), .b(s_120), .O(gate463inter1));
  and2  gate1389(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1390(.a(s_120), .O(gate463inter3));
  inv1  gate1391(.a(s_121), .O(gate463inter4));
  nand2 gate1392(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1393(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1394(.a(G23), .O(gate463inter7));
  inv1  gate1395(.a(G1198), .O(gate463inter8));
  nand2 gate1396(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1397(.a(s_121), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1398(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1399(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1400(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1471(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1472(.a(gate467inter0), .b(s_132), .O(gate467inter1));
  and2  gate1473(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1474(.a(s_132), .O(gate467inter3));
  inv1  gate1475(.a(s_133), .O(gate467inter4));
  nand2 gate1476(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1477(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1478(.a(G25), .O(gate467inter7));
  inv1  gate1479(.a(G1204), .O(gate467inter8));
  nand2 gate1480(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1481(.a(s_133), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1482(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1483(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1484(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate2899(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2900(.a(gate468inter0), .b(s_336), .O(gate468inter1));
  and2  gate2901(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2902(.a(s_336), .O(gate468inter3));
  inv1  gate2903(.a(s_337), .O(gate468inter4));
  nand2 gate2904(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2905(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2906(.a(G1108), .O(gate468inter7));
  inv1  gate2907(.a(G1204), .O(gate468inter8));
  nand2 gate2908(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2909(.a(s_337), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2910(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2911(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2912(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate673(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate674(.a(gate471inter0), .b(s_18), .O(gate471inter1));
  and2  gate675(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate676(.a(s_18), .O(gate471inter3));
  inv1  gate677(.a(s_19), .O(gate471inter4));
  nand2 gate678(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate679(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate680(.a(G27), .O(gate471inter7));
  inv1  gate681(.a(G1210), .O(gate471inter8));
  nand2 gate682(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate683(.a(s_19), .b(gate471inter3), .O(gate471inter10));
  nor2  gate684(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate685(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate686(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2059(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2060(.a(gate476inter0), .b(s_216), .O(gate476inter1));
  and2  gate2061(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2062(.a(s_216), .O(gate476inter3));
  inv1  gate2063(.a(s_217), .O(gate476inter4));
  nand2 gate2064(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2065(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2066(.a(G1120), .O(gate476inter7));
  inv1  gate2067(.a(G1216), .O(gate476inter8));
  nand2 gate2068(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2069(.a(s_217), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2070(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2071(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2072(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2843(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2844(.a(gate482inter0), .b(s_328), .O(gate482inter1));
  and2  gate2845(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2846(.a(s_328), .O(gate482inter3));
  inv1  gate2847(.a(s_329), .O(gate482inter4));
  nand2 gate2848(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2849(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2850(.a(G1129), .O(gate482inter7));
  inv1  gate2851(.a(G1225), .O(gate482inter8));
  nand2 gate2852(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2853(.a(s_329), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2854(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2855(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2856(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate687(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate688(.a(gate484inter0), .b(s_20), .O(gate484inter1));
  and2  gate689(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate690(.a(s_20), .O(gate484inter3));
  inv1  gate691(.a(s_21), .O(gate484inter4));
  nand2 gate692(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate693(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate694(.a(G1230), .O(gate484inter7));
  inv1  gate695(.a(G1231), .O(gate484inter8));
  nand2 gate696(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate697(.a(s_21), .b(gate484inter3), .O(gate484inter10));
  nor2  gate698(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate699(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate700(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1345(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1346(.a(gate487inter0), .b(s_114), .O(gate487inter1));
  and2  gate1347(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1348(.a(s_114), .O(gate487inter3));
  inv1  gate1349(.a(s_115), .O(gate487inter4));
  nand2 gate1350(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1351(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1352(.a(G1236), .O(gate487inter7));
  inv1  gate1353(.a(G1237), .O(gate487inter8));
  nand2 gate1354(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1355(.a(s_115), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1356(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1357(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1358(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate715(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate716(.a(gate497inter0), .b(s_24), .O(gate497inter1));
  and2  gate717(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate718(.a(s_24), .O(gate497inter3));
  inv1  gate719(.a(s_25), .O(gate497inter4));
  nand2 gate720(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate721(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate722(.a(G1256), .O(gate497inter7));
  inv1  gate723(.a(G1257), .O(gate497inter8));
  nand2 gate724(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate725(.a(s_25), .b(gate497inter3), .O(gate497inter10));
  nor2  gate726(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate727(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate728(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1989(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1990(.a(gate499inter0), .b(s_206), .O(gate499inter1));
  and2  gate1991(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1992(.a(s_206), .O(gate499inter3));
  inv1  gate1993(.a(s_207), .O(gate499inter4));
  nand2 gate1994(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1995(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1996(.a(G1260), .O(gate499inter7));
  inv1  gate1997(.a(G1261), .O(gate499inter8));
  nand2 gate1998(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1999(.a(s_207), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2000(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2001(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2002(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1135(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1136(.a(gate503inter0), .b(s_84), .O(gate503inter1));
  and2  gate1137(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1138(.a(s_84), .O(gate503inter3));
  inv1  gate1139(.a(s_85), .O(gate503inter4));
  nand2 gate1140(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1141(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1142(.a(G1268), .O(gate503inter7));
  inv1  gate1143(.a(G1269), .O(gate503inter8));
  nand2 gate1144(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1145(.a(s_85), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1146(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1147(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1148(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2045(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2046(.a(gate505inter0), .b(s_214), .O(gate505inter1));
  and2  gate2047(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2048(.a(s_214), .O(gate505inter3));
  inv1  gate2049(.a(s_215), .O(gate505inter4));
  nand2 gate2050(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2051(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2052(.a(G1272), .O(gate505inter7));
  inv1  gate2053(.a(G1273), .O(gate505inter8));
  nand2 gate2054(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2055(.a(s_215), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2056(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2057(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2058(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate2073(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2074(.a(gate506inter0), .b(s_218), .O(gate506inter1));
  and2  gate2075(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2076(.a(s_218), .O(gate506inter3));
  inv1  gate2077(.a(s_219), .O(gate506inter4));
  nand2 gate2078(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2079(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2080(.a(G1274), .O(gate506inter7));
  inv1  gate2081(.a(G1275), .O(gate506inter8));
  nand2 gate2082(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2083(.a(s_219), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2084(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2085(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2086(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1933(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1934(.a(gate509inter0), .b(s_198), .O(gate509inter1));
  and2  gate1935(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1936(.a(s_198), .O(gate509inter3));
  inv1  gate1937(.a(s_199), .O(gate509inter4));
  nand2 gate1938(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1939(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1940(.a(G1280), .O(gate509inter7));
  inv1  gate1941(.a(G1281), .O(gate509inter8));
  nand2 gate1942(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1943(.a(s_199), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1944(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1945(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1946(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1429(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1430(.a(gate512inter0), .b(s_126), .O(gate512inter1));
  and2  gate1431(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1432(.a(s_126), .O(gate512inter3));
  inv1  gate1433(.a(s_127), .O(gate512inter4));
  nand2 gate1434(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1435(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1436(.a(G1286), .O(gate512inter7));
  inv1  gate1437(.a(G1287), .O(gate512inter8));
  nand2 gate1438(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1439(.a(s_127), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1440(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1441(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1442(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1331(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1332(.a(gate513inter0), .b(s_112), .O(gate513inter1));
  and2  gate1333(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1334(.a(s_112), .O(gate513inter3));
  inv1  gate1335(.a(s_113), .O(gate513inter4));
  nand2 gate1336(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1337(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1338(.a(G1288), .O(gate513inter7));
  inv1  gate1339(.a(G1289), .O(gate513inter8));
  nand2 gate1340(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1341(.a(s_113), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1342(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1343(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1344(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1597(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1598(.a(gate514inter0), .b(s_150), .O(gate514inter1));
  and2  gate1599(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1600(.a(s_150), .O(gate514inter3));
  inv1  gate1601(.a(s_151), .O(gate514inter4));
  nand2 gate1602(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1603(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1604(.a(G1290), .O(gate514inter7));
  inv1  gate1605(.a(G1291), .O(gate514inter8));
  nand2 gate1606(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1607(.a(s_151), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1608(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1609(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1610(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule