module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate701(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate702(.a(gate10inter0), .b(s_22), .O(gate10inter1));
  and2  gate703(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate704(.a(s_22), .O(gate10inter3));
  inv1  gate705(.a(s_23), .O(gate10inter4));
  nand2 gate706(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate707(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate708(.a(G3), .O(gate10inter7));
  inv1  gate709(.a(G4), .O(gate10inter8));
  nand2 gate710(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate711(.a(s_23), .b(gate10inter3), .O(gate10inter10));
  nor2  gate712(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate713(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate714(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate897(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate898(.a(gate11inter0), .b(s_50), .O(gate11inter1));
  and2  gate899(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate900(.a(s_50), .O(gate11inter3));
  inv1  gate901(.a(s_51), .O(gate11inter4));
  nand2 gate902(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate903(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate904(.a(G5), .O(gate11inter7));
  inv1  gate905(.a(G6), .O(gate11inter8));
  nand2 gate906(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate907(.a(s_51), .b(gate11inter3), .O(gate11inter10));
  nor2  gate908(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate909(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate910(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1667(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1668(.a(gate12inter0), .b(s_160), .O(gate12inter1));
  and2  gate1669(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1670(.a(s_160), .O(gate12inter3));
  inv1  gate1671(.a(s_161), .O(gate12inter4));
  nand2 gate1672(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1673(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1674(.a(G7), .O(gate12inter7));
  inv1  gate1675(.a(G8), .O(gate12inter8));
  nand2 gate1676(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1677(.a(s_161), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1678(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1679(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1680(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate771(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate772(.a(gate14inter0), .b(s_32), .O(gate14inter1));
  and2  gate773(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate774(.a(s_32), .O(gate14inter3));
  inv1  gate775(.a(s_33), .O(gate14inter4));
  nand2 gate776(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate777(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate778(.a(G11), .O(gate14inter7));
  inv1  gate779(.a(G12), .O(gate14inter8));
  nand2 gate780(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate781(.a(s_33), .b(gate14inter3), .O(gate14inter10));
  nor2  gate782(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate783(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate784(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate785(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate786(.a(gate26inter0), .b(s_34), .O(gate26inter1));
  and2  gate787(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate788(.a(s_34), .O(gate26inter3));
  inv1  gate789(.a(s_35), .O(gate26inter4));
  nand2 gate790(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate791(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate792(.a(G9), .O(gate26inter7));
  inv1  gate793(.a(G13), .O(gate26inter8));
  nand2 gate794(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate795(.a(s_35), .b(gate26inter3), .O(gate26inter10));
  nor2  gate796(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate797(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate798(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate1149(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1150(.a(gate27inter0), .b(s_86), .O(gate27inter1));
  and2  gate1151(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1152(.a(s_86), .O(gate27inter3));
  inv1  gate1153(.a(s_87), .O(gate27inter4));
  nand2 gate1154(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1155(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1156(.a(G2), .O(gate27inter7));
  inv1  gate1157(.a(G6), .O(gate27inter8));
  nand2 gate1158(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1159(.a(s_87), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1160(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1161(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1162(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate995(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate996(.a(gate29inter0), .b(s_64), .O(gate29inter1));
  and2  gate997(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate998(.a(s_64), .O(gate29inter3));
  inv1  gate999(.a(s_65), .O(gate29inter4));
  nand2 gate1000(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1001(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1002(.a(G3), .O(gate29inter7));
  inv1  gate1003(.a(G7), .O(gate29inter8));
  nand2 gate1004(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1005(.a(s_65), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1006(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1007(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1008(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1107(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1108(.a(gate30inter0), .b(s_80), .O(gate30inter1));
  and2  gate1109(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1110(.a(s_80), .O(gate30inter3));
  inv1  gate1111(.a(s_81), .O(gate30inter4));
  nand2 gate1112(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1113(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1114(.a(G11), .O(gate30inter7));
  inv1  gate1115(.a(G15), .O(gate30inter8));
  nand2 gate1116(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1117(.a(s_81), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1118(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1119(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1120(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1093(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1094(.a(gate33inter0), .b(s_78), .O(gate33inter1));
  and2  gate1095(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1096(.a(s_78), .O(gate33inter3));
  inv1  gate1097(.a(s_79), .O(gate33inter4));
  nand2 gate1098(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1099(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1100(.a(G17), .O(gate33inter7));
  inv1  gate1101(.a(G21), .O(gate33inter8));
  nand2 gate1102(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1103(.a(s_79), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1104(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1105(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1106(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1079(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1080(.a(gate34inter0), .b(s_76), .O(gate34inter1));
  and2  gate1081(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1082(.a(s_76), .O(gate34inter3));
  inv1  gate1083(.a(s_77), .O(gate34inter4));
  nand2 gate1084(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1085(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1086(.a(G25), .O(gate34inter7));
  inv1  gate1087(.a(G29), .O(gate34inter8));
  nand2 gate1088(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1089(.a(s_77), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1090(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1091(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1092(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate855(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate856(.a(gate41inter0), .b(s_44), .O(gate41inter1));
  and2  gate857(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate858(.a(s_44), .O(gate41inter3));
  inv1  gate859(.a(s_45), .O(gate41inter4));
  nand2 gate860(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate861(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate862(.a(G1), .O(gate41inter7));
  inv1  gate863(.a(G266), .O(gate41inter8));
  nand2 gate864(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate865(.a(s_45), .b(gate41inter3), .O(gate41inter10));
  nor2  gate866(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate867(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate868(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate631(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate632(.a(gate66inter0), .b(s_12), .O(gate66inter1));
  and2  gate633(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate634(.a(s_12), .O(gate66inter3));
  inv1  gate635(.a(s_13), .O(gate66inter4));
  nand2 gate636(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate637(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate638(.a(G26), .O(gate66inter7));
  inv1  gate639(.a(G302), .O(gate66inter8));
  nand2 gate640(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate641(.a(s_13), .b(gate66inter3), .O(gate66inter10));
  nor2  gate642(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate643(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate644(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1429(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1430(.a(gate67inter0), .b(s_126), .O(gate67inter1));
  and2  gate1431(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1432(.a(s_126), .O(gate67inter3));
  inv1  gate1433(.a(s_127), .O(gate67inter4));
  nand2 gate1434(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1435(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1436(.a(G27), .O(gate67inter7));
  inv1  gate1437(.a(G305), .O(gate67inter8));
  nand2 gate1438(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1439(.a(s_127), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1440(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1441(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1442(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate911(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate912(.a(gate74inter0), .b(s_52), .O(gate74inter1));
  and2  gate913(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate914(.a(s_52), .O(gate74inter3));
  inv1  gate915(.a(s_53), .O(gate74inter4));
  nand2 gate916(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate917(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate918(.a(G5), .O(gate74inter7));
  inv1  gate919(.a(G314), .O(gate74inter8));
  nand2 gate920(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate921(.a(s_53), .b(gate74inter3), .O(gate74inter10));
  nor2  gate922(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate923(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate924(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1443(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1444(.a(gate75inter0), .b(s_128), .O(gate75inter1));
  and2  gate1445(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1446(.a(s_128), .O(gate75inter3));
  inv1  gate1447(.a(s_129), .O(gate75inter4));
  nand2 gate1448(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1449(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1450(.a(G9), .O(gate75inter7));
  inv1  gate1451(.a(G317), .O(gate75inter8));
  nand2 gate1452(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1453(.a(s_129), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1454(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1455(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1456(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate743(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate744(.a(gate80inter0), .b(s_28), .O(gate80inter1));
  and2  gate745(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate746(.a(s_28), .O(gate80inter3));
  inv1  gate747(.a(s_29), .O(gate80inter4));
  nand2 gate748(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate749(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate750(.a(G14), .O(gate80inter7));
  inv1  gate751(.a(G323), .O(gate80inter8));
  nand2 gate752(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate753(.a(s_29), .b(gate80inter3), .O(gate80inter10));
  nor2  gate754(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate755(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate756(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate659(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate660(.a(gate84inter0), .b(s_16), .O(gate84inter1));
  and2  gate661(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate662(.a(s_16), .O(gate84inter3));
  inv1  gate663(.a(s_17), .O(gate84inter4));
  nand2 gate664(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate665(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate666(.a(G15), .O(gate84inter7));
  inv1  gate667(.a(G329), .O(gate84inter8));
  nand2 gate668(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate669(.a(s_17), .b(gate84inter3), .O(gate84inter10));
  nor2  gate670(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate671(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate672(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1261(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1262(.a(gate89inter0), .b(s_102), .O(gate89inter1));
  and2  gate1263(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1264(.a(s_102), .O(gate89inter3));
  inv1  gate1265(.a(s_103), .O(gate89inter4));
  nand2 gate1266(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1267(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1268(.a(G17), .O(gate89inter7));
  inv1  gate1269(.a(G338), .O(gate89inter8));
  nand2 gate1270(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1271(.a(s_103), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1272(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1273(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1274(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1247(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1248(.a(gate98inter0), .b(s_100), .O(gate98inter1));
  and2  gate1249(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1250(.a(s_100), .O(gate98inter3));
  inv1  gate1251(.a(s_101), .O(gate98inter4));
  nand2 gate1252(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1253(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1254(.a(G23), .O(gate98inter7));
  inv1  gate1255(.a(G350), .O(gate98inter8));
  nand2 gate1256(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1257(.a(s_101), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1258(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1259(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1260(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1583(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1584(.a(gate99inter0), .b(s_148), .O(gate99inter1));
  and2  gate1585(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1586(.a(s_148), .O(gate99inter3));
  inv1  gate1587(.a(s_149), .O(gate99inter4));
  nand2 gate1588(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1589(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1590(.a(G27), .O(gate99inter7));
  inv1  gate1591(.a(G353), .O(gate99inter8));
  nand2 gate1592(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1593(.a(s_149), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1594(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1595(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1596(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate939(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate940(.a(gate108inter0), .b(s_56), .O(gate108inter1));
  and2  gate941(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate942(.a(s_56), .O(gate108inter3));
  inv1  gate943(.a(s_57), .O(gate108inter4));
  nand2 gate944(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate945(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate946(.a(G368), .O(gate108inter7));
  inv1  gate947(.a(G369), .O(gate108inter8));
  nand2 gate948(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate949(.a(s_57), .b(gate108inter3), .O(gate108inter10));
  nor2  gate950(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate951(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate952(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1345(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1346(.a(gate115inter0), .b(s_114), .O(gate115inter1));
  and2  gate1347(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1348(.a(s_114), .O(gate115inter3));
  inv1  gate1349(.a(s_115), .O(gate115inter4));
  nand2 gate1350(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1351(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1352(.a(G382), .O(gate115inter7));
  inv1  gate1353(.a(G383), .O(gate115inter8));
  nand2 gate1354(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1355(.a(s_115), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1356(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1357(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1358(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1373(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1374(.a(gate116inter0), .b(s_118), .O(gate116inter1));
  and2  gate1375(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1376(.a(s_118), .O(gate116inter3));
  inv1  gate1377(.a(s_119), .O(gate116inter4));
  nand2 gate1378(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1379(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1380(.a(G384), .O(gate116inter7));
  inv1  gate1381(.a(G385), .O(gate116inter8));
  nand2 gate1382(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1383(.a(s_119), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1384(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1385(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1386(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate883(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate884(.a(gate145inter0), .b(s_48), .O(gate145inter1));
  and2  gate885(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate886(.a(s_48), .O(gate145inter3));
  inv1  gate887(.a(s_49), .O(gate145inter4));
  nand2 gate888(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate889(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate890(.a(G474), .O(gate145inter7));
  inv1  gate891(.a(G477), .O(gate145inter8));
  nand2 gate892(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate893(.a(s_49), .b(gate145inter3), .O(gate145inter10));
  nor2  gate894(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate895(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate896(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate729(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate730(.a(gate150inter0), .b(s_26), .O(gate150inter1));
  and2  gate731(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate732(.a(s_26), .O(gate150inter3));
  inv1  gate733(.a(s_27), .O(gate150inter4));
  nand2 gate734(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate735(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate736(.a(G504), .O(gate150inter7));
  inv1  gate737(.a(G507), .O(gate150inter8));
  nand2 gate738(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate739(.a(s_27), .b(gate150inter3), .O(gate150inter10));
  nor2  gate740(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate741(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate742(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate575(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate576(.a(gate155inter0), .b(s_4), .O(gate155inter1));
  and2  gate577(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate578(.a(s_4), .O(gate155inter3));
  inv1  gate579(.a(s_5), .O(gate155inter4));
  nand2 gate580(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate581(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate582(.a(G432), .O(gate155inter7));
  inv1  gate583(.a(G525), .O(gate155inter8));
  nand2 gate584(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate585(.a(s_5), .b(gate155inter3), .O(gate155inter10));
  nor2  gate586(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate587(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate588(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1331(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1332(.a(gate172inter0), .b(s_112), .O(gate172inter1));
  and2  gate1333(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1334(.a(s_112), .O(gate172inter3));
  inv1  gate1335(.a(s_113), .O(gate172inter4));
  nand2 gate1336(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1337(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1338(.a(G483), .O(gate172inter7));
  inv1  gate1339(.a(G549), .O(gate172inter8));
  nand2 gate1340(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1341(.a(s_113), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1342(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1343(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1344(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1135(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1136(.a(gate183inter0), .b(s_84), .O(gate183inter1));
  and2  gate1137(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1138(.a(s_84), .O(gate183inter3));
  inv1  gate1139(.a(s_85), .O(gate183inter4));
  nand2 gate1140(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1141(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1142(.a(G516), .O(gate183inter7));
  inv1  gate1143(.a(G567), .O(gate183inter8));
  nand2 gate1144(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1145(.a(s_85), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1146(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1147(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1148(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1191(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1192(.a(gate184inter0), .b(s_92), .O(gate184inter1));
  and2  gate1193(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1194(.a(s_92), .O(gate184inter3));
  inv1  gate1195(.a(s_93), .O(gate184inter4));
  nand2 gate1196(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1197(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1198(.a(G519), .O(gate184inter7));
  inv1  gate1199(.a(G567), .O(gate184inter8));
  nand2 gate1200(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1201(.a(s_93), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1202(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1203(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1204(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1471(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1472(.a(gate185inter0), .b(s_132), .O(gate185inter1));
  and2  gate1473(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1474(.a(s_132), .O(gate185inter3));
  inv1  gate1475(.a(s_133), .O(gate185inter4));
  nand2 gate1476(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1477(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1478(.a(G570), .O(gate185inter7));
  inv1  gate1479(.a(G571), .O(gate185inter8));
  nand2 gate1480(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1481(.a(s_133), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1482(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1483(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1484(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate589(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate590(.a(gate187inter0), .b(s_6), .O(gate187inter1));
  and2  gate591(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate592(.a(s_6), .O(gate187inter3));
  inv1  gate593(.a(s_7), .O(gate187inter4));
  nand2 gate594(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate595(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate596(.a(G574), .O(gate187inter7));
  inv1  gate597(.a(G575), .O(gate187inter8));
  nand2 gate598(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate599(.a(s_7), .b(gate187inter3), .O(gate187inter10));
  nor2  gate600(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate601(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate602(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate953(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate954(.a(gate190inter0), .b(s_58), .O(gate190inter1));
  and2  gate955(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate956(.a(s_58), .O(gate190inter3));
  inv1  gate957(.a(s_59), .O(gate190inter4));
  nand2 gate958(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate959(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate960(.a(G580), .O(gate190inter7));
  inv1  gate961(.a(G581), .O(gate190inter8));
  nand2 gate962(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate963(.a(s_59), .b(gate190inter3), .O(gate190inter10));
  nor2  gate964(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate965(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate966(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1317(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1318(.a(gate196inter0), .b(s_110), .O(gate196inter1));
  and2  gate1319(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1320(.a(s_110), .O(gate196inter3));
  inv1  gate1321(.a(s_111), .O(gate196inter4));
  nand2 gate1322(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1323(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1324(.a(G592), .O(gate196inter7));
  inv1  gate1325(.a(G593), .O(gate196inter8));
  nand2 gate1326(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1327(.a(s_111), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1328(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1329(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1330(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate617(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate618(.a(gate200inter0), .b(s_10), .O(gate200inter1));
  and2  gate619(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate620(.a(s_10), .O(gate200inter3));
  inv1  gate621(.a(s_11), .O(gate200inter4));
  nand2 gate622(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate623(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate624(.a(G600), .O(gate200inter7));
  inv1  gate625(.a(G601), .O(gate200inter8));
  nand2 gate626(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate627(.a(s_11), .b(gate200inter3), .O(gate200inter10));
  nor2  gate628(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate629(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate630(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1387(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1388(.a(gate213inter0), .b(s_120), .O(gate213inter1));
  and2  gate1389(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1390(.a(s_120), .O(gate213inter3));
  inv1  gate1391(.a(s_121), .O(gate213inter4));
  nand2 gate1392(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1393(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1394(.a(G602), .O(gate213inter7));
  inv1  gate1395(.a(G672), .O(gate213inter8));
  nand2 gate1396(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1397(.a(s_121), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1398(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1399(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1400(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1121(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1122(.a(gate215inter0), .b(s_82), .O(gate215inter1));
  and2  gate1123(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1124(.a(s_82), .O(gate215inter3));
  inv1  gate1125(.a(s_83), .O(gate215inter4));
  nand2 gate1126(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1127(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1128(.a(G607), .O(gate215inter7));
  inv1  gate1129(.a(G675), .O(gate215inter8));
  nand2 gate1130(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1131(.a(s_83), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1132(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1133(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1134(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1219(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1220(.a(gate234inter0), .b(s_96), .O(gate234inter1));
  and2  gate1221(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1222(.a(s_96), .O(gate234inter3));
  inv1  gate1223(.a(s_97), .O(gate234inter4));
  nand2 gate1224(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1225(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1226(.a(G245), .O(gate234inter7));
  inv1  gate1227(.a(G721), .O(gate234inter8));
  nand2 gate1228(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1229(.a(s_97), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1230(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1231(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1232(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1555(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1556(.a(gate237inter0), .b(s_144), .O(gate237inter1));
  and2  gate1557(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1558(.a(s_144), .O(gate237inter3));
  inv1  gate1559(.a(s_145), .O(gate237inter4));
  nand2 gate1560(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1561(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1562(.a(G254), .O(gate237inter7));
  inv1  gate1563(.a(G706), .O(gate237inter8));
  nand2 gate1564(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1565(.a(s_145), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1566(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1567(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1568(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1485(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1486(.a(gate241inter0), .b(s_134), .O(gate241inter1));
  and2  gate1487(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1488(.a(s_134), .O(gate241inter3));
  inv1  gate1489(.a(s_135), .O(gate241inter4));
  nand2 gate1490(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1491(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1492(.a(G242), .O(gate241inter7));
  inv1  gate1493(.a(G730), .O(gate241inter8));
  nand2 gate1494(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1495(.a(s_135), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1496(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1497(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1498(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1065(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1066(.a(gate243inter0), .b(s_74), .O(gate243inter1));
  and2  gate1067(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1068(.a(s_74), .O(gate243inter3));
  inv1  gate1069(.a(s_75), .O(gate243inter4));
  nand2 gate1070(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1071(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1072(.a(G245), .O(gate243inter7));
  inv1  gate1073(.a(G733), .O(gate243inter8));
  nand2 gate1074(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1075(.a(s_75), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1076(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1077(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1078(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1611(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1612(.a(gate247inter0), .b(s_152), .O(gate247inter1));
  and2  gate1613(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1614(.a(s_152), .O(gate247inter3));
  inv1  gate1615(.a(s_153), .O(gate247inter4));
  nand2 gate1616(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1617(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1618(.a(G251), .O(gate247inter7));
  inv1  gate1619(.a(G739), .O(gate247inter8));
  nand2 gate1620(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1621(.a(s_153), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1622(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1623(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1624(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1569(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1570(.a(gate251inter0), .b(s_146), .O(gate251inter1));
  and2  gate1571(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1572(.a(s_146), .O(gate251inter3));
  inv1  gate1573(.a(s_147), .O(gate251inter4));
  nand2 gate1574(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1575(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1576(.a(G257), .O(gate251inter7));
  inv1  gate1577(.a(G745), .O(gate251inter8));
  nand2 gate1578(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1579(.a(s_147), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1580(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1581(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1582(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate925(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate926(.a(gate253inter0), .b(s_54), .O(gate253inter1));
  and2  gate927(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate928(.a(s_54), .O(gate253inter3));
  inv1  gate929(.a(s_55), .O(gate253inter4));
  nand2 gate930(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate931(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate932(.a(G260), .O(gate253inter7));
  inv1  gate933(.a(G748), .O(gate253inter8));
  nand2 gate934(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate935(.a(s_55), .b(gate253inter3), .O(gate253inter10));
  nor2  gate936(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate937(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate938(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1359(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1360(.a(gate254inter0), .b(s_116), .O(gate254inter1));
  and2  gate1361(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1362(.a(s_116), .O(gate254inter3));
  inv1  gate1363(.a(s_117), .O(gate254inter4));
  nand2 gate1364(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1365(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1366(.a(G712), .O(gate254inter7));
  inv1  gate1367(.a(G748), .O(gate254inter8));
  nand2 gate1368(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1369(.a(s_117), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1370(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1371(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1372(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate981(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate982(.a(gate255inter0), .b(s_62), .O(gate255inter1));
  and2  gate983(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate984(.a(s_62), .O(gate255inter3));
  inv1  gate985(.a(s_63), .O(gate255inter4));
  nand2 gate986(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate987(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate988(.a(G263), .O(gate255inter7));
  inv1  gate989(.a(G751), .O(gate255inter8));
  nand2 gate990(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate991(.a(s_63), .b(gate255inter3), .O(gate255inter10));
  nor2  gate992(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate993(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate994(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1163(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1164(.a(gate256inter0), .b(s_88), .O(gate256inter1));
  and2  gate1165(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1166(.a(s_88), .O(gate256inter3));
  inv1  gate1167(.a(s_89), .O(gate256inter4));
  nand2 gate1168(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1169(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1170(.a(G715), .O(gate256inter7));
  inv1  gate1171(.a(G751), .O(gate256inter8));
  nand2 gate1172(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1173(.a(s_89), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1174(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1175(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1176(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1233(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1234(.a(gate258inter0), .b(s_98), .O(gate258inter1));
  and2  gate1235(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1236(.a(s_98), .O(gate258inter3));
  inv1  gate1237(.a(s_99), .O(gate258inter4));
  nand2 gate1238(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1239(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1240(.a(G756), .O(gate258inter7));
  inv1  gate1241(.a(G757), .O(gate258inter8));
  nand2 gate1242(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1243(.a(s_99), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1244(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1245(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1246(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1653(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1654(.a(gate268inter0), .b(s_158), .O(gate268inter1));
  and2  gate1655(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1656(.a(s_158), .O(gate268inter3));
  inv1  gate1657(.a(s_159), .O(gate268inter4));
  nand2 gate1658(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1659(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1660(.a(G651), .O(gate268inter7));
  inv1  gate1661(.a(G779), .O(gate268inter8));
  nand2 gate1662(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1663(.a(s_159), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1664(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1665(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1666(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate841(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate842(.a(gate271inter0), .b(s_42), .O(gate271inter1));
  and2  gate843(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate844(.a(s_42), .O(gate271inter3));
  inv1  gate845(.a(s_43), .O(gate271inter4));
  nand2 gate846(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate847(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate848(.a(G660), .O(gate271inter7));
  inv1  gate849(.a(G788), .O(gate271inter8));
  nand2 gate850(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate851(.a(s_43), .b(gate271inter3), .O(gate271inter10));
  nor2  gate852(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate853(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate854(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate673(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate674(.a(gate274inter0), .b(s_18), .O(gate274inter1));
  and2  gate675(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate676(.a(s_18), .O(gate274inter3));
  inv1  gate677(.a(s_19), .O(gate274inter4));
  nand2 gate678(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate679(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate680(.a(G770), .O(gate274inter7));
  inv1  gate681(.a(G794), .O(gate274inter8));
  nand2 gate682(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate683(.a(s_19), .b(gate274inter3), .O(gate274inter10));
  nor2  gate684(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate685(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate686(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1177(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1178(.a(gate279inter0), .b(s_90), .O(gate279inter1));
  and2  gate1179(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1180(.a(s_90), .O(gate279inter3));
  inv1  gate1181(.a(s_91), .O(gate279inter4));
  nand2 gate1182(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1183(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1184(.a(G651), .O(gate279inter7));
  inv1  gate1185(.a(G803), .O(gate279inter8));
  nand2 gate1186(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1187(.a(s_91), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1188(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1189(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1190(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1625(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1626(.a(gate285inter0), .b(s_154), .O(gate285inter1));
  and2  gate1627(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1628(.a(s_154), .O(gate285inter3));
  inv1  gate1629(.a(s_155), .O(gate285inter4));
  nand2 gate1630(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1631(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1632(.a(G660), .O(gate285inter7));
  inv1  gate1633(.a(G812), .O(gate285inter8));
  nand2 gate1634(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1635(.a(s_155), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1636(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1637(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1638(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1275(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1276(.a(gate292inter0), .b(s_104), .O(gate292inter1));
  and2  gate1277(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1278(.a(s_104), .O(gate292inter3));
  inv1  gate1279(.a(s_105), .O(gate292inter4));
  nand2 gate1280(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1281(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1282(.a(G824), .O(gate292inter7));
  inv1  gate1283(.a(G825), .O(gate292inter8));
  nand2 gate1284(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1285(.a(s_105), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1286(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1287(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1288(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1037(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1038(.a(gate295inter0), .b(s_70), .O(gate295inter1));
  and2  gate1039(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1040(.a(s_70), .O(gate295inter3));
  inv1  gate1041(.a(s_71), .O(gate295inter4));
  nand2 gate1042(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1043(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1044(.a(G830), .O(gate295inter7));
  inv1  gate1045(.a(G831), .O(gate295inter8));
  nand2 gate1046(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1047(.a(s_71), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1048(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1049(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1050(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1639(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1640(.a(gate392inter0), .b(s_156), .O(gate392inter1));
  and2  gate1641(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1642(.a(s_156), .O(gate392inter3));
  inv1  gate1643(.a(s_157), .O(gate392inter4));
  nand2 gate1644(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1645(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1646(.a(G6), .O(gate392inter7));
  inv1  gate1647(.a(G1051), .O(gate392inter8));
  nand2 gate1648(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1649(.a(s_157), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1650(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1651(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1652(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1303(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1304(.a(gate393inter0), .b(s_108), .O(gate393inter1));
  and2  gate1305(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1306(.a(s_108), .O(gate393inter3));
  inv1  gate1307(.a(s_109), .O(gate393inter4));
  nand2 gate1308(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1309(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1310(.a(G7), .O(gate393inter7));
  inv1  gate1311(.a(G1054), .O(gate393inter8));
  nand2 gate1312(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1313(.a(s_109), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1314(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1315(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1316(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1051(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1052(.a(gate402inter0), .b(s_72), .O(gate402inter1));
  and2  gate1053(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1054(.a(s_72), .O(gate402inter3));
  inv1  gate1055(.a(s_73), .O(gate402inter4));
  nand2 gate1056(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1057(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1058(.a(G16), .O(gate402inter7));
  inv1  gate1059(.a(G1081), .O(gate402inter8));
  nand2 gate1060(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1061(.a(s_73), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1062(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1063(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1064(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1597(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1598(.a(gate404inter0), .b(s_150), .O(gate404inter1));
  and2  gate1599(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1600(.a(s_150), .O(gate404inter3));
  inv1  gate1601(.a(s_151), .O(gate404inter4));
  nand2 gate1602(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1603(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1604(.a(G18), .O(gate404inter7));
  inv1  gate1605(.a(G1087), .O(gate404inter8));
  nand2 gate1606(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1607(.a(s_151), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1608(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1609(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1610(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate757(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate758(.a(gate407inter0), .b(s_30), .O(gate407inter1));
  and2  gate759(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate760(.a(s_30), .O(gate407inter3));
  inv1  gate761(.a(s_31), .O(gate407inter4));
  nand2 gate762(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate763(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate764(.a(G21), .O(gate407inter7));
  inv1  gate765(.a(G1096), .O(gate407inter8));
  nand2 gate766(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate767(.a(s_31), .b(gate407inter3), .O(gate407inter10));
  nor2  gate768(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate769(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate770(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1527(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1528(.a(gate408inter0), .b(s_140), .O(gate408inter1));
  and2  gate1529(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1530(.a(s_140), .O(gate408inter3));
  inv1  gate1531(.a(s_141), .O(gate408inter4));
  nand2 gate1532(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1533(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1534(.a(G22), .O(gate408inter7));
  inv1  gate1535(.a(G1099), .O(gate408inter8));
  nand2 gate1536(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1537(.a(s_141), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1538(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1539(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1540(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate715(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate716(.a(gate410inter0), .b(s_24), .O(gate410inter1));
  and2  gate717(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate718(.a(s_24), .O(gate410inter3));
  inv1  gate719(.a(s_25), .O(gate410inter4));
  nand2 gate720(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate721(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate722(.a(G24), .O(gate410inter7));
  inv1  gate723(.a(G1105), .O(gate410inter8));
  nand2 gate724(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate725(.a(s_25), .b(gate410inter3), .O(gate410inter10));
  nor2  gate726(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate727(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate728(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1401(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1402(.a(gate419inter0), .b(s_122), .O(gate419inter1));
  and2  gate1403(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1404(.a(s_122), .O(gate419inter3));
  inv1  gate1405(.a(s_123), .O(gate419inter4));
  nand2 gate1406(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1407(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1408(.a(G1), .O(gate419inter7));
  inv1  gate1409(.a(G1132), .O(gate419inter8));
  nand2 gate1410(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1411(.a(s_123), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1412(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1413(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1414(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1205(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1206(.a(gate430inter0), .b(s_94), .O(gate430inter1));
  and2  gate1207(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1208(.a(s_94), .O(gate430inter3));
  inv1  gate1209(.a(s_95), .O(gate430inter4));
  nand2 gate1210(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1211(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1212(.a(G1051), .O(gate430inter7));
  inv1  gate1213(.a(G1147), .O(gate430inter8));
  nand2 gate1214(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1215(.a(s_95), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1216(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1217(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1218(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1541(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1542(.a(gate433inter0), .b(s_142), .O(gate433inter1));
  and2  gate1543(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1544(.a(s_142), .O(gate433inter3));
  inv1  gate1545(.a(s_143), .O(gate433inter4));
  nand2 gate1546(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1547(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1548(.a(G8), .O(gate433inter7));
  inv1  gate1549(.a(G1153), .O(gate433inter8));
  nand2 gate1550(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1551(.a(s_143), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1552(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1553(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1554(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate799(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate800(.a(gate436inter0), .b(s_36), .O(gate436inter1));
  and2  gate801(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate802(.a(s_36), .O(gate436inter3));
  inv1  gate803(.a(s_37), .O(gate436inter4));
  nand2 gate804(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate805(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate806(.a(G1060), .O(gate436inter7));
  inv1  gate807(.a(G1156), .O(gate436inter8));
  nand2 gate808(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate809(.a(s_37), .b(gate436inter3), .O(gate436inter10));
  nor2  gate810(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate811(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate812(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1499(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1500(.a(gate438inter0), .b(s_136), .O(gate438inter1));
  and2  gate1501(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1502(.a(s_136), .O(gate438inter3));
  inv1  gate1503(.a(s_137), .O(gate438inter4));
  nand2 gate1504(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1505(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1506(.a(G1063), .O(gate438inter7));
  inv1  gate1507(.a(G1159), .O(gate438inter8));
  nand2 gate1508(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1509(.a(s_137), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1510(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1511(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1512(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate967(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate968(.a(gate444inter0), .b(s_60), .O(gate444inter1));
  and2  gate969(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate970(.a(s_60), .O(gate444inter3));
  inv1  gate971(.a(s_61), .O(gate444inter4));
  nand2 gate972(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate973(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate974(.a(G1072), .O(gate444inter7));
  inv1  gate975(.a(G1168), .O(gate444inter8));
  nand2 gate976(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate977(.a(s_61), .b(gate444inter3), .O(gate444inter10));
  nor2  gate978(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate979(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate980(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate645(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate646(.a(gate449inter0), .b(s_14), .O(gate449inter1));
  and2  gate647(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate648(.a(s_14), .O(gate449inter3));
  inv1  gate649(.a(s_15), .O(gate449inter4));
  nand2 gate650(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate651(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate652(.a(G16), .O(gate449inter7));
  inv1  gate653(.a(G1177), .O(gate449inter8));
  nand2 gate654(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate655(.a(s_15), .b(gate449inter3), .O(gate449inter10));
  nor2  gate656(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate657(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate658(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1415(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1416(.a(gate456inter0), .b(s_124), .O(gate456inter1));
  and2  gate1417(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1418(.a(s_124), .O(gate456inter3));
  inv1  gate1419(.a(s_125), .O(gate456inter4));
  nand2 gate1420(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1421(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1422(.a(G1090), .O(gate456inter7));
  inv1  gate1423(.a(G1186), .O(gate456inter8));
  nand2 gate1424(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1425(.a(s_125), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1426(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1427(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1428(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate687(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate688(.a(gate471inter0), .b(s_20), .O(gate471inter1));
  and2  gate689(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate690(.a(s_20), .O(gate471inter3));
  inv1  gate691(.a(s_21), .O(gate471inter4));
  nand2 gate692(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate693(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate694(.a(G27), .O(gate471inter7));
  inv1  gate695(.a(G1210), .O(gate471inter8));
  nand2 gate696(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate697(.a(s_21), .b(gate471inter3), .O(gate471inter10));
  nor2  gate698(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate699(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate700(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate547(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate548(.a(gate474inter0), .b(s_0), .O(gate474inter1));
  and2  gate549(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate550(.a(s_0), .O(gate474inter3));
  inv1  gate551(.a(s_1), .O(gate474inter4));
  nand2 gate552(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate553(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate554(.a(G1117), .O(gate474inter7));
  inv1  gate555(.a(G1213), .O(gate474inter8));
  nand2 gate556(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate557(.a(s_1), .b(gate474inter3), .O(gate474inter10));
  nor2  gate558(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate559(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate560(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate561(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate562(.a(gate478inter0), .b(s_2), .O(gate478inter1));
  and2  gate563(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate564(.a(s_2), .O(gate478inter3));
  inv1  gate565(.a(s_3), .O(gate478inter4));
  nand2 gate566(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate567(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate568(.a(G1123), .O(gate478inter7));
  inv1  gate569(.a(G1219), .O(gate478inter8));
  nand2 gate570(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate571(.a(s_3), .b(gate478inter3), .O(gate478inter10));
  nor2  gate572(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate573(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate574(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1009(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1010(.a(gate481inter0), .b(s_66), .O(gate481inter1));
  and2  gate1011(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1012(.a(s_66), .O(gate481inter3));
  inv1  gate1013(.a(s_67), .O(gate481inter4));
  nand2 gate1014(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1015(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1016(.a(G32), .O(gate481inter7));
  inv1  gate1017(.a(G1225), .O(gate481inter8));
  nand2 gate1018(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1019(.a(s_67), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1020(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1021(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1022(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1289(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1290(.a(gate483inter0), .b(s_106), .O(gate483inter1));
  and2  gate1291(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1292(.a(s_106), .O(gate483inter3));
  inv1  gate1293(.a(s_107), .O(gate483inter4));
  nand2 gate1294(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1295(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1296(.a(G1228), .O(gate483inter7));
  inv1  gate1297(.a(G1229), .O(gate483inter8));
  nand2 gate1298(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1299(.a(s_107), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1300(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1301(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1302(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate827(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate828(.a(gate494inter0), .b(s_40), .O(gate494inter1));
  and2  gate829(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate830(.a(s_40), .O(gate494inter3));
  inv1  gate831(.a(s_41), .O(gate494inter4));
  nand2 gate832(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate833(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate834(.a(G1250), .O(gate494inter7));
  inv1  gate835(.a(G1251), .O(gate494inter8));
  nand2 gate836(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate837(.a(s_41), .b(gate494inter3), .O(gate494inter10));
  nor2  gate838(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate839(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate840(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate869(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate870(.a(gate496inter0), .b(s_46), .O(gate496inter1));
  and2  gate871(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate872(.a(s_46), .O(gate496inter3));
  inv1  gate873(.a(s_47), .O(gate496inter4));
  nand2 gate874(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate875(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate876(.a(G1254), .O(gate496inter7));
  inv1  gate877(.a(G1255), .O(gate496inter8));
  nand2 gate878(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate879(.a(s_47), .b(gate496inter3), .O(gate496inter10));
  nor2  gate880(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate881(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate882(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1513(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1514(.a(gate500inter0), .b(s_138), .O(gate500inter1));
  and2  gate1515(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1516(.a(s_138), .O(gate500inter3));
  inv1  gate1517(.a(s_139), .O(gate500inter4));
  nand2 gate1518(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1519(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1520(.a(G1262), .O(gate500inter7));
  inv1  gate1521(.a(G1263), .O(gate500inter8));
  nand2 gate1522(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1523(.a(s_139), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1524(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1525(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1526(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate813(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate814(.a(gate501inter0), .b(s_38), .O(gate501inter1));
  and2  gate815(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate816(.a(s_38), .O(gate501inter3));
  inv1  gate817(.a(s_39), .O(gate501inter4));
  nand2 gate818(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate819(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate820(.a(G1264), .O(gate501inter7));
  inv1  gate821(.a(G1265), .O(gate501inter8));
  nand2 gate822(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate823(.a(s_39), .b(gate501inter3), .O(gate501inter10));
  nor2  gate824(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate825(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate826(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1457(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1458(.a(gate505inter0), .b(s_130), .O(gate505inter1));
  and2  gate1459(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1460(.a(s_130), .O(gate505inter3));
  inv1  gate1461(.a(s_131), .O(gate505inter4));
  nand2 gate1462(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1463(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1464(.a(G1272), .O(gate505inter7));
  inv1  gate1465(.a(G1273), .O(gate505inter8));
  nand2 gate1466(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1467(.a(s_131), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1468(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1469(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1470(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1023(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1024(.a(gate510inter0), .b(s_68), .O(gate510inter1));
  and2  gate1025(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1026(.a(s_68), .O(gate510inter3));
  inv1  gate1027(.a(s_69), .O(gate510inter4));
  nand2 gate1028(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1029(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1030(.a(G1282), .O(gate510inter7));
  inv1  gate1031(.a(G1283), .O(gate510inter8));
  nand2 gate1032(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1033(.a(s_69), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1034(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1035(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1036(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate603(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate604(.a(gate514inter0), .b(s_8), .O(gate514inter1));
  and2  gate605(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate606(.a(s_8), .O(gate514inter3));
  inv1  gate607(.a(s_9), .O(gate514inter4));
  nand2 gate608(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate609(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate610(.a(G1290), .O(gate514inter7));
  inv1  gate611(.a(G1291), .O(gate514inter8));
  nand2 gate612(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate613(.a(s_9), .b(gate514inter3), .O(gate514inter10));
  nor2  gate614(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate615(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate616(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule