module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12;

  xor2  gate259(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate260(.a(gate1inter0), .b(s_8), .O(gate1inter1));
  and2  gate261(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate262(.a(s_8), .O(gate1inter3));
  inv1  gate263(.a(s_9), .O(gate1inter4));
  nand2 gate264(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate265(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate266(.a(N1), .O(gate1inter7));
  inv1  gate267(.a(N5), .O(gate1inter8));
  nand2 gate268(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate269(.a(s_9), .b(gate1inter3), .O(gate1inter10));
  nor2  gate270(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate271(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate272(.a(gate1inter12), .b(gate1inter1), .O(N250));

  xor2  gate609(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate610(.a(gate2inter0), .b(s_58), .O(gate2inter1));
  and2  gate611(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate612(.a(s_58), .O(gate2inter3));
  inv1  gate613(.a(s_59), .O(gate2inter4));
  nand2 gate614(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate615(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate616(.a(N9), .O(gate2inter7));
  inv1  gate617(.a(N13), .O(gate2inter8));
  nand2 gate618(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate619(.a(s_59), .b(gate2inter3), .O(gate2inter10));
  nor2  gate620(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate621(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate622(.a(gate2inter12), .b(gate2inter1), .O(N251));
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate301(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate302(.a(gate4inter0), .b(s_14), .O(gate4inter1));
  and2  gate303(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate304(.a(s_14), .O(gate4inter3));
  inv1  gate305(.a(s_15), .O(gate4inter4));
  nand2 gate306(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate307(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate308(.a(N25), .O(gate4inter7));
  inv1  gate309(.a(N29), .O(gate4inter8));
  nand2 gate310(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate311(.a(s_15), .b(gate4inter3), .O(gate4inter10));
  nor2  gate312(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate313(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate314(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate595(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate596(.a(gate6inter0), .b(s_56), .O(gate6inter1));
  and2  gate597(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate598(.a(s_56), .O(gate6inter3));
  inv1  gate599(.a(s_57), .O(gate6inter4));
  nand2 gate600(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate601(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate602(.a(N41), .O(gate6inter7));
  inv1  gate603(.a(N45), .O(gate6inter8));
  nand2 gate604(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate605(.a(s_57), .b(gate6inter3), .O(gate6inter10));
  nor2  gate606(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate607(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate608(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );

  xor2  gate763(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate764(.a(gate10inter0), .b(s_80), .O(gate10inter1));
  and2  gate765(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate766(.a(s_80), .O(gate10inter3));
  inv1  gate767(.a(s_81), .O(gate10inter4));
  nand2 gate768(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate769(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate770(.a(N73), .O(gate10inter7));
  inv1  gate771(.a(N77), .O(gate10inter8));
  nand2 gate772(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate773(.a(s_81), .b(gate10inter3), .O(gate10inter10));
  nor2  gate774(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate775(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate776(.a(gate10inter12), .b(gate10inter1), .O(N259));

  xor2  gate329(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate330(.a(gate11inter0), .b(s_18), .O(gate11inter1));
  and2  gate331(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate332(.a(s_18), .O(gate11inter3));
  inv1  gate333(.a(s_19), .O(gate11inter4));
  nand2 gate334(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate335(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate336(.a(N81), .O(gate11inter7));
  inv1  gate337(.a(N85), .O(gate11inter8));
  nand2 gate338(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate339(.a(s_19), .b(gate11inter3), .O(gate11inter10));
  nor2  gate340(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate341(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate342(.a(gate11inter12), .b(gate11inter1), .O(N260));
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );

  xor2  gate427(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate428(.a(gate15inter0), .b(s_32), .O(gate15inter1));
  and2  gate429(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate430(.a(s_32), .O(gate15inter3));
  inv1  gate431(.a(s_33), .O(gate15inter4));
  nand2 gate432(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate433(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate434(.a(N113), .O(gate15inter7));
  inv1  gate435(.a(N117), .O(gate15inter8));
  nand2 gate436(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate437(.a(s_33), .b(gate15inter3), .O(gate15inter10));
  nor2  gate438(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate439(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate440(.a(gate15inter12), .b(gate15inter1), .O(N264));
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );

  xor2  gate679(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate680(.a(gate26inter0), .b(s_68), .O(gate26inter1));
  and2  gate681(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate682(.a(s_68), .O(gate26inter3));
  inv1  gate683(.a(s_69), .O(gate26inter4));
  nand2 gate684(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate685(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate686(.a(N33), .O(gate26inter7));
  inv1  gate687(.a(N49), .O(gate26inter8));
  nand2 gate688(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate689(.a(s_69), .b(gate26inter3), .O(gate26inter10));
  nor2  gate690(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate691(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate692(.a(gate26inter12), .b(gate26inter1), .O(N275));

  xor2  gate693(.a(N21), .b(N5), .O(gate27inter0));
  nand2 gate694(.a(gate27inter0), .b(s_70), .O(gate27inter1));
  and2  gate695(.a(N21), .b(N5), .O(gate27inter2));
  inv1  gate696(.a(s_70), .O(gate27inter3));
  inv1  gate697(.a(s_71), .O(gate27inter4));
  nand2 gate698(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate699(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate700(.a(N5), .O(gate27inter7));
  inv1  gate701(.a(N21), .O(gate27inter8));
  nand2 gate702(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate703(.a(s_71), .b(gate27inter3), .O(gate27inter10));
  nor2  gate704(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate705(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate706(.a(gate27inter12), .b(gate27inter1), .O(N276));

  xor2  gate315(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate316(.a(gate28inter0), .b(s_16), .O(gate28inter1));
  and2  gate317(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate318(.a(s_16), .O(gate28inter3));
  inv1  gate319(.a(s_17), .O(gate28inter4));
  nand2 gate320(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate321(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate322(.a(N37), .O(gate28inter7));
  inv1  gate323(.a(N53), .O(gate28inter8));
  nand2 gate324(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate325(.a(s_17), .b(gate28inter3), .O(gate28inter10));
  nor2  gate326(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate327(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate328(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );

  xor2  gate749(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate750(.a(gate33inter0), .b(s_78), .O(gate33inter1));
  and2  gate751(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate752(.a(s_78), .O(gate33inter3));
  inv1  gate753(.a(s_79), .O(gate33inter4));
  nand2 gate754(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate755(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate756(.a(N65), .O(gate33inter7));
  inv1  gate757(.a(N81), .O(gate33inter8));
  nand2 gate758(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate759(.a(s_79), .b(gate33inter3), .O(gate33inter10));
  nor2  gate760(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate761(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate762(.a(gate33inter12), .b(gate33inter1), .O(N282));

  xor2  gate231(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate232(.a(gate34inter0), .b(s_4), .O(gate34inter1));
  and2  gate233(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate234(.a(s_4), .O(gate34inter3));
  inv1  gate235(.a(s_5), .O(gate34inter4));
  nand2 gate236(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate237(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate238(.a(N97), .O(gate34inter7));
  inv1  gate239(.a(N113), .O(gate34inter8));
  nand2 gate240(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate241(.a(s_5), .b(gate34inter3), .O(gate34inter10));
  nor2  gate242(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate243(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate244(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );

  xor2  gate287(.a(N93), .b(N77), .O(gate39inter0));
  nand2 gate288(.a(gate39inter0), .b(s_12), .O(gate39inter1));
  and2  gate289(.a(N93), .b(N77), .O(gate39inter2));
  inv1  gate290(.a(s_12), .O(gate39inter3));
  inv1  gate291(.a(s_13), .O(gate39inter4));
  nand2 gate292(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate293(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate294(.a(N77), .O(gate39inter7));
  inv1  gate295(.a(N93), .O(gate39inter8));
  nand2 gate296(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate297(.a(s_13), .b(gate39inter3), .O(gate39inter10));
  nor2  gate298(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate299(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate300(.a(gate39inter12), .b(gate39inter1), .O(N288));

  xor2  gate665(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate666(.a(gate40inter0), .b(s_66), .O(gate40inter1));
  and2  gate667(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate668(.a(s_66), .O(gate40inter3));
  inv1  gate669(.a(s_67), .O(gate40inter4));
  nand2 gate670(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate671(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate672(.a(N109), .O(gate40inter7));
  inv1  gate673(.a(N125), .O(gate40inter8));
  nand2 gate674(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate675(.a(s_67), .b(gate40inter3), .O(gate40inter10));
  nor2  gate676(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate677(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate678(.a(gate40inter12), .b(gate40inter1), .O(N289));
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate203(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate204(.a(gate47inter0), .b(s_0), .O(gate47inter1));
  and2  gate205(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate206(.a(s_0), .O(gate47inter3));
  inv1  gate207(.a(s_1), .O(gate47inter4));
  nand2 gate208(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate209(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate210(.a(N262), .O(gate47inter7));
  inv1  gate211(.a(N263), .O(gate47inter8));
  nand2 gate212(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate213(.a(s_1), .b(gate47inter3), .O(gate47inter10));
  nor2  gate214(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate215(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate216(.a(gate47inter12), .b(gate47inter1), .O(N308));
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );

  xor2  gate581(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate582(.a(gate54inter0), .b(s_54), .O(gate54inter1));
  and2  gate583(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate584(.a(s_54), .O(gate54inter3));
  inv1  gate585(.a(s_55), .O(gate54inter4));
  nand2 gate586(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate587(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate588(.a(N284), .O(gate54inter7));
  inv1  gate589(.a(N285), .O(gate54inter8));
  nand2 gate590(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate591(.a(s_55), .b(gate54inter3), .O(gate54inter10));
  nor2  gate592(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate593(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate594(.a(gate54inter12), .b(gate54inter1), .O(N319));

  xor2  gate385(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate386(.a(gate55inter0), .b(s_26), .O(gate55inter1));
  and2  gate387(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate388(.a(s_26), .O(gate55inter3));
  inv1  gate389(.a(s_27), .O(gate55inter4));
  nand2 gate390(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate391(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate392(.a(N286), .O(gate55inter7));
  inv1  gate393(.a(N287), .O(gate55inter8));
  nand2 gate394(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate395(.a(s_27), .b(gate55inter3), .O(gate55inter10));
  nor2  gate396(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate397(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate398(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate371(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate372(.a(gate59inter0), .b(s_24), .O(gate59inter1));
  and2  gate373(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate374(.a(s_24), .O(gate59inter3));
  inv1  gate375(.a(s_25), .O(gate59inter4));
  nand2 gate376(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate377(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate378(.a(N290), .O(gate59inter7));
  inv1  gate379(.a(N296), .O(gate59inter8));
  nand2 gate380(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate381(.a(s_25), .b(gate59inter3), .O(gate59inter10));
  nor2  gate382(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate383(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate384(.a(gate59inter12), .b(gate59inter1), .O(N340));

  xor2  gate469(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate470(.a(gate60inter0), .b(s_38), .O(gate60inter1));
  and2  gate471(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate472(.a(s_38), .O(gate60inter3));
  inv1  gate473(.a(s_39), .O(gate60inter4));
  nand2 gate474(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate475(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate476(.a(N293), .O(gate60inter7));
  inv1  gate477(.a(N299), .O(gate60inter8));
  nand2 gate478(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate479(.a(s_39), .b(gate60inter3), .O(gate60inter10));
  nor2  gate480(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate481(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate482(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate343(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate344(.a(gate62inter0), .b(s_20), .O(gate62inter1));
  and2  gate345(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate346(.a(s_20), .O(gate62inter3));
  inv1  gate347(.a(s_21), .O(gate62inter4));
  nand2 gate348(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate349(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate350(.a(N308), .O(gate62inter7));
  inv1  gate351(.a(N311), .O(gate62inter8));
  nand2 gate352(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate353(.a(s_21), .b(gate62inter3), .O(gate62inter10));
  nor2  gate354(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate355(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate356(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );

  xor2  gate413(.a(N345), .b(N269), .O(gate68inter0));
  nand2 gate414(.a(gate68inter0), .b(s_30), .O(gate68inter1));
  and2  gate415(.a(N345), .b(N269), .O(gate68inter2));
  inv1  gate416(.a(s_30), .O(gate68inter3));
  inv1  gate417(.a(s_31), .O(gate68inter4));
  nand2 gate418(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate419(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate420(.a(N269), .O(gate68inter7));
  inv1  gate421(.a(N345), .O(gate68inter8));
  nand2 gate422(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate423(.a(s_31), .b(gate68inter3), .O(gate68inter10));
  nor2  gate424(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate425(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate426(.a(gate68inter12), .b(gate68inter1), .O(N349));
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate217(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate218(.a(gate70inter0), .b(s_2), .O(gate70inter1));
  and2  gate219(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate220(.a(s_2), .O(gate70inter3));
  inv1  gate221(.a(s_3), .O(gate70inter4));
  nand2 gate222(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate223(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate224(.a(N271), .O(gate70inter7));
  inv1  gate225(.a(N339), .O(gate70inter8));
  nand2 gate226(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate227(.a(s_3), .b(gate70inter3), .O(gate70inter10));
  nor2  gate228(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate229(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate230(.a(gate70inter12), .b(gate70inter1), .O(N351));

  xor2  gate539(.a(N340), .b(N272), .O(gate71inter0));
  nand2 gate540(.a(gate71inter0), .b(s_48), .O(gate71inter1));
  and2  gate541(.a(N340), .b(N272), .O(gate71inter2));
  inv1  gate542(.a(s_48), .O(gate71inter3));
  inv1  gate543(.a(s_49), .O(gate71inter4));
  nand2 gate544(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate545(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate546(.a(N272), .O(gate71inter7));
  inv1  gate547(.a(N340), .O(gate71inter8));
  nand2 gate548(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate549(.a(s_49), .b(gate71inter3), .O(gate71inter10));
  nor2  gate550(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate551(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate552(.a(gate71inter12), .b(gate71inter1), .O(N352));
xor2 gate72( .a(N273), .b(N341), .O(N353) );

  xor2  gate497(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate498(.a(gate73inter0), .b(s_42), .O(gate73inter1));
  and2  gate499(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate500(.a(s_42), .O(gate73inter3));
  inv1  gate501(.a(s_43), .O(gate73inter4));
  nand2 gate502(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate503(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate504(.a(N314), .O(gate73inter7));
  inv1  gate505(.a(N346), .O(gate73inter8));
  nand2 gate506(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate507(.a(s_43), .b(gate73inter3), .O(gate73inter10));
  nor2  gate508(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate509(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate510(.a(gate73inter12), .b(gate73inter1), .O(N354));
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate735(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate736(.a(gate75inter0), .b(s_76), .O(gate75inter1));
  and2  gate737(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate738(.a(s_76), .O(gate75inter3));
  inv1  gate739(.a(s_77), .O(gate75inter4));
  nand2 gate740(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate741(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate742(.a(N316), .O(gate75inter7));
  inv1  gate743(.a(N348), .O(gate75inter8));
  nand2 gate744(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate745(.a(s_77), .b(gate75inter3), .O(gate75inter10));
  nor2  gate746(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate747(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate748(.a(gate75inter12), .b(gate75inter1), .O(N380));

  xor2  gate721(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate722(.a(gate76inter0), .b(s_74), .O(gate76inter1));
  and2  gate723(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate724(.a(s_74), .O(gate76inter3));
  inv1  gate725(.a(s_75), .O(gate76inter4));
  nand2 gate726(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate727(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate728(.a(N317), .O(gate76inter7));
  inv1  gate729(.a(N349), .O(gate76inter8));
  nand2 gate730(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate731(.a(s_75), .b(gate76inter3), .O(gate76inter10));
  nor2  gate732(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate733(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate734(.a(gate76inter12), .b(gate76inter1), .O(N393));

  xor2  gate553(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate554(.a(gate77inter0), .b(s_50), .O(gate77inter1));
  and2  gate555(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate556(.a(s_50), .O(gate77inter3));
  inv1  gate557(.a(s_51), .O(gate77inter4));
  nand2 gate558(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate559(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate560(.a(N318), .O(gate77inter7));
  inv1  gate561(.a(N350), .O(gate77inter8));
  nand2 gate562(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate563(.a(s_51), .b(gate77inter3), .O(gate77inter10));
  nor2  gate564(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate565(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate566(.a(gate77inter12), .b(gate77inter1), .O(N406));
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate399(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate400(.a(gate80inter0), .b(s_28), .O(gate80inter1));
  and2  gate401(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate402(.a(s_28), .O(gate80inter3));
  inv1  gate403(.a(s_29), .O(gate80inter4));
  nand2 gate404(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate405(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate406(.a(N321), .O(gate80inter7));
  inv1  gate407(.a(N353), .O(gate80inter8));
  nand2 gate408(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate409(.a(s_29), .b(gate80inter3), .O(gate80inter10));
  nor2  gate410(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate411(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate412(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );

  xor2  gate273(.a(N692), .b(N1), .O(gate171inter0));
  nand2 gate274(.a(gate171inter0), .b(s_10), .O(gate171inter1));
  and2  gate275(.a(N692), .b(N1), .O(gate171inter2));
  inv1  gate276(.a(s_10), .O(gate171inter3));
  inv1  gate277(.a(s_11), .O(gate171inter4));
  nand2 gate278(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate279(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate280(.a(N1), .O(gate171inter7));
  inv1  gate281(.a(N692), .O(gate171inter8));
  nand2 gate282(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate283(.a(s_11), .b(gate171inter3), .O(gate171inter10));
  nor2  gate284(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate285(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate286(.a(gate171inter12), .b(gate171inter1), .O(N724));

  xor2  gate455(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate456(.a(gate172inter0), .b(s_36), .O(gate172inter1));
  and2  gate457(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate458(.a(s_36), .O(gate172inter3));
  inv1  gate459(.a(s_37), .O(gate172inter4));
  nand2 gate460(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate461(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate462(.a(N5), .O(gate172inter7));
  inv1  gate463(.a(N693), .O(gate172inter8));
  nand2 gate464(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate465(.a(s_37), .b(gate172inter3), .O(gate172inter10));
  nor2  gate466(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate467(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate468(.a(gate172inter12), .b(gate172inter1), .O(N725));

  xor2  gate357(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate358(.a(gate173inter0), .b(s_22), .O(gate173inter1));
  and2  gate359(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate360(.a(s_22), .O(gate173inter3));
  inv1  gate361(.a(s_23), .O(gate173inter4));
  nand2 gate362(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate363(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate364(.a(N9), .O(gate173inter7));
  inv1  gate365(.a(N694), .O(gate173inter8));
  nand2 gate366(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate367(.a(s_23), .b(gate173inter3), .O(gate173inter10));
  nor2  gate368(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate369(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate370(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );

  xor2  gate651(.a(N696), .b(N17), .O(gate175inter0));
  nand2 gate652(.a(gate175inter0), .b(s_64), .O(gate175inter1));
  and2  gate653(.a(N696), .b(N17), .O(gate175inter2));
  inv1  gate654(.a(s_64), .O(gate175inter3));
  inv1  gate655(.a(s_65), .O(gate175inter4));
  nand2 gate656(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate657(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate658(.a(N17), .O(gate175inter7));
  inv1  gate659(.a(N696), .O(gate175inter8));
  nand2 gate660(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate661(.a(s_65), .b(gate175inter3), .O(gate175inter10));
  nor2  gate662(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate663(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate664(.a(gate175inter12), .b(gate175inter1), .O(N728));
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );

  xor2  gate567(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate568(.a(gate178inter0), .b(s_52), .O(gate178inter1));
  and2  gate569(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate570(.a(s_52), .O(gate178inter3));
  inv1  gate571(.a(s_53), .O(gate178inter4));
  nand2 gate572(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate573(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate574(.a(N29), .O(gate178inter7));
  inv1  gate575(.a(N699), .O(gate178inter8));
  nand2 gate576(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate577(.a(s_53), .b(gate178inter3), .O(gate178inter10));
  nor2  gate578(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate579(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate580(.a(gate178inter12), .b(gate178inter1), .O(N731));

  xor2  gate707(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate708(.a(gate179inter0), .b(s_72), .O(gate179inter1));
  and2  gate709(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate710(.a(s_72), .O(gate179inter3));
  inv1  gate711(.a(s_73), .O(gate179inter4));
  nand2 gate712(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate713(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate714(.a(N33), .O(gate179inter7));
  inv1  gate715(.a(N700), .O(gate179inter8));
  nand2 gate716(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate717(.a(s_73), .b(gate179inter3), .O(gate179inter10));
  nor2  gate718(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate719(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate720(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );

  xor2  gate623(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate624(.a(gate185inter0), .b(s_60), .O(gate185inter1));
  and2  gate625(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate626(.a(s_60), .O(gate185inter3));
  inv1  gate627(.a(s_61), .O(gate185inter4));
  nand2 gate628(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate629(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate630(.a(N57), .O(gate185inter7));
  inv1  gate631(.a(N706), .O(gate185inter8));
  nand2 gate632(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate633(.a(s_61), .b(gate185inter3), .O(gate185inter10));
  nor2  gate634(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate635(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate636(.a(gate185inter12), .b(gate185inter1), .O(N738));
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );

  xor2  gate441(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate442(.a(gate189inter0), .b(s_34), .O(gate189inter1));
  and2  gate443(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate444(.a(s_34), .O(gate189inter3));
  inv1  gate445(.a(s_35), .O(gate189inter4));
  nand2 gate446(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate447(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate448(.a(N73), .O(gate189inter7));
  inv1  gate449(.a(N710), .O(gate189inter8));
  nand2 gate450(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate451(.a(s_35), .b(gate189inter3), .O(gate189inter10));
  nor2  gate452(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate453(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate454(.a(gate189inter12), .b(gate189inter1), .O(N742));
xor2 gate190( .a(N77), .b(N711), .O(N743) );

  xor2  gate637(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate638(.a(gate191inter0), .b(s_62), .O(gate191inter1));
  and2  gate639(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate640(.a(s_62), .O(gate191inter3));
  inv1  gate641(.a(s_63), .O(gate191inter4));
  nand2 gate642(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate643(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate644(.a(N81), .O(gate191inter7));
  inv1  gate645(.a(N712), .O(gate191inter8));
  nand2 gate646(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate647(.a(s_63), .b(gate191inter3), .O(gate191inter10));
  nor2  gate648(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate649(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate650(.a(gate191inter12), .b(gate191inter1), .O(N744));
xor2 gate192( .a(N85), .b(N713), .O(N745) );

  xor2  gate525(.a(N714), .b(N89), .O(gate193inter0));
  nand2 gate526(.a(gate193inter0), .b(s_46), .O(gate193inter1));
  and2  gate527(.a(N714), .b(N89), .O(gate193inter2));
  inv1  gate528(.a(s_46), .O(gate193inter3));
  inv1  gate529(.a(s_47), .O(gate193inter4));
  nand2 gate530(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate531(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate532(.a(N89), .O(gate193inter7));
  inv1  gate533(.a(N714), .O(gate193inter8));
  nand2 gate534(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate535(.a(s_47), .b(gate193inter3), .O(gate193inter10));
  nor2  gate536(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate537(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate538(.a(gate193inter12), .b(gate193inter1), .O(N746));
xor2 gate194( .a(N93), .b(N715), .O(N747) );

  xor2  gate245(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate246(.a(gate195inter0), .b(s_6), .O(gate195inter1));
  and2  gate247(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate248(.a(s_6), .O(gate195inter3));
  inv1  gate249(.a(s_7), .O(gate195inter4));
  nand2 gate250(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate251(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate252(.a(N97), .O(gate195inter7));
  inv1  gate253(.a(N716), .O(gate195inter8));
  nand2 gate254(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate255(.a(s_7), .b(gate195inter3), .O(gate195inter10));
  nor2  gate256(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate257(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate258(.a(gate195inter12), .b(gate195inter1), .O(N748));
xor2 gate196( .a(N101), .b(N717), .O(N749) );

  xor2  gate483(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate484(.a(gate197inter0), .b(s_40), .O(gate197inter1));
  and2  gate485(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate486(.a(s_40), .O(gate197inter3));
  inv1  gate487(.a(s_41), .O(gate197inter4));
  nand2 gate488(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate489(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate490(.a(N105), .O(gate197inter7));
  inv1  gate491(.a(N718), .O(gate197inter8));
  nand2 gate492(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate493(.a(s_41), .b(gate197inter3), .O(gate197inter10));
  nor2  gate494(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate495(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate496(.a(gate197inter12), .b(gate197inter1), .O(N750));
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );

  xor2  gate511(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate512(.a(gate202inter0), .b(s_44), .O(gate202inter1));
  and2  gate513(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate514(.a(s_44), .O(gate202inter3));
  inv1  gate515(.a(s_45), .O(gate202inter4));
  nand2 gate516(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate517(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate518(.a(N125), .O(gate202inter7));
  inv1  gate519(.a(N723), .O(gate202inter8));
  nand2 gate520(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate521(.a(s_45), .b(gate202inter3), .O(gate202inter10));
  nor2  gate522(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate523(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate524(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule