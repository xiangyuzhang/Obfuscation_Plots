module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1303(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1304(.a(gate17inter0), .b(s_108), .O(gate17inter1));
  and2  gate1305(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1306(.a(s_108), .O(gate17inter3));
  inv1  gate1307(.a(s_109), .O(gate17inter4));
  nand2 gate1308(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1309(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1310(.a(G17), .O(gate17inter7));
  inv1  gate1311(.a(G18), .O(gate17inter8));
  nand2 gate1312(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1313(.a(s_109), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1314(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1315(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1316(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1233(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1234(.a(gate26inter0), .b(s_98), .O(gate26inter1));
  and2  gate1235(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1236(.a(s_98), .O(gate26inter3));
  inv1  gate1237(.a(s_99), .O(gate26inter4));
  nand2 gate1238(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1239(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1240(.a(G9), .O(gate26inter7));
  inv1  gate1241(.a(G13), .O(gate26inter8));
  nand2 gate1242(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1243(.a(s_99), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1244(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1245(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1246(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate729(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate730(.a(gate29inter0), .b(s_26), .O(gate29inter1));
  and2  gate731(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate732(.a(s_26), .O(gate29inter3));
  inv1  gate733(.a(s_27), .O(gate29inter4));
  nand2 gate734(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate735(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate736(.a(G3), .O(gate29inter7));
  inv1  gate737(.a(G7), .O(gate29inter8));
  nand2 gate738(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate739(.a(s_27), .b(gate29inter3), .O(gate29inter10));
  nor2  gate740(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate741(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate742(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate631(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate632(.a(gate31inter0), .b(s_12), .O(gate31inter1));
  and2  gate633(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate634(.a(s_12), .O(gate31inter3));
  inv1  gate635(.a(s_13), .O(gate31inter4));
  nand2 gate636(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate637(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate638(.a(G4), .O(gate31inter7));
  inv1  gate639(.a(G8), .O(gate31inter8));
  nand2 gate640(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate641(.a(s_13), .b(gate31inter3), .O(gate31inter10));
  nor2  gate642(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate643(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate644(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1023(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1024(.a(gate32inter0), .b(s_68), .O(gate32inter1));
  and2  gate1025(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1026(.a(s_68), .O(gate32inter3));
  inv1  gate1027(.a(s_69), .O(gate32inter4));
  nand2 gate1028(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1029(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1030(.a(G12), .O(gate32inter7));
  inv1  gate1031(.a(G16), .O(gate32inter8));
  nand2 gate1032(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1033(.a(s_69), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1034(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1035(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1036(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1317(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1318(.a(gate43inter0), .b(s_110), .O(gate43inter1));
  and2  gate1319(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1320(.a(s_110), .O(gate43inter3));
  inv1  gate1321(.a(s_111), .O(gate43inter4));
  nand2 gate1322(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1323(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1324(.a(G3), .O(gate43inter7));
  inv1  gate1325(.a(G269), .O(gate43inter8));
  nand2 gate1326(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1327(.a(s_111), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1328(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1329(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1330(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1611(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1612(.a(gate48inter0), .b(s_152), .O(gate48inter1));
  and2  gate1613(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1614(.a(s_152), .O(gate48inter3));
  inv1  gate1615(.a(s_153), .O(gate48inter4));
  nand2 gate1616(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1617(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1618(.a(G8), .O(gate48inter7));
  inv1  gate1619(.a(G275), .O(gate48inter8));
  nand2 gate1620(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1621(.a(s_153), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1622(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1623(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1624(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1975(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1976(.a(gate55inter0), .b(s_204), .O(gate55inter1));
  and2  gate1977(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1978(.a(s_204), .O(gate55inter3));
  inv1  gate1979(.a(s_205), .O(gate55inter4));
  nand2 gate1980(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1981(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1982(.a(G15), .O(gate55inter7));
  inv1  gate1983(.a(G287), .O(gate55inter8));
  nand2 gate1984(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1985(.a(s_205), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1986(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1987(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1988(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1065(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1066(.a(gate59inter0), .b(s_74), .O(gate59inter1));
  and2  gate1067(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1068(.a(s_74), .O(gate59inter3));
  inv1  gate1069(.a(s_75), .O(gate59inter4));
  nand2 gate1070(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1071(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1072(.a(G19), .O(gate59inter7));
  inv1  gate1073(.a(G293), .O(gate59inter8));
  nand2 gate1074(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1075(.a(s_75), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1076(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1077(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1078(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1709(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1710(.a(gate62inter0), .b(s_166), .O(gate62inter1));
  and2  gate1711(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1712(.a(s_166), .O(gate62inter3));
  inv1  gate1713(.a(s_167), .O(gate62inter4));
  nand2 gate1714(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1715(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1716(.a(G22), .O(gate62inter7));
  inv1  gate1717(.a(G296), .O(gate62inter8));
  nand2 gate1718(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1719(.a(s_167), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1720(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1721(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1722(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1681(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1682(.a(gate74inter0), .b(s_162), .O(gate74inter1));
  and2  gate1683(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1684(.a(s_162), .O(gate74inter3));
  inv1  gate1685(.a(s_163), .O(gate74inter4));
  nand2 gate1686(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1687(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1688(.a(G5), .O(gate74inter7));
  inv1  gate1689(.a(G314), .O(gate74inter8));
  nand2 gate1690(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1691(.a(s_163), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1692(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1693(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1694(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1835(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1836(.a(gate77inter0), .b(s_184), .O(gate77inter1));
  and2  gate1837(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1838(.a(s_184), .O(gate77inter3));
  inv1  gate1839(.a(s_185), .O(gate77inter4));
  nand2 gate1840(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1841(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1842(.a(G2), .O(gate77inter7));
  inv1  gate1843(.a(G320), .O(gate77inter8));
  nand2 gate1844(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1845(.a(s_185), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1846(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1847(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1848(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1639(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1640(.a(gate92inter0), .b(s_156), .O(gate92inter1));
  and2  gate1641(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1642(.a(s_156), .O(gate92inter3));
  inv1  gate1643(.a(s_157), .O(gate92inter4));
  nand2 gate1644(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1645(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1646(.a(G29), .O(gate92inter7));
  inv1  gate1647(.a(G341), .O(gate92inter8));
  nand2 gate1648(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1649(.a(s_157), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1650(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1651(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1652(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1219(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1220(.a(gate97inter0), .b(s_96), .O(gate97inter1));
  and2  gate1221(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1222(.a(s_96), .O(gate97inter3));
  inv1  gate1223(.a(s_97), .O(gate97inter4));
  nand2 gate1224(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1225(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1226(.a(G19), .O(gate97inter7));
  inv1  gate1227(.a(G350), .O(gate97inter8));
  nand2 gate1228(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1229(.a(s_97), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1230(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1231(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1232(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1541(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1542(.a(gate99inter0), .b(s_142), .O(gate99inter1));
  and2  gate1543(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1544(.a(s_142), .O(gate99inter3));
  inv1  gate1545(.a(s_143), .O(gate99inter4));
  nand2 gate1546(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1547(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1548(.a(G27), .O(gate99inter7));
  inv1  gate1549(.a(G353), .O(gate99inter8));
  nand2 gate1550(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1551(.a(s_143), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1552(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1553(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1554(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1667(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1668(.a(gate100inter0), .b(s_160), .O(gate100inter1));
  and2  gate1669(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1670(.a(s_160), .O(gate100inter3));
  inv1  gate1671(.a(s_161), .O(gate100inter4));
  nand2 gate1672(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1673(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1674(.a(G31), .O(gate100inter7));
  inv1  gate1675(.a(G353), .O(gate100inter8));
  nand2 gate1676(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1677(.a(s_161), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1678(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1679(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1680(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2017(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2018(.a(gate104inter0), .b(s_210), .O(gate104inter1));
  and2  gate2019(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2020(.a(s_210), .O(gate104inter3));
  inv1  gate2021(.a(s_211), .O(gate104inter4));
  nand2 gate2022(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2023(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2024(.a(G32), .O(gate104inter7));
  inv1  gate2025(.a(G359), .O(gate104inter8));
  nand2 gate2026(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2027(.a(s_211), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2028(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2029(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2030(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1163(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1164(.a(gate110inter0), .b(s_88), .O(gate110inter1));
  and2  gate1165(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1166(.a(s_88), .O(gate110inter3));
  inv1  gate1167(.a(s_89), .O(gate110inter4));
  nand2 gate1168(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1169(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1170(.a(G372), .O(gate110inter7));
  inv1  gate1171(.a(G373), .O(gate110inter8));
  nand2 gate1172(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1173(.a(s_89), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1174(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1175(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1176(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1387(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1388(.a(gate111inter0), .b(s_120), .O(gate111inter1));
  and2  gate1389(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1390(.a(s_120), .O(gate111inter3));
  inv1  gate1391(.a(s_121), .O(gate111inter4));
  nand2 gate1392(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1393(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1394(.a(G374), .O(gate111inter7));
  inv1  gate1395(.a(G375), .O(gate111inter8));
  nand2 gate1396(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1397(.a(s_121), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1398(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1399(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1400(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1527(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1528(.a(gate114inter0), .b(s_140), .O(gate114inter1));
  and2  gate1529(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1530(.a(s_140), .O(gate114inter3));
  inv1  gate1531(.a(s_141), .O(gate114inter4));
  nand2 gate1532(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1533(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1534(.a(G380), .O(gate114inter7));
  inv1  gate1535(.a(G381), .O(gate114inter8));
  nand2 gate1536(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1537(.a(s_141), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1538(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1539(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1540(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate743(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate744(.a(gate117inter0), .b(s_28), .O(gate117inter1));
  and2  gate745(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate746(.a(s_28), .O(gate117inter3));
  inv1  gate747(.a(s_29), .O(gate117inter4));
  nand2 gate748(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate749(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate750(.a(G386), .O(gate117inter7));
  inv1  gate751(.a(G387), .O(gate117inter8));
  nand2 gate752(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate753(.a(s_29), .b(gate117inter3), .O(gate117inter10));
  nor2  gate754(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate755(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate756(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1289(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1290(.a(gate121inter0), .b(s_106), .O(gate121inter1));
  and2  gate1291(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1292(.a(s_106), .O(gate121inter3));
  inv1  gate1293(.a(s_107), .O(gate121inter4));
  nand2 gate1294(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1295(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1296(.a(G394), .O(gate121inter7));
  inv1  gate1297(.a(G395), .O(gate121inter8));
  nand2 gate1298(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1299(.a(s_107), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1300(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1301(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1302(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2003(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2004(.a(gate125inter0), .b(s_208), .O(gate125inter1));
  and2  gate2005(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2006(.a(s_208), .O(gate125inter3));
  inv1  gate2007(.a(s_209), .O(gate125inter4));
  nand2 gate2008(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2009(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2010(.a(G402), .O(gate125inter7));
  inv1  gate2011(.a(G403), .O(gate125inter8));
  nand2 gate2012(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2013(.a(s_209), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2014(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2015(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2016(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1079(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1080(.a(gate132inter0), .b(s_76), .O(gate132inter1));
  and2  gate1081(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1082(.a(s_76), .O(gate132inter3));
  inv1  gate1083(.a(s_77), .O(gate132inter4));
  nand2 gate1084(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1085(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1086(.a(G416), .O(gate132inter7));
  inv1  gate1087(.a(G417), .O(gate132inter8));
  nand2 gate1088(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1089(.a(s_77), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1090(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1091(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1092(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1443(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1444(.a(gate133inter0), .b(s_128), .O(gate133inter1));
  and2  gate1445(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1446(.a(s_128), .O(gate133inter3));
  inv1  gate1447(.a(s_129), .O(gate133inter4));
  nand2 gate1448(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1449(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1450(.a(G418), .O(gate133inter7));
  inv1  gate1451(.a(G419), .O(gate133inter8));
  nand2 gate1452(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1453(.a(s_129), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1454(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1455(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1456(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1121(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1122(.a(gate136inter0), .b(s_82), .O(gate136inter1));
  and2  gate1123(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1124(.a(s_82), .O(gate136inter3));
  inv1  gate1125(.a(s_83), .O(gate136inter4));
  nand2 gate1126(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1127(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1128(.a(G424), .O(gate136inter7));
  inv1  gate1129(.a(G425), .O(gate136inter8));
  nand2 gate1130(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1131(.a(s_83), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1132(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1133(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1134(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1485(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1486(.a(gate139inter0), .b(s_134), .O(gate139inter1));
  and2  gate1487(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1488(.a(s_134), .O(gate139inter3));
  inv1  gate1489(.a(s_135), .O(gate139inter4));
  nand2 gate1490(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1491(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1492(.a(G438), .O(gate139inter7));
  inv1  gate1493(.a(G441), .O(gate139inter8));
  nand2 gate1494(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1495(.a(s_135), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1496(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1497(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1498(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1247(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1248(.a(gate140inter0), .b(s_100), .O(gate140inter1));
  and2  gate1249(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1250(.a(s_100), .O(gate140inter3));
  inv1  gate1251(.a(s_101), .O(gate140inter4));
  nand2 gate1252(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1253(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1254(.a(G444), .O(gate140inter7));
  inv1  gate1255(.a(G447), .O(gate140inter8));
  nand2 gate1256(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1257(.a(s_101), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1258(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1259(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1260(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1751(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1752(.a(gate143inter0), .b(s_172), .O(gate143inter1));
  and2  gate1753(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1754(.a(s_172), .O(gate143inter3));
  inv1  gate1755(.a(s_173), .O(gate143inter4));
  nand2 gate1756(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1757(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1758(.a(G462), .O(gate143inter7));
  inv1  gate1759(.a(G465), .O(gate143inter8));
  nand2 gate1760(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1761(.a(s_173), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1762(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1763(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1764(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate673(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate674(.a(gate144inter0), .b(s_18), .O(gate144inter1));
  and2  gate675(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate676(.a(s_18), .O(gate144inter3));
  inv1  gate677(.a(s_19), .O(gate144inter4));
  nand2 gate678(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate679(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate680(.a(G468), .O(gate144inter7));
  inv1  gate681(.a(G471), .O(gate144inter8));
  nand2 gate682(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate683(.a(s_19), .b(gate144inter3), .O(gate144inter10));
  nor2  gate684(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate685(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate686(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate701(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate702(.a(gate145inter0), .b(s_22), .O(gate145inter1));
  and2  gate703(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate704(.a(s_22), .O(gate145inter3));
  inv1  gate705(.a(s_23), .O(gate145inter4));
  nand2 gate706(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate707(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate708(.a(G474), .O(gate145inter7));
  inv1  gate709(.a(G477), .O(gate145inter8));
  nand2 gate710(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate711(.a(s_23), .b(gate145inter3), .O(gate145inter10));
  nor2  gate712(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate713(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate714(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1737(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1738(.a(gate148inter0), .b(s_170), .O(gate148inter1));
  and2  gate1739(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1740(.a(s_170), .O(gate148inter3));
  inv1  gate1741(.a(s_171), .O(gate148inter4));
  nand2 gate1742(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1743(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1744(.a(G492), .O(gate148inter7));
  inv1  gate1745(.a(G495), .O(gate148inter8));
  nand2 gate1746(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1747(.a(s_171), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1748(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1749(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1750(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1919(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1920(.a(gate151inter0), .b(s_196), .O(gate151inter1));
  and2  gate1921(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1922(.a(s_196), .O(gate151inter3));
  inv1  gate1923(.a(s_197), .O(gate151inter4));
  nand2 gate1924(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1925(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1926(.a(G510), .O(gate151inter7));
  inv1  gate1927(.a(G513), .O(gate151inter8));
  nand2 gate1928(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1929(.a(s_197), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1930(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1931(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1932(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1779(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1780(.a(gate155inter0), .b(s_176), .O(gate155inter1));
  and2  gate1781(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1782(.a(s_176), .O(gate155inter3));
  inv1  gate1783(.a(s_177), .O(gate155inter4));
  nand2 gate1784(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1785(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1786(.a(G432), .O(gate155inter7));
  inv1  gate1787(.a(G525), .O(gate155inter8));
  nand2 gate1788(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1789(.a(s_177), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1790(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1791(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1792(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate799(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate800(.a(gate157inter0), .b(s_36), .O(gate157inter1));
  and2  gate801(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate802(.a(s_36), .O(gate157inter3));
  inv1  gate803(.a(s_37), .O(gate157inter4));
  nand2 gate804(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate805(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate806(.a(G438), .O(gate157inter7));
  inv1  gate807(.a(G528), .O(gate157inter8));
  nand2 gate808(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate809(.a(s_37), .b(gate157inter3), .O(gate157inter10));
  nor2  gate810(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate811(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate812(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1093(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1094(.a(gate174inter0), .b(s_78), .O(gate174inter1));
  and2  gate1095(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1096(.a(s_78), .O(gate174inter3));
  inv1  gate1097(.a(s_79), .O(gate174inter4));
  nand2 gate1098(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1099(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1100(.a(G489), .O(gate174inter7));
  inv1  gate1101(.a(G552), .O(gate174inter8));
  nand2 gate1102(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1103(.a(s_79), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1104(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1105(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1106(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1401(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1402(.a(gate190inter0), .b(s_122), .O(gate190inter1));
  and2  gate1403(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1404(.a(s_122), .O(gate190inter3));
  inv1  gate1405(.a(s_123), .O(gate190inter4));
  nand2 gate1406(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1407(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1408(.a(G580), .O(gate190inter7));
  inv1  gate1409(.a(G581), .O(gate190inter8));
  nand2 gate1410(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1411(.a(s_123), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1412(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1413(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1414(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate995(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate996(.a(gate192inter0), .b(s_64), .O(gate192inter1));
  and2  gate997(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate998(.a(s_64), .O(gate192inter3));
  inv1  gate999(.a(s_65), .O(gate192inter4));
  nand2 gate1000(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1001(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1002(.a(G584), .O(gate192inter7));
  inv1  gate1003(.a(G585), .O(gate192inter8));
  nand2 gate1004(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1005(.a(s_65), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1006(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1007(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1008(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1471(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1472(.a(gate194inter0), .b(s_132), .O(gate194inter1));
  and2  gate1473(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1474(.a(s_132), .O(gate194inter3));
  inv1  gate1475(.a(s_133), .O(gate194inter4));
  nand2 gate1476(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1477(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1478(.a(G588), .O(gate194inter7));
  inv1  gate1479(.a(G589), .O(gate194inter8));
  nand2 gate1480(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1481(.a(s_133), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1482(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1483(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1484(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1191(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1192(.a(gate203inter0), .b(s_92), .O(gate203inter1));
  and2  gate1193(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1194(.a(s_92), .O(gate203inter3));
  inv1  gate1195(.a(s_93), .O(gate203inter4));
  nand2 gate1196(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1197(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1198(.a(G602), .O(gate203inter7));
  inv1  gate1199(.a(G612), .O(gate203inter8));
  nand2 gate1200(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1201(.a(s_93), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1202(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1203(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1204(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1849(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1850(.a(gate204inter0), .b(s_186), .O(gate204inter1));
  and2  gate1851(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1852(.a(s_186), .O(gate204inter3));
  inv1  gate1853(.a(s_187), .O(gate204inter4));
  nand2 gate1854(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1855(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1856(.a(G607), .O(gate204inter7));
  inv1  gate1857(.a(G617), .O(gate204inter8));
  nand2 gate1858(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1859(.a(s_187), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1860(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1861(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1862(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1583(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1584(.a(gate212inter0), .b(s_148), .O(gate212inter1));
  and2  gate1585(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1586(.a(s_148), .O(gate212inter3));
  inv1  gate1587(.a(s_149), .O(gate212inter4));
  nand2 gate1588(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1589(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1590(.a(G617), .O(gate212inter7));
  inv1  gate1591(.a(G669), .O(gate212inter8));
  nand2 gate1592(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1593(.a(s_149), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1594(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1595(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1596(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate603(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate604(.a(gate216inter0), .b(s_8), .O(gate216inter1));
  and2  gate605(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate606(.a(s_8), .O(gate216inter3));
  inv1  gate607(.a(s_9), .O(gate216inter4));
  nand2 gate608(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate609(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate610(.a(G617), .O(gate216inter7));
  inv1  gate611(.a(G675), .O(gate216inter8));
  nand2 gate612(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate613(.a(s_9), .b(gate216inter3), .O(gate216inter10));
  nor2  gate614(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate615(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate616(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate785(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate786(.a(gate219inter0), .b(s_34), .O(gate219inter1));
  and2  gate787(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate788(.a(s_34), .O(gate219inter3));
  inv1  gate789(.a(s_35), .O(gate219inter4));
  nand2 gate790(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate791(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate792(.a(G632), .O(gate219inter7));
  inv1  gate793(.a(G681), .O(gate219inter8));
  nand2 gate794(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate795(.a(s_35), .b(gate219inter3), .O(gate219inter10));
  nor2  gate796(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate797(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate798(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate617(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate618(.a(gate220inter0), .b(s_10), .O(gate220inter1));
  and2  gate619(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate620(.a(s_10), .O(gate220inter3));
  inv1  gate621(.a(s_11), .O(gate220inter4));
  nand2 gate622(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate623(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate624(.a(G637), .O(gate220inter7));
  inv1  gate625(.a(G681), .O(gate220inter8));
  nand2 gate626(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate627(.a(s_11), .b(gate220inter3), .O(gate220inter10));
  nor2  gate628(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate629(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate630(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1807(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1808(.a(gate222inter0), .b(s_180), .O(gate222inter1));
  and2  gate1809(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1810(.a(s_180), .O(gate222inter3));
  inv1  gate1811(.a(s_181), .O(gate222inter4));
  nand2 gate1812(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1813(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1814(.a(G632), .O(gate222inter7));
  inv1  gate1815(.a(G684), .O(gate222inter8));
  nand2 gate1816(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1817(.a(s_181), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1818(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1819(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1820(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate813(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate814(.a(gate223inter0), .b(s_38), .O(gate223inter1));
  and2  gate815(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate816(.a(s_38), .O(gate223inter3));
  inv1  gate817(.a(s_39), .O(gate223inter4));
  nand2 gate818(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate819(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate820(.a(G627), .O(gate223inter7));
  inv1  gate821(.a(G687), .O(gate223inter8));
  nand2 gate822(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate823(.a(s_39), .b(gate223inter3), .O(gate223inter10));
  nor2  gate824(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate825(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate826(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1625(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1626(.a(gate227inter0), .b(s_154), .O(gate227inter1));
  and2  gate1627(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1628(.a(s_154), .O(gate227inter3));
  inv1  gate1629(.a(s_155), .O(gate227inter4));
  nand2 gate1630(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1631(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1632(.a(G694), .O(gate227inter7));
  inv1  gate1633(.a(G695), .O(gate227inter8));
  nand2 gate1634(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1635(.a(s_155), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1636(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1637(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1638(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate715(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate716(.a(gate229inter0), .b(s_24), .O(gate229inter1));
  and2  gate717(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate718(.a(s_24), .O(gate229inter3));
  inv1  gate719(.a(s_25), .O(gate229inter4));
  nand2 gate720(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate721(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate722(.a(G698), .O(gate229inter7));
  inv1  gate723(.a(G699), .O(gate229inter8));
  nand2 gate724(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate725(.a(s_25), .b(gate229inter3), .O(gate229inter10));
  nor2  gate726(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate727(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate728(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1331(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1332(.a(gate231inter0), .b(s_112), .O(gate231inter1));
  and2  gate1333(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1334(.a(s_112), .O(gate231inter3));
  inv1  gate1335(.a(s_113), .O(gate231inter4));
  nand2 gate1336(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1337(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1338(.a(G702), .O(gate231inter7));
  inv1  gate1339(.a(G703), .O(gate231inter8));
  nand2 gate1340(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1341(.a(s_113), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1342(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1343(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1344(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1947(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1948(.a(gate233inter0), .b(s_200), .O(gate233inter1));
  and2  gate1949(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1950(.a(s_200), .O(gate233inter3));
  inv1  gate1951(.a(s_201), .O(gate233inter4));
  nand2 gate1952(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1953(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1954(.a(G242), .O(gate233inter7));
  inv1  gate1955(.a(G718), .O(gate233inter8));
  nand2 gate1956(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1957(.a(s_201), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1958(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1959(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1960(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1555(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1556(.a(gate242inter0), .b(s_144), .O(gate242inter1));
  and2  gate1557(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1558(.a(s_144), .O(gate242inter3));
  inv1  gate1559(.a(s_145), .O(gate242inter4));
  nand2 gate1560(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1561(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1562(.a(G718), .O(gate242inter7));
  inv1  gate1563(.a(G730), .O(gate242inter8));
  nand2 gate1564(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1565(.a(s_145), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1566(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1567(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1568(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1149(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1150(.a(gate244inter0), .b(s_86), .O(gate244inter1));
  and2  gate1151(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1152(.a(s_86), .O(gate244inter3));
  inv1  gate1153(.a(s_87), .O(gate244inter4));
  nand2 gate1154(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1155(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1156(.a(G721), .O(gate244inter7));
  inv1  gate1157(.a(G733), .O(gate244inter8));
  nand2 gate1158(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1159(.a(s_87), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1160(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1161(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1162(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1891(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1892(.a(gate245inter0), .b(s_192), .O(gate245inter1));
  and2  gate1893(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1894(.a(s_192), .O(gate245inter3));
  inv1  gate1895(.a(s_193), .O(gate245inter4));
  nand2 gate1896(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1897(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1898(.a(G248), .O(gate245inter7));
  inv1  gate1899(.a(G736), .O(gate245inter8));
  nand2 gate1900(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1901(.a(s_193), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1902(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1903(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1904(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate757(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate758(.a(gate259inter0), .b(s_30), .O(gate259inter1));
  and2  gate759(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate760(.a(s_30), .O(gate259inter3));
  inv1  gate761(.a(s_31), .O(gate259inter4));
  nand2 gate762(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate763(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate764(.a(G758), .O(gate259inter7));
  inv1  gate765(.a(G759), .O(gate259inter8));
  nand2 gate766(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate767(.a(s_31), .b(gate259inter3), .O(gate259inter10));
  nor2  gate768(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate769(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate770(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate925(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate926(.a(gate261inter0), .b(s_54), .O(gate261inter1));
  and2  gate927(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate928(.a(s_54), .O(gate261inter3));
  inv1  gate929(.a(s_55), .O(gate261inter4));
  nand2 gate930(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate931(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate932(.a(G762), .O(gate261inter7));
  inv1  gate933(.a(G763), .O(gate261inter8));
  nand2 gate934(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate935(.a(s_55), .b(gate261inter3), .O(gate261inter10));
  nor2  gate936(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate937(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate938(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate953(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate954(.a(gate262inter0), .b(s_58), .O(gate262inter1));
  and2  gate955(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate956(.a(s_58), .O(gate262inter3));
  inv1  gate957(.a(s_59), .O(gate262inter4));
  nand2 gate958(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate959(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate960(.a(G764), .O(gate262inter7));
  inv1  gate961(.a(G765), .O(gate262inter8));
  nand2 gate962(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate963(.a(s_59), .b(gate262inter3), .O(gate262inter10));
  nor2  gate964(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate965(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate966(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1863(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1864(.a(gate265inter0), .b(s_188), .O(gate265inter1));
  and2  gate1865(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1866(.a(s_188), .O(gate265inter3));
  inv1  gate1867(.a(s_189), .O(gate265inter4));
  nand2 gate1868(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1869(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1870(.a(G642), .O(gate265inter7));
  inv1  gate1871(.a(G770), .O(gate265inter8));
  nand2 gate1872(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1873(.a(s_189), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1874(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1875(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1876(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate897(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate898(.a(gate267inter0), .b(s_50), .O(gate267inter1));
  and2  gate899(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate900(.a(s_50), .O(gate267inter3));
  inv1  gate901(.a(s_51), .O(gate267inter4));
  nand2 gate902(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate903(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate904(.a(G648), .O(gate267inter7));
  inv1  gate905(.a(G776), .O(gate267inter8));
  nand2 gate906(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate907(.a(s_51), .b(gate267inter3), .O(gate267inter10));
  nor2  gate908(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate909(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate910(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1933(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1934(.a(gate271inter0), .b(s_198), .O(gate271inter1));
  and2  gate1935(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1936(.a(s_198), .O(gate271inter3));
  inv1  gate1937(.a(s_199), .O(gate271inter4));
  nand2 gate1938(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1939(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1940(.a(G660), .O(gate271inter7));
  inv1  gate1941(.a(G788), .O(gate271inter8));
  nand2 gate1942(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1943(.a(s_199), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1944(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1945(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1946(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate575(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate576(.a(gate273inter0), .b(s_4), .O(gate273inter1));
  and2  gate577(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate578(.a(s_4), .O(gate273inter3));
  inv1  gate579(.a(s_5), .O(gate273inter4));
  nand2 gate580(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate581(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate582(.a(G642), .O(gate273inter7));
  inv1  gate583(.a(G794), .O(gate273inter8));
  nand2 gate584(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate585(.a(s_5), .b(gate273inter3), .O(gate273inter10));
  nor2  gate586(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate587(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate588(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate561(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate562(.a(gate275inter0), .b(s_2), .O(gate275inter1));
  and2  gate563(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate564(.a(s_2), .O(gate275inter3));
  inv1  gate565(.a(s_3), .O(gate275inter4));
  nand2 gate566(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate567(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate568(.a(G645), .O(gate275inter7));
  inv1  gate569(.a(G797), .O(gate275inter8));
  nand2 gate570(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate571(.a(s_3), .b(gate275inter3), .O(gate275inter10));
  nor2  gate572(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate573(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate574(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1275(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1276(.a(gate280inter0), .b(s_104), .O(gate280inter1));
  and2  gate1277(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1278(.a(s_104), .O(gate280inter3));
  inv1  gate1279(.a(s_105), .O(gate280inter4));
  nand2 gate1280(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1281(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1282(.a(G779), .O(gate280inter7));
  inv1  gate1283(.a(G803), .O(gate280inter8));
  nand2 gate1284(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1285(.a(s_105), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1286(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1287(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1288(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate645(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate646(.a(gate281inter0), .b(s_14), .O(gate281inter1));
  and2  gate647(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate648(.a(s_14), .O(gate281inter3));
  inv1  gate649(.a(s_15), .O(gate281inter4));
  nand2 gate650(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate651(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate652(.a(G654), .O(gate281inter7));
  inv1  gate653(.a(G806), .O(gate281inter8));
  nand2 gate654(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate655(.a(s_15), .b(gate281inter3), .O(gate281inter10));
  nor2  gate656(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate657(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate658(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1037(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1038(.a(gate282inter0), .b(s_70), .O(gate282inter1));
  and2  gate1039(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1040(.a(s_70), .O(gate282inter3));
  inv1  gate1041(.a(s_71), .O(gate282inter4));
  nand2 gate1042(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1043(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1044(.a(G782), .O(gate282inter7));
  inv1  gate1045(.a(G806), .O(gate282inter8));
  nand2 gate1046(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1047(.a(s_71), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1048(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1049(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1050(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1821(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1822(.a(gate283inter0), .b(s_182), .O(gate283inter1));
  and2  gate1823(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1824(.a(s_182), .O(gate283inter3));
  inv1  gate1825(.a(s_183), .O(gate283inter4));
  nand2 gate1826(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1827(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1828(.a(G657), .O(gate283inter7));
  inv1  gate1829(.a(G809), .O(gate283inter8));
  nand2 gate1830(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1831(.a(s_183), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1832(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1833(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1834(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate659(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate660(.a(gate284inter0), .b(s_16), .O(gate284inter1));
  and2  gate661(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate662(.a(s_16), .O(gate284inter3));
  inv1  gate663(.a(s_17), .O(gate284inter4));
  nand2 gate664(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate665(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate666(.a(G785), .O(gate284inter7));
  inv1  gate667(.a(G809), .O(gate284inter8));
  nand2 gate668(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate669(.a(s_17), .b(gate284inter3), .O(gate284inter10));
  nor2  gate670(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate671(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate672(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1765(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1766(.a(gate287inter0), .b(s_174), .O(gate287inter1));
  and2  gate1767(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1768(.a(s_174), .O(gate287inter3));
  inv1  gate1769(.a(s_175), .O(gate287inter4));
  nand2 gate1770(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1771(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1772(.a(G663), .O(gate287inter7));
  inv1  gate1773(.a(G815), .O(gate287inter8));
  nand2 gate1774(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1775(.a(s_175), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1776(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1777(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1778(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate869(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate870(.a(gate291inter0), .b(s_46), .O(gate291inter1));
  and2  gate871(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate872(.a(s_46), .O(gate291inter3));
  inv1  gate873(.a(s_47), .O(gate291inter4));
  nand2 gate874(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate875(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate876(.a(G822), .O(gate291inter7));
  inv1  gate877(.a(G823), .O(gate291inter8));
  nand2 gate878(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate879(.a(s_47), .b(gate291inter3), .O(gate291inter10));
  nor2  gate880(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate881(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate882(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate827(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate828(.a(gate292inter0), .b(s_40), .O(gate292inter1));
  and2  gate829(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate830(.a(s_40), .O(gate292inter3));
  inv1  gate831(.a(s_41), .O(gate292inter4));
  nand2 gate832(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate833(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate834(.a(G824), .O(gate292inter7));
  inv1  gate835(.a(G825), .O(gate292inter8));
  nand2 gate836(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate837(.a(s_41), .b(gate292inter3), .O(gate292inter10));
  nor2  gate838(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate839(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate840(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate771(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate772(.a(gate293inter0), .b(s_32), .O(gate293inter1));
  and2  gate773(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate774(.a(s_32), .O(gate293inter3));
  inv1  gate775(.a(s_33), .O(gate293inter4));
  nand2 gate776(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate777(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate778(.a(G828), .O(gate293inter7));
  inv1  gate779(.a(G829), .O(gate293inter8));
  nand2 gate780(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate781(.a(s_33), .b(gate293inter3), .O(gate293inter10));
  nor2  gate782(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate783(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate784(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1989(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1990(.a(gate390inter0), .b(s_206), .O(gate390inter1));
  and2  gate1991(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1992(.a(s_206), .O(gate390inter3));
  inv1  gate1993(.a(s_207), .O(gate390inter4));
  nand2 gate1994(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1995(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1996(.a(G4), .O(gate390inter7));
  inv1  gate1997(.a(G1045), .O(gate390inter8));
  nand2 gate1998(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1999(.a(s_207), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2000(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2001(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2002(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1345(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1346(.a(gate392inter0), .b(s_114), .O(gate392inter1));
  and2  gate1347(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1348(.a(s_114), .O(gate392inter3));
  inv1  gate1349(.a(s_115), .O(gate392inter4));
  nand2 gate1350(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1351(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1352(.a(G6), .O(gate392inter7));
  inv1  gate1353(.a(G1051), .O(gate392inter8));
  nand2 gate1354(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1355(.a(s_115), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1356(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1357(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1358(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate911(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate912(.a(gate395inter0), .b(s_52), .O(gate395inter1));
  and2  gate913(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate914(.a(s_52), .O(gate395inter3));
  inv1  gate915(.a(s_53), .O(gate395inter4));
  nand2 gate916(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate917(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate918(.a(G9), .O(gate395inter7));
  inv1  gate919(.a(G1060), .O(gate395inter8));
  nand2 gate920(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate921(.a(s_53), .b(gate395inter3), .O(gate395inter10));
  nor2  gate922(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate923(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate924(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1499(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1500(.a(gate398inter0), .b(s_136), .O(gate398inter1));
  and2  gate1501(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1502(.a(s_136), .O(gate398inter3));
  inv1  gate1503(.a(s_137), .O(gate398inter4));
  nand2 gate1504(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1505(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1506(.a(G12), .O(gate398inter7));
  inv1  gate1507(.a(G1069), .O(gate398inter8));
  nand2 gate1508(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1509(.a(s_137), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1510(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1511(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1512(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1205(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1206(.a(gate402inter0), .b(s_94), .O(gate402inter1));
  and2  gate1207(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1208(.a(s_94), .O(gate402inter3));
  inv1  gate1209(.a(s_95), .O(gate402inter4));
  nand2 gate1210(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1211(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1212(.a(G16), .O(gate402inter7));
  inv1  gate1213(.a(G1081), .O(gate402inter8));
  nand2 gate1214(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1215(.a(s_95), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1216(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1217(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1218(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1429(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1430(.a(gate403inter0), .b(s_126), .O(gate403inter1));
  and2  gate1431(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1432(.a(s_126), .O(gate403inter3));
  inv1  gate1433(.a(s_127), .O(gate403inter4));
  nand2 gate1434(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1435(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1436(.a(G17), .O(gate403inter7));
  inv1  gate1437(.a(G1084), .O(gate403inter8));
  nand2 gate1438(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1439(.a(s_127), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1440(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1441(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1442(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1051(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1052(.a(gate404inter0), .b(s_72), .O(gate404inter1));
  and2  gate1053(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1054(.a(s_72), .O(gate404inter3));
  inv1  gate1055(.a(s_73), .O(gate404inter4));
  nand2 gate1056(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1057(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1058(.a(G18), .O(gate404inter7));
  inv1  gate1059(.a(G1087), .O(gate404inter8));
  nand2 gate1060(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1061(.a(s_73), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1062(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1063(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1064(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1905(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1906(.a(gate408inter0), .b(s_194), .O(gate408inter1));
  and2  gate1907(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1908(.a(s_194), .O(gate408inter3));
  inv1  gate1909(.a(s_195), .O(gate408inter4));
  nand2 gate1910(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1911(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1912(.a(G22), .O(gate408inter7));
  inv1  gate1913(.a(G1099), .O(gate408inter8));
  nand2 gate1914(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1915(.a(s_195), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1916(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1917(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1918(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1359(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1360(.a(gate411inter0), .b(s_116), .O(gate411inter1));
  and2  gate1361(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1362(.a(s_116), .O(gate411inter3));
  inv1  gate1363(.a(s_117), .O(gate411inter4));
  nand2 gate1364(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1365(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1366(.a(G25), .O(gate411inter7));
  inv1  gate1367(.a(G1108), .O(gate411inter8));
  nand2 gate1368(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1369(.a(s_117), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1370(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1371(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1372(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate939(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate940(.a(gate414inter0), .b(s_56), .O(gate414inter1));
  and2  gate941(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate942(.a(s_56), .O(gate414inter3));
  inv1  gate943(.a(s_57), .O(gate414inter4));
  nand2 gate944(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate945(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate946(.a(G28), .O(gate414inter7));
  inv1  gate947(.a(G1117), .O(gate414inter8));
  nand2 gate948(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate949(.a(s_57), .b(gate414inter3), .O(gate414inter10));
  nor2  gate950(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate951(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate952(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1723(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1724(.a(gate415inter0), .b(s_168), .O(gate415inter1));
  and2  gate1725(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1726(.a(s_168), .O(gate415inter3));
  inv1  gate1727(.a(s_169), .O(gate415inter4));
  nand2 gate1728(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1729(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1730(.a(G29), .O(gate415inter7));
  inv1  gate1731(.a(G1120), .O(gate415inter8));
  nand2 gate1732(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1733(.a(s_169), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1734(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1735(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1736(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1961(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1962(.a(gate420inter0), .b(s_202), .O(gate420inter1));
  and2  gate1963(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1964(.a(s_202), .O(gate420inter3));
  inv1  gate1965(.a(s_203), .O(gate420inter4));
  nand2 gate1966(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1967(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1968(.a(G1036), .O(gate420inter7));
  inv1  gate1969(.a(G1132), .O(gate420inter8));
  nand2 gate1970(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1971(.a(s_203), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1972(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1973(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1974(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1457(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1458(.a(gate422inter0), .b(s_130), .O(gate422inter1));
  and2  gate1459(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1460(.a(s_130), .O(gate422inter3));
  inv1  gate1461(.a(s_131), .O(gate422inter4));
  nand2 gate1462(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1463(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1464(.a(G1039), .O(gate422inter7));
  inv1  gate1465(.a(G1135), .O(gate422inter8));
  nand2 gate1466(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1467(.a(s_131), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1468(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1469(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1470(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate589(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate590(.a(gate430inter0), .b(s_6), .O(gate430inter1));
  and2  gate591(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate592(.a(s_6), .O(gate430inter3));
  inv1  gate593(.a(s_7), .O(gate430inter4));
  nand2 gate594(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate595(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate596(.a(G1051), .O(gate430inter7));
  inv1  gate597(.a(G1147), .O(gate430inter8));
  nand2 gate598(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate599(.a(s_7), .b(gate430inter3), .O(gate430inter10));
  nor2  gate600(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate601(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate602(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1877(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1878(.a(gate432inter0), .b(s_190), .O(gate432inter1));
  and2  gate1879(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1880(.a(s_190), .O(gate432inter3));
  inv1  gate1881(.a(s_191), .O(gate432inter4));
  nand2 gate1882(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1883(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1884(.a(G1054), .O(gate432inter7));
  inv1  gate1885(.a(G1150), .O(gate432inter8));
  nand2 gate1886(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1887(.a(s_191), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1888(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1889(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1890(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1695(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1696(.a(gate441inter0), .b(s_164), .O(gate441inter1));
  and2  gate1697(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1698(.a(s_164), .O(gate441inter3));
  inv1  gate1699(.a(s_165), .O(gate441inter4));
  nand2 gate1700(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1701(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1702(.a(G12), .O(gate441inter7));
  inv1  gate1703(.a(G1165), .O(gate441inter8));
  nand2 gate1704(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1705(.a(s_165), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1706(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1707(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1708(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate841(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate842(.a(gate445inter0), .b(s_42), .O(gate445inter1));
  and2  gate843(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate844(.a(s_42), .O(gate445inter3));
  inv1  gate845(.a(s_43), .O(gate445inter4));
  nand2 gate846(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate847(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate848(.a(G14), .O(gate445inter7));
  inv1  gate849(.a(G1171), .O(gate445inter8));
  nand2 gate850(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate851(.a(s_43), .b(gate445inter3), .O(gate445inter10));
  nor2  gate852(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate853(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate854(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate687(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate688(.a(gate451inter0), .b(s_20), .O(gate451inter1));
  and2  gate689(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate690(.a(s_20), .O(gate451inter3));
  inv1  gate691(.a(s_21), .O(gate451inter4));
  nand2 gate692(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate693(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate694(.a(G17), .O(gate451inter7));
  inv1  gate695(.a(G1180), .O(gate451inter8));
  nand2 gate696(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate697(.a(s_21), .b(gate451inter3), .O(gate451inter10));
  nor2  gate698(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate699(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate700(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate981(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate982(.a(gate455inter0), .b(s_62), .O(gate455inter1));
  and2  gate983(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate984(.a(s_62), .O(gate455inter3));
  inv1  gate985(.a(s_63), .O(gate455inter4));
  nand2 gate986(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate987(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate988(.a(G19), .O(gate455inter7));
  inv1  gate989(.a(G1186), .O(gate455inter8));
  nand2 gate990(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate991(.a(s_63), .b(gate455inter3), .O(gate455inter10));
  nor2  gate992(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate993(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate994(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1793(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1794(.a(gate470inter0), .b(s_178), .O(gate470inter1));
  and2  gate1795(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1796(.a(s_178), .O(gate470inter3));
  inv1  gate1797(.a(s_179), .O(gate470inter4));
  nand2 gate1798(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1799(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1800(.a(G1111), .O(gate470inter7));
  inv1  gate1801(.a(G1207), .O(gate470inter8));
  nand2 gate1802(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1803(.a(s_179), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1804(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1805(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1806(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1177(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1178(.a(gate472inter0), .b(s_90), .O(gate472inter1));
  and2  gate1179(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1180(.a(s_90), .O(gate472inter3));
  inv1  gate1181(.a(s_91), .O(gate472inter4));
  nand2 gate1182(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1183(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1184(.a(G1114), .O(gate472inter7));
  inv1  gate1185(.a(G1210), .O(gate472inter8));
  nand2 gate1186(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1187(.a(s_91), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1188(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1189(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1190(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1009(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1010(.a(gate480inter0), .b(s_66), .O(gate480inter1));
  and2  gate1011(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1012(.a(s_66), .O(gate480inter3));
  inv1  gate1013(.a(s_67), .O(gate480inter4));
  nand2 gate1014(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1015(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1016(.a(G1126), .O(gate480inter7));
  inv1  gate1017(.a(G1222), .O(gate480inter8));
  nand2 gate1018(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1019(.a(s_67), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1020(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1021(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1022(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1513(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1514(.a(gate481inter0), .b(s_138), .O(gate481inter1));
  and2  gate1515(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1516(.a(s_138), .O(gate481inter3));
  inv1  gate1517(.a(s_139), .O(gate481inter4));
  nand2 gate1518(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1519(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1520(.a(G32), .O(gate481inter7));
  inv1  gate1521(.a(G1225), .O(gate481inter8));
  nand2 gate1522(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1523(.a(s_139), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1524(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1525(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1526(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1597(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1598(.a(gate482inter0), .b(s_150), .O(gate482inter1));
  and2  gate1599(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1600(.a(s_150), .O(gate482inter3));
  inv1  gate1601(.a(s_151), .O(gate482inter4));
  nand2 gate1602(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1603(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1604(.a(G1129), .O(gate482inter7));
  inv1  gate1605(.a(G1225), .O(gate482inter8));
  nand2 gate1606(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1607(.a(s_151), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1608(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1609(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1610(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate883(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate884(.a(gate484inter0), .b(s_48), .O(gate484inter1));
  and2  gate885(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate886(.a(s_48), .O(gate484inter3));
  inv1  gate887(.a(s_49), .O(gate484inter4));
  nand2 gate888(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate889(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate890(.a(G1230), .O(gate484inter7));
  inv1  gate891(.a(G1231), .O(gate484inter8));
  nand2 gate892(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate893(.a(s_49), .b(gate484inter3), .O(gate484inter10));
  nor2  gate894(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate895(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate896(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1415(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1416(.a(gate486inter0), .b(s_124), .O(gate486inter1));
  and2  gate1417(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1418(.a(s_124), .O(gate486inter3));
  inv1  gate1419(.a(s_125), .O(gate486inter4));
  nand2 gate1420(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1421(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1422(.a(G1234), .O(gate486inter7));
  inv1  gate1423(.a(G1235), .O(gate486inter8));
  nand2 gate1424(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1425(.a(s_125), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1426(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1427(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1428(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1653(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1654(.a(gate489inter0), .b(s_158), .O(gate489inter1));
  and2  gate1655(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1656(.a(s_158), .O(gate489inter3));
  inv1  gate1657(.a(s_159), .O(gate489inter4));
  nand2 gate1658(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1659(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1660(.a(G1240), .O(gate489inter7));
  inv1  gate1661(.a(G1241), .O(gate489inter8));
  nand2 gate1662(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1663(.a(s_159), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1664(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1665(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1666(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate855(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate856(.a(gate493inter0), .b(s_44), .O(gate493inter1));
  and2  gate857(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate858(.a(s_44), .O(gate493inter3));
  inv1  gate859(.a(s_45), .O(gate493inter4));
  nand2 gate860(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate861(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate862(.a(G1248), .O(gate493inter7));
  inv1  gate863(.a(G1249), .O(gate493inter8));
  nand2 gate864(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate865(.a(s_45), .b(gate493inter3), .O(gate493inter10));
  nor2  gate866(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate867(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate868(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1261(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1262(.a(gate499inter0), .b(s_102), .O(gate499inter1));
  and2  gate1263(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1264(.a(s_102), .O(gate499inter3));
  inv1  gate1265(.a(s_103), .O(gate499inter4));
  nand2 gate1266(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1267(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1268(.a(G1260), .O(gate499inter7));
  inv1  gate1269(.a(G1261), .O(gate499inter8));
  nand2 gate1270(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1271(.a(s_103), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1272(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1273(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1274(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate967(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate968(.a(gate504inter0), .b(s_60), .O(gate504inter1));
  and2  gate969(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate970(.a(s_60), .O(gate504inter3));
  inv1  gate971(.a(s_61), .O(gate504inter4));
  nand2 gate972(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate973(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate974(.a(G1270), .O(gate504inter7));
  inv1  gate975(.a(G1271), .O(gate504inter8));
  nand2 gate976(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate977(.a(s_61), .b(gate504inter3), .O(gate504inter10));
  nor2  gate978(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate979(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate980(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate547(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate548(.a(gate505inter0), .b(s_0), .O(gate505inter1));
  and2  gate549(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate550(.a(s_0), .O(gate505inter3));
  inv1  gate551(.a(s_1), .O(gate505inter4));
  nand2 gate552(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate553(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate554(.a(G1272), .O(gate505inter7));
  inv1  gate555(.a(G1273), .O(gate505inter8));
  nand2 gate556(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate557(.a(s_1), .b(gate505inter3), .O(gate505inter10));
  nor2  gate558(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate559(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate560(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1107(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1108(.a(gate509inter0), .b(s_80), .O(gate509inter1));
  and2  gate1109(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1110(.a(s_80), .O(gate509inter3));
  inv1  gate1111(.a(s_81), .O(gate509inter4));
  nand2 gate1112(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1113(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1114(.a(G1280), .O(gate509inter7));
  inv1  gate1115(.a(G1281), .O(gate509inter8));
  nand2 gate1116(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1117(.a(s_81), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1118(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1119(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1120(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1569(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1570(.a(gate510inter0), .b(s_146), .O(gate510inter1));
  and2  gate1571(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1572(.a(s_146), .O(gate510inter3));
  inv1  gate1573(.a(s_147), .O(gate510inter4));
  nand2 gate1574(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1575(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1576(.a(G1282), .O(gate510inter7));
  inv1  gate1577(.a(G1283), .O(gate510inter8));
  nand2 gate1578(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1579(.a(s_147), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1580(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1581(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1582(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1135(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1136(.a(gate511inter0), .b(s_84), .O(gate511inter1));
  and2  gate1137(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1138(.a(s_84), .O(gate511inter3));
  inv1  gate1139(.a(s_85), .O(gate511inter4));
  nand2 gate1140(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1141(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1142(.a(G1284), .O(gate511inter7));
  inv1  gate1143(.a(G1285), .O(gate511inter8));
  nand2 gate1144(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1145(.a(s_85), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1146(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1147(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1148(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1373(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1374(.a(gate514inter0), .b(s_118), .O(gate514inter1));
  and2  gate1375(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1376(.a(s_118), .O(gate514inter3));
  inv1  gate1377(.a(s_119), .O(gate514inter4));
  nand2 gate1378(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1379(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1380(.a(G1290), .O(gate514inter7));
  inv1  gate1381(.a(G1291), .O(gate514inter8));
  nand2 gate1382(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1383(.a(s_119), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1384(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1385(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1386(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule