module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1555(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1556(.a(gate12inter0), .b(s_144), .O(gate12inter1));
  and2  gate1557(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1558(.a(s_144), .O(gate12inter3));
  inv1  gate1559(.a(s_145), .O(gate12inter4));
  nand2 gate1560(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1561(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1562(.a(G7), .O(gate12inter7));
  inv1  gate1563(.a(G8), .O(gate12inter8));
  nand2 gate1564(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1565(.a(s_145), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1566(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1567(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1568(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate883(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate884(.a(gate13inter0), .b(s_48), .O(gate13inter1));
  and2  gate885(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate886(.a(s_48), .O(gate13inter3));
  inv1  gate887(.a(s_49), .O(gate13inter4));
  nand2 gate888(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate889(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate890(.a(G9), .O(gate13inter7));
  inv1  gate891(.a(G10), .O(gate13inter8));
  nand2 gate892(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate893(.a(s_49), .b(gate13inter3), .O(gate13inter10));
  nor2  gate894(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate895(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate896(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1569(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1570(.a(gate15inter0), .b(s_146), .O(gate15inter1));
  and2  gate1571(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1572(.a(s_146), .O(gate15inter3));
  inv1  gate1573(.a(s_147), .O(gate15inter4));
  nand2 gate1574(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1575(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1576(.a(G13), .O(gate15inter7));
  inv1  gate1577(.a(G14), .O(gate15inter8));
  nand2 gate1578(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1579(.a(s_147), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1580(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1581(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1582(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2269(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2270(.a(gate16inter0), .b(s_246), .O(gate16inter1));
  and2  gate2271(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2272(.a(s_246), .O(gate16inter3));
  inv1  gate2273(.a(s_247), .O(gate16inter4));
  nand2 gate2274(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2275(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2276(.a(G15), .O(gate16inter7));
  inv1  gate2277(.a(G16), .O(gate16inter8));
  nand2 gate2278(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2279(.a(s_247), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2280(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2281(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2282(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2563(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2564(.a(gate17inter0), .b(s_288), .O(gate17inter1));
  and2  gate2565(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2566(.a(s_288), .O(gate17inter3));
  inv1  gate2567(.a(s_289), .O(gate17inter4));
  nand2 gate2568(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2569(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2570(.a(G17), .O(gate17inter7));
  inv1  gate2571(.a(G18), .O(gate17inter8));
  nand2 gate2572(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2573(.a(s_289), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2574(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2575(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2576(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1751(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1752(.a(gate19inter0), .b(s_172), .O(gate19inter1));
  and2  gate1753(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1754(.a(s_172), .O(gate19inter3));
  inv1  gate1755(.a(s_173), .O(gate19inter4));
  nand2 gate1756(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1757(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1758(.a(G21), .O(gate19inter7));
  inv1  gate1759(.a(G22), .O(gate19inter8));
  nand2 gate1760(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1761(.a(s_173), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1762(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1763(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1764(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2493(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2494(.a(gate20inter0), .b(s_278), .O(gate20inter1));
  and2  gate2495(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2496(.a(s_278), .O(gate20inter3));
  inv1  gate2497(.a(s_279), .O(gate20inter4));
  nand2 gate2498(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2499(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2500(.a(G23), .O(gate20inter7));
  inv1  gate2501(.a(G24), .O(gate20inter8));
  nand2 gate2502(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2503(.a(s_279), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2504(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2505(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2506(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1401(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1402(.a(gate26inter0), .b(s_122), .O(gate26inter1));
  and2  gate1403(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1404(.a(s_122), .O(gate26inter3));
  inv1  gate1405(.a(s_123), .O(gate26inter4));
  nand2 gate1406(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1407(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1408(.a(G9), .O(gate26inter7));
  inv1  gate1409(.a(G13), .O(gate26inter8));
  nand2 gate1410(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1411(.a(s_123), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1412(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1413(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1414(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2101(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2102(.a(gate29inter0), .b(s_222), .O(gate29inter1));
  and2  gate2103(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2104(.a(s_222), .O(gate29inter3));
  inv1  gate2105(.a(s_223), .O(gate29inter4));
  nand2 gate2106(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2107(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2108(.a(G3), .O(gate29inter7));
  inv1  gate2109(.a(G7), .O(gate29inter8));
  nand2 gate2110(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2111(.a(s_223), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2112(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2113(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2114(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2577(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2578(.a(gate31inter0), .b(s_290), .O(gate31inter1));
  and2  gate2579(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2580(.a(s_290), .O(gate31inter3));
  inv1  gate2581(.a(s_291), .O(gate31inter4));
  nand2 gate2582(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2583(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2584(.a(G4), .O(gate31inter7));
  inv1  gate2585(.a(G8), .O(gate31inter8));
  nand2 gate2586(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2587(.a(s_291), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2588(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2589(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2590(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1583(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1584(.a(gate33inter0), .b(s_148), .O(gate33inter1));
  and2  gate1585(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1586(.a(s_148), .O(gate33inter3));
  inv1  gate1587(.a(s_149), .O(gate33inter4));
  nand2 gate1588(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1589(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1590(.a(G17), .O(gate33inter7));
  inv1  gate1591(.a(G21), .O(gate33inter8));
  nand2 gate1592(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1593(.a(s_149), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1594(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1595(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1596(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2059(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2060(.a(gate38inter0), .b(s_216), .O(gate38inter1));
  and2  gate2061(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2062(.a(s_216), .O(gate38inter3));
  inv1  gate2063(.a(s_217), .O(gate38inter4));
  nand2 gate2064(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2065(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2066(.a(G27), .O(gate38inter7));
  inv1  gate2067(.a(G31), .O(gate38inter8));
  nand2 gate2068(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2069(.a(s_217), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2070(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2071(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2072(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1121(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1122(.a(gate40inter0), .b(s_82), .O(gate40inter1));
  and2  gate1123(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1124(.a(s_82), .O(gate40inter3));
  inv1  gate1125(.a(s_83), .O(gate40inter4));
  nand2 gate1126(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1127(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1128(.a(G28), .O(gate40inter7));
  inv1  gate1129(.a(G32), .O(gate40inter8));
  nand2 gate1130(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1131(.a(s_83), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1132(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1133(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1134(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate715(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate716(.a(gate42inter0), .b(s_24), .O(gate42inter1));
  and2  gate717(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate718(.a(s_24), .O(gate42inter3));
  inv1  gate719(.a(s_25), .O(gate42inter4));
  nand2 gate720(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate721(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate722(.a(G2), .O(gate42inter7));
  inv1  gate723(.a(G266), .O(gate42inter8));
  nand2 gate724(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate725(.a(s_25), .b(gate42inter3), .O(gate42inter10));
  nor2  gate726(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate727(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate728(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1597(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1598(.a(gate43inter0), .b(s_150), .O(gate43inter1));
  and2  gate1599(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1600(.a(s_150), .O(gate43inter3));
  inv1  gate1601(.a(s_151), .O(gate43inter4));
  nand2 gate1602(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1603(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1604(.a(G3), .O(gate43inter7));
  inv1  gate1605(.a(G269), .O(gate43inter8));
  nand2 gate1606(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1607(.a(s_151), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1608(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1609(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1610(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate925(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate926(.a(gate46inter0), .b(s_54), .O(gate46inter1));
  and2  gate927(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate928(.a(s_54), .O(gate46inter3));
  inv1  gate929(.a(s_55), .O(gate46inter4));
  nand2 gate930(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate931(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate932(.a(G6), .O(gate46inter7));
  inv1  gate933(.a(G272), .O(gate46inter8));
  nand2 gate934(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate935(.a(s_55), .b(gate46inter3), .O(gate46inter10));
  nor2  gate936(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate937(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate938(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1345(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1346(.a(gate55inter0), .b(s_114), .O(gate55inter1));
  and2  gate1347(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1348(.a(s_114), .O(gate55inter3));
  inv1  gate1349(.a(s_115), .O(gate55inter4));
  nand2 gate1350(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1351(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1352(.a(G15), .O(gate55inter7));
  inv1  gate1353(.a(G287), .O(gate55inter8));
  nand2 gate1354(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1355(.a(s_115), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1356(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1357(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1358(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2451(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2452(.a(gate59inter0), .b(s_272), .O(gate59inter1));
  and2  gate2453(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2454(.a(s_272), .O(gate59inter3));
  inv1  gate2455(.a(s_273), .O(gate59inter4));
  nand2 gate2456(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2457(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2458(.a(G19), .O(gate59inter7));
  inv1  gate2459(.a(G293), .O(gate59inter8));
  nand2 gate2460(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2461(.a(s_273), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2462(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2463(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2464(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1471(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1472(.a(gate61inter0), .b(s_132), .O(gate61inter1));
  and2  gate1473(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1474(.a(s_132), .O(gate61inter3));
  inv1  gate1475(.a(s_133), .O(gate61inter4));
  nand2 gate1476(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1477(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1478(.a(G21), .O(gate61inter7));
  inv1  gate1479(.a(G296), .O(gate61inter8));
  nand2 gate1480(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1481(.a(s_133), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1482(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1483(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1484(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate2255(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2256(.a(gate63inter0), .b(s_244), .O(gate63inter1));
  and2  gate2257(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2258(.a(s_244), .O(gate63inter3));
  inv1  gate2259(.a(s_245), .O(gate63inter4));
  nand2 gate2260(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2261(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2262(.a(G23), .O(gate63inter7));
  inv1  gate2263(.a(G299), .O(gate63inter8));
  nand2 gate2264(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2265(.a(s_245), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2266(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2267(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2268(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1625(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1626(.a(gate64inter0), .b(s_154), .O(gate64inter1));
  and2  gate1627(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1628(.a(s_154), .O(gate64inter3));
  inv1  gate1629(.a(s_155), .O(gate64inter4));
  nand2 gate1630(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1631(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1632(.a(G24), .O(gate64inter7));
  inv1  gate1633(.a(G299), .O(gate64inter8));
  nand2 gate1634(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1635(.a(s_155), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1636(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1637(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1638(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1611(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1612(.a(gate65inter0), .b(s_152), .O(gate65inter1));
  and2  gate1613(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1614(.a(s_152), .O(gate65inter3));
  inv1  gate1615(.a(s_153), .O(gate65inter4));
  nand2 gate1616(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1617(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1618(.a(G25), .O(gate65inter7));
  inv1  gate1619(.a(G302), .O(gate65inter8));
  nand2 gate1620(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1621(.a(s_153), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1622(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1623(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1624(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1723(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1724(.a(gate67inter0), .b(s_168), .O(gate67inter1));
  and2  gate1725(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1726(.a(s_168), .O(gate67inter3));
  inv1  gate1727(.a(s_169), .O(gate67inter4));
  nand2 gate1728(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1729(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1730(.a(G27), .O(gate67inter7));
  inv1  gate1731(.a(G305), .O(gate67inter8));
  nand2 gate1732(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1733(.a(s_169), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1734(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1735(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1736(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1247(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1248(.a(gate68inter0), .b(s_100), .O(gate68inter1));
  and2  gate1249(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1250(.a(s_100), .O(gate68inter3));
  inv1  gate1251(.a(s_101), .O(gate68inter4));
  nand2 gate1252(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1253(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1254(.a(G28), .O(gate68inter7));
  inv1  gate1255(.a(G305), .O(gate68inter8));
  nand2 gate1256(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1257(.a(s_101), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1258(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1259(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1260(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate1359(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1360(.a(gate69inter0), .b(s_116), .O(gate69inter1));
  and2  gate1361(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1362(.a(s_116), .O(gate69inter3));
  inv1  gate1363(.a(s_117), .O(gate69inter4));
  nand2 gate1364(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1365(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1366(.a(G29), .O(gate69inter7));
  inv1  gate1367(.a(G308), .O(gate69inter8));
  nand2 gate1368(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1369(.a(s_117), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1370(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1371(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1372(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2325(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2326(.a(gate72inter0), .b(s_254), .O(gate72inter1));
  and2  gate2327(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2328(.a(s_254), .O(gate72inter3));
  inv1  gate2329(.a(s_255), .O(gate72inter4));
  nand2 gate2330(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2331(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2332(.a(G32), .O(gate72inter7));
  inv1  gate2333(.a(G311), .O(gate72inter8));
  nand2 gate2334(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2335(.a(s_255), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2336(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2337(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2338(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate561(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate562(.a(gate73inter0), .b(s_2), .O(gate73inter1));
  and2  gate563(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate564(.a(s_2), .O(gate73inter3));
  inv1  gate565(.a(s_3), .O(gate73inter4));
  nand2 gate566(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate567(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate568(.a(G1), .O(gate73inter7));
  inv1  gate569(.a(G314), .O(gate73inter8));
  nand2 gate570(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate571(.a(s_3), .b(gate73inter3), .O(gate73inter10));
  nor2  gate572(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate573(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate574(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate827(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate828(.a(gate75inter0), .b(s_40), .O(gate75inter1));
  and2  gate829(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate830(.a(s_40), .O(gate75inter3));
  inv1  gate831(.a(s_41), .O(gate75inter4));
  nand2 gate832(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate833(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate834(.a(G9), .O(gate75inter7));
  inv1  gate835(.a(G317), .O(gate75inter8));
  nand2 gate836(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate837(.a(s_41), .b(gate75inter3), .O(gate75inter10));
  nor2  gate838(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate839(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate840(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate645(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate646(.a(gate77inter0), .b(s_14), .O(gate77inter1));
  and2  gate647(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate648(.a(s_14), .O(gate77inter3));
  inv1  gate649(.a(s_15), .O(gate77inter4));
  nand2 gate650(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate651(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate652(.a(G2), .O(gate77inter7));
  inv1  gate653(.a(G320), .O(gate77inter8));
  nand2 gate654(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate655(.a(s_15), .b(gate77inter3), .O(gate77inter10));
  nor2  gate656(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate657(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate658(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate981(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate982(.a(gate78inter0), .b(s_62), .O(gate78inter1));
  and2  gate983(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate984(.a(s_62), .O(gate78inter3));
  inv1  gate985(.a(s_63), .O(gate78inter4));
  nand2 gate986(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate987(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate988(.a(G6), .O(gate78inter7));
  inv1  gate989(.a(G320), .O(gate78inter8));
  nand2 gate990(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate991(.a(s_63), .b(gate78inter3), .O(gate78inter10));
  nor2  gate992(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate993(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate994(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1527(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1528(.a(gate80inter0), .b(s_140), .O(gate80inter1));
  and2  gate1529(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1530(.a(s_140), .O(gate80inter3));
  inv1  gate1531(.a(s_141), .O(gate80inter4));
  nand2 gate1532(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1533(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1534(.a(G14), .O(gate80inter7));
  inv1  gate1535(.a(G323), .O(gate80inter8));
  nand2 gate1536(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1537(.a(s_141), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1538(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1539(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1540(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1541(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1542(.a(gate81inter0), .b(s_142), .O(gate81inter1));
  and2  gate1543(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1544(.a(s_142), .O(gate81inter3));
  inv1  gate1545(.a(s_143), .O(gate81inter4));
  nand2 gate1546(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1547(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1548(.a(G3), .O(gate81inter7));
  inv1  gate1549(.a(G326), .O(gate81inter8));
  nand2 gate1550(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1551(.a(s_143), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1552(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1553(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1554(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2241(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2242(.a(gate86inter0), .b(s_242), .O(gate86inter1));
  and2  gate2243(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2244(.a(s_242), .O(gate86inter3));
  inv1  gate2245(.a(s_243), .O(gate86inter4));
  nand2 gate2246(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2247(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2248(.a(G8), .O(gate86inter7));
  inv1  gate2249(.a(G332), .O(gate86inter8));
  nand2 gate2250(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2251(.a(s_243), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2252(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2253(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2254(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2521(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2522(.a(gate88inter0), .b(s_282), .O(gate88inter1));
  and2  gate2523(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2524(.a(s_282), .O(gate88inter3));
  inv1  gate2525(.a(s_283), .O(gate88inter4));
  nand2 gate2526(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2527(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2528(.a(G16), .O(gate88inter7));
  inv1  gate2529(.a(G335), .O(gate88inter8));
  nand2 gate2530(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2531(.a(s_283), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2532(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2533(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2534(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1107(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1108(.a(gate89inter0), .b(s_80), .O(gate89inter1));
  and2  gate1109(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1110(.a(s_80), .O(gate89inter3));
  inv1  gate1111(.a(s_81), .O(gate89inter4));
  nand2 gate1112(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1113(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1114(.a(G17), .O(gate89inter7));
  inv1  gate1115(.a(G338), .O(gate89inter8));
  nand2 gate1116(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1117(.a(s_81), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1118(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1119(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1120(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate2157(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2158(.a(gate90inter0), .b(s_230), .O(gate90inter1));
  and2  gate2159(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2160(.a(s_230), .O(gate90inter3));
  inv1  gate2161(.a(s_231), .O(gate90inter4));
  nand2 gate2162(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2163(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2164(.a(G21), .O(gate90inter7));
  inv1  gate2165(.a(G338), .O(gate90inter8));
  nand2 gate2166(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2167(.a(s_231), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2168(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2169(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2170(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1415(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1416(.a(gate92inter0), .b(s_124), .O(gate92inter1));
  and2  gate1417(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1418(.a(s_124), .O(gate92inter3));
  inv1  gate1419(.a(s_125), .O(gate92inter4));
  nand2 gate1420(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1421(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1422(.a(G29), .O(gate92inter7));
  inv1  gate1423(.a(G341), .O(gate92inter8));
  nand2 gate1424(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1425(.a(s_125), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1426(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1427(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1428(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1135(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1136(.a(gate97inter0), .b(s_84), .O(gate97inter1));
  and2  gate1137(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1138(.a(s_84), .O(gate97inter3));
  inv1  gate1139(.a(s_85), .O(gate97inter4));
  nand2 gate1140(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1141(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1142(.a(G19), .O(gate97inter7));
  inv1  gate1143(.a(G350), .O(gate97inter8));
  nand2 gate1144(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1145(.a(s_85), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1146(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1147(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1148(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate729(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate730(.a(gate98inter0), .b(s_26), .O(gate98inter1));
  and2  gate731(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate732(.a(s_26), .O(gate98inter3));
  inv1  gate733(.a(s_27), .O(gate98inter4));
  nand2 gate734(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate735(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate736(.a(G23), .O(gate98inter7));
  inv1  gate737(.a(G350), .O(gate98inter8));
  nand2 gate738(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate739(.a(s_27), .b(gate98inter3), .O(gate98inter10));
  nor2  gate740(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate741(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate742(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate659(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate660(.a(gate99inter0), .b(s_16), .O(gate99inter1));
  and2  gate661(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate662(.a(s_16), .O(gate99inter3));
  inv1  gate663(.a(s_17), .O(gate99inter4));
  nand2 gate664(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate665(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate666(.a(G27), .O(gate99inter7));
  inv1  gate667(.a(G353), .O(gate99inter8));
  nand2 gate668(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate669(.a(s_17), .b(gate99inter3), .O(gate99inter10));
  nor2  gate670(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate671(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate672(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2479(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2480(.a(gate102inter0), .b(s_276), .O(gate102inter1));
  and2  gate2481(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2482(.a(s_276), .O(gate102inter3));
  inv1  gate2483(.a(s_277), .O(gate102inter4));
  nand2 gate2484(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2485(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2486(.a(G24), .O(gate102inter7));
  inv1  gate2487(.a(G356), .O(gate102inter8));
  nand2 gate2488(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2489(.a(s_277), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2490(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2491(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2492(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate939(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate940(.a(gate104inter0), .b(s_56), .O(gate104inter1));
  and2  gate941(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate942(.a(s_56), .O(gate104inter3));
  inv1  gate943(.a(s_57), .O(gate104inter4));
  nand2 gate944(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate945(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate946(.a(G32), .O(gate104inter7));
  inv1  gate947(.a(G359), .O(gate104inter8));
  nand2 gate948(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate949(.a(s_57), .b(gate104inter3), .O(gate104inter10));
  nor2  gate950(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate951(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate952(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2339(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2340(.a(gate107inter0), .b(s_256), .O(gate107inter1));
  and2  gate2341(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2342(.a(s_256), .O(gate107inter3));
  inv1  gate2343(.a(s_257), .O(gate107inter4));
  nand2 gate2344(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2345(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2346(.a(G366), .O(gate107inter7));
  inv1  gate2347(.a(G367), .O(gate107inter8));
  nand2 gate2348(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2349(.a(s_257), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2350(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2351(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2352(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate2311(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2312(.a(gate108inter0), .b(s_252), .O(gate108inter1));
  and2  gate2313(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2314(.a(s_252), .O(gate108inter3));
  inv1  gate2315(.a(s_253), .O(gate108inter4));
  nand2 gate2316(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2317(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2318(.a(G368), .O(gate108inter7));
  inv1  gate2319(.a(G369), .O(gate108inter8));
  nand2 gate2320(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2321(.a(s_253), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2322(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2323(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2324(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1905(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1906(.a(gate110inter0), .b(s_194), .O(gate110inter1));
  and2  gate1907(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1908(.a(s_194), .O(gate110inter3));
  inv1  gate1909(.a(s_195), .O(gate110inter4));
  nand2 gate1910(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1911(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1912(.a(G372), .O(gate110inter7));
  inv1  gate1913(.a(G373), .O(gate110inter8));
  nand2 gate1914(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1915(.a(s_195), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1916(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1917(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1918(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1821(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1822(.a(gate111inter0), .b(s_182), .O(gate111inter1));
  and2  gate1823(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1824(.a(s_182), .O(gate111inter3));
  inv1  gate1825(.a(s_183), .O(gate111inter4));
  nand2 gate1826(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1827(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1828(.a(G374), .O(gate111inter7));
  inv1  gate1829(.a(G375), .O(gate111inter8));
  nand2 gate1830(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1831(.a(s_183), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1832(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1833(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1834(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1205(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1206(.a(gate112inter0), .b(s_94), .O(gate112inter1));
  and2  gate1207(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1208(.a(s_94), .O(gate112inter3));
  inv1  gate1209(.a(s_95), .O(gate112inter4));
  nand2 gate1210(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1211(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1212(.a(G376), .O(gate112inter7));
  inv1  gate1213(.a(G377), .O(gate112inter8));
  nand2 gate1214(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1215(.a(s_95), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1216(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1217(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1218(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1149(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1150(.a(gate114inter0), .b(s_86), .O(gate114inter1));
  and2  gate1151(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1152(.a(s_86), .O(gate114inter3));
  inv1  gate1153(.a(s_87), .O(gate114inter4));
  nand2 gate1154(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1155(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1156(.a(G380), .O(gate114inter7));
  inv1  gate1157(.a(G381), .O(gate114inter8));
  nand2 gate1158(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1159(.a(s_87), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1160(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1161(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1162(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1037(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1038(.a(gate116inter0), .b(s_70), .O(gate116inter1));
  and2  gate1039(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1040(.a(s_70), .O(gate116inter3));
  inv1  gate1041(.a(s_71), .O(gate116inter4));
  nand2 gate1042(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1043(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1044(.a(G384), .O(gate116inter7));
  inv1  gate1045(.a(G385), .O(gate116inter8));
  nand2 gate1046(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1047(.a(s_71), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1048(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1049(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1050(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2227(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2228(.a(gate119inter0), .b(s_240), .O(gate119inter1));
  and2  gate2229(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2230(.a(s_240), .O(gate119inter3));
  inv1  gate2231(.a(s_241), .O(gate119inter4));
  nand2 gate2232(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2233(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2234(.a(G390), .O(gate119inter7));
  inv1  gate2235(.a(G391), .O(gate119inter8));
  nand2 gate2236(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2237(.a(s_241), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2238(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2239(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2240(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1681(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1682(.a(gate132inter0), .b(s_162), .O(gate132inter1));
  and2  gate1683(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1684(.a(s_162), .O(gate132inter3));
  inv1  gate1685(.a(s_163), .O(gate132inter4));
  nand2 gate1686(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1687(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1688(.a(G416), .O(gate132inter7));
  inv1  gate1689(.a(G417), .O(gate132inter8));
  nand2 gate1690(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1691(.a(s_163), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1692(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1693(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1694(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2507(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2508(.a(gate136inter0), .b(s_280), .O(gate136inter1));
  and2  gate2509(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2510(.a(s_280), .O(gate136inter3));
  inv1  gate2511(.a(s_281), .O(gate136inter4));
  nand2 gate2512(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2513(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2514(.a(G424), .O(gate136inter7));
  inv1  gate2515(.a(G425), .O(gate136inter8));
  nand2 gate2516(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2517(.a(s_281), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2518(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2519(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2520(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2143(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2144(.a(gate139inter0), .b(s_228), .O(gate139inter1));
  and2  gate2145(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2146(.a(s_228), .O(gate139inter3));
  inv1  gate2147(.a(s_229), .O(gate139inter4));
  nand2 gate2148(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2149(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2150(.a(G438), .O(gate139inter7));
  inv1  gate2151(.a(G441), .O(gate139inter8));
  nand2 gate2152(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2153(.a(s_229), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2154(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2155(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2156(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1289(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1290(.a(gate142inter0), .b(s_106), .O(gate142inter1));
  and2  gate1291(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1292(.a(s_106), .O(gate142inter3));
  inv1  gate1293(.a(s_107), .O(gate142inter4));
  nand2 gate1294(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1295(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1296(.a(G456), .O(gate142inter7));
  inv1  gate1297(.a(G459), .O(gate142inter8));
  nand2 gate1298(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1299(.a(s_107), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1300(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1301(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1302(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate855(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate856(.a(gate146inter0), .b(s_44), .O(gate146inter1));
  and2  gate857(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate858(.a(s_44), .O(gate146inter3));
  inv1  gate859(.a(s_45), .O(gate146inter4));
  nand2 gate860(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate861(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate862(.a(G480), .O(gate146inter7));
  inv1  gate863(.a(G483), .O(gate146inter8));
  nand2 gate864(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate865(.a(s_45), .b(gate146inter3), .O(gate146inter10));
  nor2  gate866(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate867(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate868(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1079(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1080(.a(gate149inter0), .b(s_76), .O(gate149inter1));
  and2  gate1081(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1082(.a(s_76), .O(gate149inter3));
  inv1  gate1083(.a(s_77), .O(gate149inter4));
  nand2 gate1084(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1085(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1086(.a(G498), .O(gate149inter7));
  inv1  gate1087(.a(G501), .O(gate149inter8));
  nand2 gate1088(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1089(.a(s_77), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1090(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1091(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1092(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1695(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1696(.a(gate150inter0), .b(s_164), .O(gate150inter1));
  and2  gate1697(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1698(.a(s_164), .O(gate150inter3));
  inv1  gate1699(.a(s_165), .O(gate150inter4));
  nand2 gate1700(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1701(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1702(.a(G504), .O(gate150inter7));
  inv1  gate1703(.a(G507), .O(gate150inter8));
  nand2 gate1704(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1705(.a(s_165), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1706(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1707(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1708(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2549(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2550(.a(gate151inter0), .b(s_286), .O(gate151inter1));
  and2  gate2551(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2552(.a(s_286), .O(gate151inter3));
  inv1  gate2553(.a(s_287), .O(gate151inter4));
  nand2 gate2554(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2555(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2556(.a(G510), .O(gate151inter7));
  inv1  gate2557(.a(G513), .O(gate151inter8));
  nand2 gate2558(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2559(.a(s_287), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2560(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2561(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2562(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1485(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1486(.a(gate154inter0), .b(s_134), .O(gate154inter1));
  and2  gate1487(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1488(.a(s_134), .O(gate154inter3));
  inv1  gate1489(.a(s_135), .O(gate154inter4));
  nand2 gate1490(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1491(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1492(.a(G429), .O(gate154inter7));
  inv1  gate1493(.a(G522), .O(gate154inter8));
  nand2 gate1494(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1495(.a(s_135), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1496(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1497(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1498(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate589(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate590(.a(gate160inter0), .b(s_6), .O(gate160inter1));
  and2  gate591(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate592(.a(s_6), .O(gate160inter3));
  inv1  gate593(.a(s_7), .O(gate160inter4));
  nand2 gate594(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate595(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate596(.a(G447), .O(gate160inter7));
  inv1  gate597(.a(G531), .O(gate160inter8));
  nand2 gate598(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate599(.a(s_7), .b(gate160inter3), .O(gate160inter10));
  nor2  gate600(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate601(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate602(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate701(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate702(.a(gate163inter0), .b(s_22), .O(gate163inter1));
  and2  gate703(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate704(.a(s_22), .O(gate163inter3));
  inv1  gate705(.a(s_23), .O(gate163inter4));
  nand2 gate706(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate707(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate708(.a(G456), .O(gate163inter7));
  inv1  gate709(.a(G537), .O(gate163inter8));
  nand2 gate710(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate711(.a(s_23), .b(gate163inter3), .O(gate163inter10));
  nor2  gate712(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate713(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate714(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate785(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate786(.a(gate164inter0), .b(s_34), .O(gate164inter1));
  and2  gate787(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate788(.a(s_34), .O(gate164inter3));
  inv1  gate789(.a(s_35), .O(gate164inter4));
  nand2 gate790(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate791(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate792(.a(G459), .O(gate164inter7));
  inv1  gate793(.a(G537), .O(gate164inter8));
  nand2 gate794(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate795(.a(s_35), .b(gate164inter3), .O(gate164inter10));
  nor2  gate796(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate797(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate798(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate995(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate996(.a(gate165inter0), .b(s_64), .O(gate165inter1));
  and2  gate997(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate998(.a(s_64), .O(gate165inter3));
  inv1  gate999(.a(s_65), .O(gate165inter4));
  nand2 gate1000(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1001(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1002(.a(G462), .O(gate165inter7));
  inv1  gate1003(.a(G540), .O(gate165inter8));
  nand2 gate1004(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1005(.a(s_65), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1006(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1007(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1008(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1219(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1220(.a(gate167inter0), .b(s_96), .O(gate167inter1));
  and2  gate1221(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1222(.a(s_96), .O(gate167inter3));
  inv1  gate1223(.a(s_97), .O(gate167inter4));
  nand2 gate1224(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1225(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1226(.a(G468), .O(gate167inter7));
  inv1  gate1227(.a(G543), .O(gate167inter8));
  nand2 gate1228(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1229(.a(s_97), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1230(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1231(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1232(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate897(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate898(.a(gate176inter0), .b(s_50), .O(gate176inter1));
  and2  gate899(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate900(.a(s_50), .O(gate176inter3));
  inv1  gate901(.a(s_51), .O(gate176inter4));
  nand2 gate902(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate903(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate904(.a(G495), .O(gate176inter7));
  inv1  gate905(.a(G555), .O(gate176inter8));
  nand2 gate906(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate907(.a(s_51), .b(gate176inter3), .O(gate176inter10));
  nor2  gate908(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate909(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate910(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate617(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate618(.a(gate180inter0), .b(s_10), .O(gate180inter1));
  and2  gate619(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate620(.a(s_10), .O(gate180inter3));
  inv1  gate621(.a(s_11), .O(gate180inter4));
  nand2 gate622(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate623(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate624(.a(G507), .O(gate180inter7));
  inv1  gate625(.a(G561), .O(gate180inter8));
  nand2 gate626(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate627(.a(s_11), .b(gate180inter3), .O(gate180inter10));
  nor2  gate628(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate629(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate630(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate603(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate604(.a(gate186inter0), .b(s_8), .O(gate186inter1));
  and2  gate605(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate606(.a(s_8), .O(gate186inter3));
  inv1  gate607(.a(s_9), .O(gate186inter4));
  nand2 gate608(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate609(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate610(.a(G572), .O(gate186inter7));
  inv1  gate611(.a(G573), .O(gate186inter8));
  nand2 gate612(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate613(.a(s_9), .b(gate186inter3), .O(gate186inter10));
  nor2  gate614(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate615(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate616(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate841(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate842(.a(gate197inter0), .b(s_42), .O(gate197inter1));
  and2  gate843(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate844(.a(s_42), .O(gate197inter3));
  inv1  gate845(.a(s_43), .O(gate197inter4));
  nand2 gate846(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate847(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate848(.a(G594), .O(gate197inter7));
  inv1  gate849(.a(G595), .O(gate197inter8));
  nand2 gate850(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate851(.a(s_43), .b(gate197inter3), .O(gate197inter10));
  nor2  gate852(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate853(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate854(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1387(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1388(.a(gate200inter0), .b(s_120), .O(gate200inter1));
  and2  gate1389(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1390(.a(s_120), .O(gate200inter3));
  inv1  gate1391(.a(s_121), .O(gate200inter4));
  nand2 gate1392(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1393(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1394(.a(G600), .O(gate200inter7));
  inv1  gate1395(.a(G601), .O(gate200inter8));
  nand2 gate1396(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1397(.a(s_121), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1398(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1399(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1400(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1709(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1710(.a(gate202inter0), .b(s_166), .O(gate202inter1));
  and2  gate1711(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1712(.a(s_166), .O(gate202inter3));
  inv1  gate1713(.a(s_167), .O(gate202inter4));
  nand2 gate1714(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1715(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1716(.a(G612), .O(gate202inter7));
  inv1  gate1717(.a(G617), .O(gate202inter8));
  nand2 gate1718(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1719(.a(s_167), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1720(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1721(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1722(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1793(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1794(.a(gate203inter0), .b(s_178), .O(gate203inter1));
  and2  gate1795(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1796(.a(s_178), .O(gate203inter3));
  inv1  gate1797(.a(s_179), .O(gate203inter4));
  nand2 gate1798(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1799(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1800(.a(G602), .O(gate203inter7));
  inv1  gate1801(.a(G612), .O(gate203inter8));
  nand2 gate1802(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1803(.a(s_179), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1804(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1805(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1806(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2073(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2074(.a(gate205inter0), .b(s_218), .O(gate205inter1));
  and2  gate2075(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2076(.a(s_218), .O(gate205inter3));
  inv1  gate2077(.a(s_219), .O(gate205inter4));
  nand2 gate2078(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2079(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2080(.a(G622), .O(gate205inter7));
  inv1  gate2081(.a(G627), .O(gate205inter8));
  nand2 gate2082(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2083(.a(s_219), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2084(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2085(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2086(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate743(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate744(.a(gate213inter0), .b(s_28), .O(gate213inter1));
  and2  gate745(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate746(.a(s_28), .O(gate213inter3));
  inv1  gate747(.a(s_29), .O(gate213inter4));
  nand2 gate748(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate749(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate750(.a(G602), .O(gate213inter7));
  inv1  gate751(.a(G672), .O(gate213inter8));
  nand2 gate752(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate753(.a(s_29), .b(gate213inter3), .O(gate213inter10));
  nor2  gate754(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate755(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate756(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1877(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1878(.a(gate215inter0), .b(s_190), .O(gate215inter1));
  and2  gate1879(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1880(.a(s_190), .O(gate215inter3));
  inv1  gate1881(.a(s_191), .O(gate215inter4));
  nand2 gate1882(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1883(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1884(.a(G607), .O(gate215inter7));
  inv1  gate1885(.a(G675), .O(gate215inter8));
  nand2 gate1886(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1887(.a(s_191), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1888(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1889(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1890(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1331(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1332(.a(gate216inter0), .b(s_112), .O(gate216inter1));
  and2  gate1333(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1334(.a(s_112), .O(gate216inter3));
  inv1  gate1335(.a(s_113), .O(gate216inter4));
  nand2 gate1336(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1337(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1338(.a(G617), .O(gate216inter7));
  inv1  gate1339(.a(G675), .O(gate216inter8));
  nand2 gate1340(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1341(.a(s_113), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1342(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1343(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1344(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate869(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate870(.a(gate217inter0), .b(s_46), .O(gate217inter1));
  and2  gate871(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate872(.a(s_46), .O(gate217inter3));
  inv1  gate873(.a(s_47), .O(gate217inter4));
  nand2 gate874(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate875(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate876(.a(G622), .O(gate217inter7));
  inv1  gate877(.a(G678), .O(gate217inter8));
  nand2 gate878(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate879(.a(s_47), .b(gate217inter3), .O(gate217inter10));
  nor2  gate880(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate881(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate882(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2297(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2298(.a(gate219inter0), .b(s_250), .O(gate219inter1));
  and2  gate2299(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2300(.a(s_250), .O(gate219inter3));
  inv1  gate2301(.a(s_251), .O(gate219inter4));
  nand2 gate2302(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2303(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2304(.a(G632), .O(gate219inter7));
  inv1  gate2305(.a(G681), .O(gate219inter8));
  nand2 gate2306(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2307(.a(s_251), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2308(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2309(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2310(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2423(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2424(.a(gate222inter0), .b(s_268), .O(gate222inter1));
  and2  gate2425(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2426(.a(s_268), .O(gate222inter3));
  inv1  gate2427(.a(s_269), .O(gate222inter4));
  nand2 gate2428(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2429(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2430(.a(G632), .O(gate222inter7));
  inv1  gate2431(.a(G684), .O(gate222inter8));
  nand2 gate2432(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2433(.a(s_269), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2434(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2435(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2436(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate771(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate772(.a(gate230inter0), .b(s_32), .O(gate230inter1));
  and2  gate773(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate774(.a(s_32), .O(gate230inter3));
  inv1  gate775(.a(s_33), .O(gate230inter4));
  nand2 gate776(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate777(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate778(.a(G700), .O(gate230inter7));
  inv1  gate779(.a(G701), .O(gate230inter8));
  nand2 gate780(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate781(.a(s_33), .b(gate230inter3), .O(gate230inter10));
  nor2  gate782(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate783(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate784(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2115(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2116(.a(gate232inter0), .b(s_224), .O(gate232inter1));
  and2  gate2117(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2118(.a(s_224), .O(gate232inter3));
  inv1  gate2119(.a(s_225), .O(gate232inter4));
  nand2 gate2120(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2121(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2122(.a(G704), .O(gate232inter7));
  inv1  gate2123(.a(G705), .O(gate232inter8));
  nand2 gate2124(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2125(.a(s_225), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2126(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2127(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2128(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2381(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2382(.a(gate236inter0), .b(s_262), .O(gate236inter1));
  and2  gate2383(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2384(.a(s_262), .O(gate236inter3));
  inv1  gate2385(.a(s_263), .O(gate236inter4));
  nand2 gate2386(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2387(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2388(.a(G251), .O(gate236inter7));
  inv1  gate2389(.a(G727), .O(gate236inter8));
  nand2 gate2390(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2391(.a(s_263), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2392(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2393(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2394(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1737(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1738(.a(gate237inter0), .b(s_170), .O(gate237inter1));
  and2  gate1739(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1740(.a(s_170), .O(gate237inter3));
  inv1  gate1741(.a(s_171), .O(gate237inter4));
  nand2 gate1742(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1743(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1744(.a(G254), .O(gate237inter7));
  inv1  gate1745(.a(G706), .O(gate237inter8));
  nand2 gate1746(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1747(.a(s_171), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1748(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1749(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1750(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1667(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1668(.a(gate248inter0), .b(s_160), .O(gate248inter1));
  and2  gate1669(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1670(.a(s_160), .O(gate248inter3));
  inv1  gate1671(.a(s_161), .O(gate248inter4));
  nand2 gate1672(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1673(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1674(.a(G727), .O(gate248inter7));
  inv1  gate1675(.a(G739), .O(gate248inter8));
  nand2 gate1676(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1677(.a(s_161), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1678(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1679(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1680(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1933(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1934(.a(gate249inter0), .b(s_198), .O(gate249inter1));
  and2  gate1935(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1936(.a(s_198), .O(gate249inter3));
  inv1  gate1937(.a(s_199), .O(gate249inter4));
  nand2 gate1938(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1939(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1940(.a(G254), .O(gate249inter7));
  inv1  gate1941(.a(G742), .O(gate249inter8));
  nand2 gate1942(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1943(.a(s_199), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1944(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1945(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1946(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1807(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1808(.a(gate250inter0), .b(s_180), .O(gate250inter1));
  and2  gate1809(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1810(.a(s_180), .O(gate250inter3));
  inv1  gate1811(.a(s_181), .O(gate250inter4));
  nand2 gate1812(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1813(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1814(.a(G706), .O(gate250inter7));
  inv1  gate1815(.a(G742), .O(gate250inter8));
  nand2 gate1816(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1817(.a(s_181), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1818(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1819(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1820(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1919(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1920(.a(gate252inter0), .b(s_196), .O(gate252inter1));
  and2  gate1921(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1922(.a(s_196), .O(gate252inter3));
  inv1  gate1923(.a(s_197), .O(gate252inter4));
  nand2 gate1924(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1925(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1926(.a(G709), .O(gate252inter7));
  inv1  gate1927(.a(G745), .O(gate252inter8));
  nand2 gate1928(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1929(.a(s_197), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1930(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1931(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1932(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2409(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2410(.a(gate257inter0), .b(s_266), .O(gate257inter1));
  and2  gate2411(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2412(.a(s_266), .O(gate257inter3));
  inv1  gate2413(.a(s_267), .O(gate257inter4));
  nand2 gate2414(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2415(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2416(.a(G754), .O(gate257inter7));
  inv1  gate2417(.a(G755), .O(gate257inter8));
  nand2 gate2418(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2419(.a(s_267), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2420(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2421(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2422(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1261(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1262(.a(gate258inter0), .b(s_102), .O(gate258inter1));
  and2  gate1263(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1264(.a(s_102), .O(gate258inter3));
  inv1  gate1265(.a(s_103), .O(gate258inter4));
  nand2 gate1266(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1267(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1268(.a(G756), .O(gate258inter7));
  inv1  gate1269(.a(G757), .O(gate258inter8));
  nand2 gate1270(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1271(.a(s_103), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1272(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1273(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1274(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1191(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1192(.a(gate261inter0), .b(s_92), .O(gate261inter1));
  and2  gate1193(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1194(.a(s_92), .O(gate261inter3));
  inv1  gate1195(.a(s_93), .O(gate261inter4));
  nand2 gate1196(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1197(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1198(.a(G762), .O(gate261inter7));
  inv1  gate1199(.a(G763), .O(gate261inter8));
  nand2 gate1200(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1201(.a(s_93), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1202(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1203(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1204(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate953(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate954(.a(gate262inter0), .b(s_58), .O(gate262inter1));
  and2  gate955(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate956(.a(s_58), .O(gate262inter3));
  inv1  gate957(.a(s_59), .O(gate262inter4));
  nand2 gate958(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate959(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate960(.a(G764), .O(gate262inter7));
  inv1  gate961(.a(G765), .O(gate262inter8));
  nand2 gate962(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate963(.a(s_59), .b(gate262inter3), .O(gate262inter10));
  nor2  gate964(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate965(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate966(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1765(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1766(.a(gate267inter0), .b(s_174), .O(gate267inter1));
  and2  gate1767(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1768(.a(s_174), .O(gate267inter3));
  inv1  gate1769(.a(s_175), .O(gate267inter4));
  nand2 gate1770(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1771(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1772(.a(G648), .O(gate267inter7));
  inv1  gate1773(.a(G776), .O(gate267inter8));
  nand2 gate1774(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1775(.a(s_175), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1776(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1777(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1778(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1989(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1990(.a(gate268inter0), .b(s_206), .O(gate268inter1));
  and2  gate1991(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1992(.a(s_206), .O(gate268inter3));
  inv1  gate1993(.a(s_207), .O(gate268inter4));
  nand2 gate1994(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1995(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1996(.a(G651), .O(gate268inter7));
  inv1  gate1997(.a(G779), .O(gate268inter8));
  nand2 gate1998(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1999(.a(s_207), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2000(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2001(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2002(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2213(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2214(.a(gate269inter0), .b(s_238), .O(gate269inter1));
  and2  gate2215(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2216(.a(s_238), .O(gate269inter3));
  inv1  gate2217(.a(s_239), .O(gate269inter4));
  nand2 gate2218(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2219(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2220(.a(G654), .O(gate269inter7));
  inv1  gate2221(.a(G782), .O(gate269inter8));
  nand2 gate2222(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2223(.a(s_239), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2224(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2225(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2226(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1065(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1066(.a(gate276inter0), .b(s_74), .O(gate276inter1));
  and2  gate1067(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1068(.a(s_74), .O(gate276inter3));
  inv1  gate1069(.a(s_75), .O(gate276inter4));
  nand2 gate1070(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1071(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1072(.a(G773), .O(gate276inter7));
  inv1  gate1073(.a(G797), .O(gate276inter8));
  nand2 gate1074(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1075(.a(s_75), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1076(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1077(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1078(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2437(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2438(.a(gate278inter0), .b(s_270), .O(gate278inter1));
  and2  gate2439(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2440(.a(s_270), .O(gate278inter3));
  inv1  gate2441(.a(s_271), .O(gate278inter4));
  nand2 gate2442(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2443(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2444(.a(G776), .O(gate278inter7));
  inv1  gate2445(.a(G800), .O(gate278inter8));
  nand2 gate2446(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2447(.a(s_271), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2448(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2449(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2450(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate547(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate548(.a(gate279inter0), .b(s_0), .O(gate279inter1));
  and2  gate549(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate550(.a(s_0), .O(gate279inter3));
  inv1  gate551(.a(s_1), .O(gate279inter4));
  nand2 gate552(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate553(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate554(.a(G651), .O(gate279inter7));
  inv1  gate555(.a(G803), .O(gate279inter8));
  nand2 gate556(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate557(.a(s_1), .b(gate279inter3), .O(gate279inter10));
  nor2  gate558(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate559(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate560(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1023(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1024(.a(gate280inter0), .b(s_68), .O(gate280inter1));
  and2  gate1025(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1026(.a(s_68), .O(gate280inter3));
  inv1  gate1027(.a(s_69), .O(gate280inter4));
  nand2 gate1028(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1029(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1030(.a(G779), .O(gate280inter7));
  inv1  gate1031(.a(G803), .O(gate280inter8));
  nand2 gate1032(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1033(.a(s_69), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1034(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1035(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1036(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2017(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2018(.a(gate282inter0), .b(s_210), .O(gate282inter1));
  and2  gate2019(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2020(.a(s_210), .O(gate282inter3));
  inv1  gate2021(.a(s_211), .O(gate282inter4));
  nand2 gate2022(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2023(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2024(.a(G782), .O(gate282inter7));
  inv1  gate2025(.a(G806), .O(gate282inter8));
  nand2 gate2026(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2027(.a(s_211), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2028(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2029(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2030(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1513(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1514(.a(gate283inter0), .b(s_138), .O(gate283inter1));
  and2  gate1515(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1516(.a(s_138), .O(gate283inter3));
  inv1  gate1517(.a(s_139), .O(gate283inter4));
  nand2 gate1518(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1519(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1520(.a(G657), .O(gate283inter7));
  inv1  gate1521(.a(G809), .O(gate283inter8));
  nand2 gate1522(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1523(.a(s_139), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1524(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1525(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1526(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1499(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1500(.a(gate284inter0), .b(s_136), .O(gate284inter1));
  and2  gate1501(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1502(.a(s_136), .O(gate284inter3));
  inv1  gate1503(.a(s_137), .O(gate284inter4));
  nand2 gate1504(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1505(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1506(.a(G785), .O(gate284inter7));
  inv1  gate1507(.a(G809), .O(gate284inter8));
  nand2 gate1508(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1509(.a(s_137), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1510(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1511(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1512(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1835(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1836(.a(gate286inter0), .b(s_184), .O(gate286inter1));
  and2  gate1837(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1838(.a(s_184), .O(gate286inter3));
  inv1  gate1839(.a(s_185), .O(gate286inter4));
  nand2 gate1840(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1841(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1842(.a(G788), .O(gate286inter7));
  inv1  gate1843(.a(G812), .O(gate286inter8));
  nand2 gate1844(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1845(.a(s_185), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1846(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1847(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1848(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate799(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate800(.a(gate289inter0), .b(s_36), .O(gate289inter1));
  and2  gate801(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate802(.a(s_36), .O(gate289inter3));
  inv1  gate803(.a(s_37), .O(gate289inter4));
  nand2 gate804(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate805(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate806(.a(G818), .O(gate289inter7));
  inv1  gate807(.a(G819), .O(gate289inter8));
  nand2 gate808(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate809(.a(s_37), .b(gate289inter3), .O(gate289inter10));
  nor2  gate810(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate811(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate812(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1303(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1304(.a(gate290inter0), .b(s_108), .O(gate290inter1));
  and2  gate1305(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1306(.a(s_108), .O(gate290inter3));
  inv1  gate1307(.a(s_109), .O(gate290inter4));
  nand2 gate1308(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1309(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1310(.a(G820), .O(gate290inter7));
  inv1  gate1311(.a(G821), .O(gate290inter8));
  nand2 gate1312(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1313(.a(s_109), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1314(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1315(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1316(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2353(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2354(.a(gate293inter0), .b(s_258), .O(gate293inter1));
  and2  gate2355(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2356(.a(s_258), .O(gate293inter3));
  inv1  gate2357(.a(s_259), .O(gate293inter4));
  nand2 gate2358(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2359(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2360(.a(G828), .O(gate293inter7));
  inv1  gate2361(.a(G829), .O(gate293inter8));
  nand2 gate2362(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2363(.a(s_259), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2364(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2365(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2366(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2087(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2088(.a(gate295inter0), .b(s_220), .O(gate295inter1));
  and2  gate2089(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2090(.a(s_220), .O(gate295inter3));
  inv1  gate2091(.a(s_221), .O(gate295inter4));
  nand2 gate2092(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2093(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2094(.a(G830), .O(gate295inter7));
  inv1  gate2095(.a(G831), .O(gate295inter8));
  nand2 gate2096(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2097(.a(s_221), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2098(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2099(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2100(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1373(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1374(.a(gate388inter0), .b(s_118), .O(gate388inter1));
  and2  gate1375(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1376(.a(s_118), .O(gate388inter3));
  inv1  gate1377(.a(s_119), .O(gate388inter4));
  nand2 gate1378(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1379(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1380(.a(G2), .O(gate388inter7));
  inv1  gate1381(.a(G1039), .O(gate388inter8));
  nand2 gate1382(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1383(.a(s_119), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1384(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1385(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1386(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2199(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2200(.a(gate393inter0), .b(s_236), .O(gate393inter1));
  and2  gate2201(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2202(.a(s_236), .O(gate393inter3));
  inv1  gate2203(.a(s_237), .O(gate393inter4));
  nand2 gate2204(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2205(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2206(.a(G7), .O(gate393inter7));
  inv1  gate2207(.a(G1054), .O(gate393inter8));
  nand2 gate2208(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2209(.a(s_237), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2210(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2211(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2212(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate967(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate968(.a(gate399inter0), .b(s_60), .O(gate399inter1));
  and2  gate969(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate970(.a(s_60), .O(gate399inter3));
  inv1  gate971(.a(s_61), .O(gate399inter4));
  nand2 gate972(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate973(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate974(.a(G13), .O(gate399inter7));
  inv1  gate975(.a(G1072), .O(gate399inter8));
  nand2 gate976(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate977(.a(s_61), .b(gate399inter3), .O(gate399inter10));
  nor2  gate978(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate979(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate980(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1947(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1948(.a(gate407inter0), .b(s_200), .O(gate407inter1));
  and2  gate1949(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1950(.a(s_200), .O(gate407inter3));
  inv1  gate1951(.a(s_201), .O(gate407inter4));
  nand2 gate1952(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1953(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1954(.a(G21), .O(gate407inter7));
  inv1  gate1955(.a(G1096), .O(gate407inter8));
  nand2 gate1956(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1957(.a(s_201), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1958(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1959(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1960(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1653(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1654(.a(gate410inter0), .b(s_158), .O(gate410inter1));
  and2  gate1655(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1656(.a(s_158), .O(gate410inter3));
  inv1  gate1657(.a(s_159), .O(gate410inter4));
  nand2 gate1658(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1659(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1660(.a(G24), .O(gate410inter7));
  inv1  gate1661(.a(G1105), .O(gate410inter8));
  nand2 gate1662(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1663(.a(s_159), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1664(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1665(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1666(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate2045(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2046(.a(gate411inter0), .b(s_214), .O(gate411inter1));
  and2  gate2047(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2048(.a(s_214), .O(gate411inter3));
  inv1  gate2049(.a(s_215), .O(gate411inter4));
  nand2 gate2050(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2051(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2052(.a(G25), .O(gate411inter7));
  inv1  gate2053(.a(G1108), .O(gate411inter8));
  nand2 gate2054(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2055(.a(s_215), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2056(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2057(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2058(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2171(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2172(.a(gate412inter0), .b(s_232), .O(gate412inter1));
  and2  gate2173(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2174(.a(s_232), .O(gate412inter3));
  inv1  gate2175(.a(s_233), .O(gate412inter4));
  nand2 gate2176(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2177(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2178(.a(G26), .O(gate412inter7));
  inv1  gate2179(.a(G1111), .O(gate412inter8));
  nand2 gate2180(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2181(.a(s_233), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2182(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2183(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2184(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1233(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1234(.a(gate413inter0), .b(s_98), .O(gate413inter1));
  and2  gate1235(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1236(.a(s_98), .O(gate413inter3));
  inv1  gate1237(.a(s_99), .O(gate413inter4));
  nand2 gate1238(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1239(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1240(.a(G27), .O(gate413inter7));
  inv1  gate1241(.a(G1114), .O(gate413inter8));
  nand2 gate1242(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1243(.a(s_99), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1244(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1245(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1246(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2465(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2466(.a(gate417inter0), .b(s_274), .O(gate417inter1));
  and2  gate2467(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2468(.a(s_274), .O(gate417inter3));
  inv1  gate2469(.a(s_275), .O(gate417inter4));
  nand2 gate2470(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2471(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2472(.a(G31), .O(gate417inter7));
  inv1  gate2473(.a(G1126), .O(gate417inter8));
  nand2 gate2474(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2475(.a(s_275), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2476(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2477(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2478(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1051(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1052(.a(gate425inter0), .b(s_72), .O(gate425inter1));
  and2  gate1053(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1054(.a(s_72), .O(gate425inter3));
  inv1  gate1055(.a(s_73), .O(gate425inter4));
  nand2 gate1056(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1057(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1058(.a(G4), .O(gate425inter7));
  inv1  gate1059(.a(G1141), .O(gate425inter8));
  nand2 gate1060(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1061(.a(s_73), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1062(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1063(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1064(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1891(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1892(.a(gate434inter0), .b(s_192), .O(gate434inter1));
  and2  gate1893(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1894(.a(s_192), .O(gate434inter3));
  inv1  gate1895(.a(s_193), .O(gate434inter4));
  nand2 gate1896(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1897(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1898(.a(G1057), .O(gate434inter7));
  inv1  gate1899(.a(G1153), .O(gate434inter8));
  nand2 gate1900(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1901(.a(s_193), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1902(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1903(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1904(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate687(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate688(.a(gate435inter0), .b(s_20), .O(gate435inter1));
  and2  gate689(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate690(.a(s_20), .O(gate435inter3));
  inv1  gate691(.a(s_21), .O(gate435inter4));
  nand2 gate692(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate693(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate694(.a(G9), .O(gate435inter7));
  inv1  gate695(.a(G1156), .O(gate435inter8));
  nand2 gate696(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate697(.a(s_21), .b(gate435inter3), .O(gate435inter10));
  nor2  gate698(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate699(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate700(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1317(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1318(.a(gate437inter0), .b(s_110), .O(gate437inter1));
  and2  gate1319(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1320(.a(s_110), .O(gate437inter3));
  inv1  gate1321(.a(s_111), .O(gate437inter4));
  nand2 gate1322(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1323(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1324(.a(G10), .O(gate437inter7));
  inv1  gate1325(.a(G1159), .O(gate437inter8));
  nand2 gate1326(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1327(.a(s_111), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1328(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1329(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1330(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate813(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate814(.a(gate441inter0), .b(s_38), .O(gate441inter1));
  and2  gate815(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate816(.a(s_38), .O(gate441inter3));
  inv1  gate817(.a(s_39), .O(gate441inter4));
  nand2 gate818(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate819(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate820(.a(G12), .O(gate441inter7));
  inv1  gate821(.a(G1165), .O(gate441inter8));
  nand2 gate822(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate823(.a(s_39), .b(gate441inter3), .O(gate441inter10));
  nor2  gate824(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate825(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate826(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2395(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2396(.a(gate443inter0), .b(s_264), .O(gate443inter1));
  and2  gate2397(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2398(.a(s_264), .O(gate443inter3));
  inv1  gate2399(.a(s_265), .O(gate443inter4));
  nand2 gate2400(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2401(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2402(.a(G13), .O(gate443inter7));
  inv1  gate2403(.a(G1168), .O(gate443inter8));
  nand2 gate2404(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2405(.a(s_265), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2406(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2407(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2408(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1961(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1962(.a(gate444inter0), .b(s_202), .O(gate444inter1));
  and2  gate1963(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1964(.a(s_202), .O(gate444inter3));
  inv1  gate1965(.a(s_203), .O(gate444inter4));
  nand2 gate1966(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1967(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1968(.a(G1072), .O(gate444inter7));
  inv1  gate1969(.a(G1168), .O(gate444inter8));
  nand2 gate1970(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1971(.a(s_203), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1972(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1973(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1974(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1457(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1458(.a(gate448inter0), .b(s_130), .O(gate448inter1));
  and2  gate1459(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1460(.a(s_130), .O(gate448inter3));
  inv1  gate1461(.a(s_131), .O(gate448inter4));
  nand2 gate1462(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1463(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1464(.a(G1078), .O(gate448inter7));
  inv1  gate1465(.a(G1174), .O(gate448inter8));
  nand2 gate1466(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1467(.a(s_131), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1468(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1469(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1470(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate631(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate632(.a(gate450inter0), .b(s_12), .O(gate450inter1));
  and2  gate633(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate634(.a(s_12), .O(gate450inter3));
  inv1  gate635(.a(s_13), .O(gate450inter4));
  nand2 gate636(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate637(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate638(.a(G1081), .O(gate450inter7));
  inv1  gate639(.a(G1177), .O(gate450inter8));
  nand2 gate640(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate641(.a(s_13), .b(gate450inter3), .O(gate450inter10));
  nor2  gate642(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate643(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate644(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1429(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1430(.a(gate457inter0), .b(s_126), .O(gate457inter1));
  and2  gate1431(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1432(.a(s_126), .O(gate457inter3));
  inv1  gate1433(.a(s_127), .O(gate457inter4));
  nand2 gate1434(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1435(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1436(.a(G20), .O(gate457inter7));
  inv1  gate1437(.a(G1189), .O(gate457inter8));
  nand2 gate1438(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1439(.a(s_127), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1440(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1441(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1442(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate575(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate576(.a(gate458inter0), .b(s_4), .O(gate458inter1));
  and2  gate577(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate578(.a(s_4), .O(gate458inter3));
  inv1  gate579(.a(s_5), .O(gate458inter4));
  nand2 gate580(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate581(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate582(.a(G1093), .O(gate458inter7));
  inv1  gate583(.a(G1189), .O(gate458inter8));
  nand2 gate584(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate585(.a(s_5), .b(gate458inter3), .O(gate458inter10));
  nor2  gate586(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate587(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate588(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1275(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1276(.a(gate464inter0), .b(s_104), .O(gate464inter1));
  and2  gate1277(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1278(.a(s_104), .O(gate464inter3));
  inv1  gate1279(.a(s_105), .O(gate464inter4));
  nand2 gate1280(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1281(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1282(.a(G1102), .O(gate464inter7));
  inv1  gate1283(.a(G1198), .O(gate464inter8));
  nand2 gate1284(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1285(.a(s_105), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1286(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1287(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1288(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1443(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1444(.a(gate465inter0), .b(s_128), .O(gate465inter1));
  and2  gate1445(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1446(.a(s_128), .O(gate465inter3));
  inv1  gate1447(.a(s_129), .O(gate465inter4));
  nand2 gate1448(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1449(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1450(.a(G24), .O(gate465inter7));
  inv1  gate1451(.a(G1201), .O(gate465inter8));
  nand2 gate1452(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1453(.a(s_129), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1454(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1455(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1456(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1779(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1780(.a(gate467inter0), .b(s_176), .O(gate467inter1));
  and2  gate1781(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1782(.a(s_176), .O(gate467inter3));
  inv1  gate1783(.a(s_177), .O(gate467inter4));
  nand2 gate1784(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1785(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1786(.a(G25), .O(gate467inter7));
  inv1  gate1787(.a(G1204), .O(gate467inter8));
  nand2 gate1788(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1789(.a(s_177), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1790(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1791(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1792(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1009(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1010(.a(gate468inter0), .b(s_66), .O(gate468inter1));
  and2  gate1011(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1012(.a(s_66), .O(gate468inter3));
  inv1  gate1013(.a(s_67), .O(gate468inter4));
  nand2 gate1014(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1015(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1016(.a(G1108), .O(gate468inter7));
  inv1  gate1017(.a(G1204), .O(gate468inter8));
  nand2 gate1018(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1019(.a(s_67), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1020(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1021(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1022(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate911(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate912(.a(gate469inter0), .b(s_52), .O(gate469inter1));
  and2  gate913(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate914(.a(s_52), .O(gate469inter3));
  inv1  gate915(.a(s_53), .O(gate469inter4));
  nand2 gate916(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate917(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate918(.a(G26), .O(gate469inter7));
  inv1  gate919(.a(G1207), .O(gate469inter8));
  nand2 gate920(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate921(.a(s_53), .b(gate469inter3), .O(gate469inter10));
  nor2  gate922(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate923(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate924(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate757(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate758(.a(gate470inter0), .b(s_30), .O(gate470inter1));
  and2  gate759(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate760(.a(s_30), .O(gate470inter3));
  inv1  gate761(.a(s_31), .O(gate470inter4));
  nand2 gate762(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate763(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate764(.a(G1111), .O(gate470inter7));
  inv1  gate765(.a(G1207), .O(gate470inter8));
  nand2 gate766(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate767(.a(s_31), .b(gate470inter3), .O(gate470inter10));
  nor2  gate768(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate769(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate770(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2367(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2368(.a(gate477inter0), .b(s_260), .O(gate477inter1));
  and2  gate2369(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2370(.a(s_260), .O(gate477inter3));
  inv1  gate2371(.a(s_261), .O(gate477inter4));
  nand2 gate2372(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2373(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2374(.a(G30), .O(gate477inter7));
  inv1  gate2375(.a(G1219), .O(gate477inter8));
  nand2 gate2376(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2377(.a(s_261), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2378(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2379(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2380(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate673(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate674(.a(gate480inter0), .b(s_18), .O(gate480inter1));
  and2  gate675(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate676(.a(s_18), .O(gate480inter3));
  inv1  gate677(.a(s_19), .O(gate480inter4));
  nand2 gate678(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate679(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate680(.a(G1126), .O(gate480inter7));
  inv1  gate681(.a(G1222), .O(gate480inter8));
  nand2 gate682(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate683(.a(s_19), .b(gate480inter3), .O(gate480inter10));
  nor2  gate684(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate685(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate686(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1093(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1094(.a(gate482inter0), .b(s_78), .O(gate482inter1));
  and2  gate1095(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1096(.a(s_78), .O(gate482inter3));
  inv1  gate1097(.a(s_79), .O(gate482inter4));
  nand2 gate1098(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1099(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1100(.a(G1129), .O(gate482inter7));
  inv1  gate1101(.a(G1225), .O(gate482inter8));
  nand2 gate1102(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1103(.a(s_79), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1104(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1105(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1106(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate2003(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2004(.a(gate483inter0), .b(s_208), .O(gate483inter1));
  and2  gate2005(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2006(.a(s_208), .O(gate483inter3));
  inv1  gate2007(.a(s_209), .O(gate483inter4));
  nand2 gate2008(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2009(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2010(.a(G1228), .O(gate483inter7));
  inv1  gate2011(.a(G1229), .O(gate483inter8));
  nand2 gate2012(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2013(.a(s_209), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2014(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2015(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2016(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1177(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1178(.a(gate484inter0), .b(s_90), .O(gate484inter1));
  and2  gate1179(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1180(.a(s_90), .O(gate484inter3));
  inv1  gate1181(.a(s_91), .O(gate484inter4));
  nand2 gate1182(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1183(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1184(.a(G1230), .O(gate484inter7));
  inv1  gate1185(.a(G1231), .O(gate484inter8));
  nand2 gate1186(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1187(.a(s_91), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1188(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1189(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1190(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1975(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1976(.a(gate487inter0), .b(s_204), .O(gate487inter1));
  and2  gate1977(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1978(.a(s_204), .O(gate487inter3));
  inv1  gate1979(.a(s_205), .O(gate487inter4));
  nand2 gate1980(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1981(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1982(.a(G1236), .O(gate487inter7));
  inv1  gate1983(.a(G1237), .O(gate487inter8));
  nand2 gate1984(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1985(.a(s_205), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1986(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1987(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1988(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2031(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2032(.a(gate488inter0), .b(s_212), .O(gate488inter1));
  and2  gate2033(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2034(.a(s_212), .O(gate488inter3));
  inv1  gate2035(.a(s_213), .O(gate488inter4));
  nand2 gate2036(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2037(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2038(.a(G1238), .O(gate488inter7));
  inv1  gate2039(.a(G1239), .O(gate488inter8));
  nand2 gate2040(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2041(.a(s_213), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2042(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2043(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2044(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2283(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2284(.a(gate490inter0), .b(s_248), .O(gate490inter1));
  and2  gate2285(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2286(.a(s_248), .O(gate490inter3));
  inv1  gate2287(.a(s_249), .O(gate490inter4));
  nand2 gate2288(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2289(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2290(.a(G1242), .O(gate490inter7));
  inv1  gate2291(.a(G1243), .O(gate490inter8));
  nand2 gate2292(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2293(.a(s_249), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2294(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2295(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2296(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2185(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2186(.a(gate496inter0), .b(s_234), .O(gate496inter1));
  and2  gate2187(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2188(.a(s_234), .O(gate496inter3));
  inv1  gate2189(.a(s_235), .O(gate496inter4));
  nand2 gate2190(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2191(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2192(.a(G1254), .O(gate496inter7));
  inv1  gate2193(.a(G1255), .O(gate496inter8));
  nand2 gate2194(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2195(.a(s_235), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2196(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2197(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2198(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1863(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1864(.a(gate500inter0), .b(s_188), .O(gate500inter1));
  and2  gate1865(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1866(.a(s_188), .O(gate500inter3));
  inv1  gate1867(.a(s_189), .O(gate500inter4));
  nand2 gate1868(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1869(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1870(.a(G1262), .O(gate500inter7));
  inv1  gate1871(.a(G1263), .O(gate500inter8));
  nand2 gate1872(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1873(.a(s_189), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1874(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1875(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1876(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1639(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1640(.a(gate501inter0), .b(s_156), .O(gate501inter1));
  and2  gate1641(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1642(.a(s_156), .O(gate501inter3));
  inv1  gate1643(.a(s_157), .O(gate501inter4));
  nand2 gate1644(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1645(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1646(.a(G1264), .O(gate501inter7));
  inv1  gate1647(.a(G1265), .O(gate501inter8));
  nand2 gate1648(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1649(.a(s_157), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1650(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1651(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1652(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1163(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1164(.a(gate503inter0), .b(s_88), .O(gate503inter1));
  and2  gate1165(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1166(.a(s_88), .O(gate503inter3));
  inv1  gate1167(.a(s_89), .O(gate503inter4));
  nand2 gate1168(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1169(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1170(.a(G1268), .O(gate503inter7));
  inv1  gate1171(.a(G1269), .O(gate503inter8));
  nand2 gate1172(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1173(.a(s_89), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1174(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1175(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1176(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2129(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2130(.a(gate506inter0), .b(s_226), .O(gate506inter1));
  and2  gate2131(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2132(.a(s_226), .O(gate506inter3));
  inv1  gate2133(.a(s_227), .O(gate506inter4));
  nand2 gate2134(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2135(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2136(.a(G1274), .O(gate506inter7));
  inv1  gate2137(.a(G1275), .O(gate506inter8));
  nand2 gate2138(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2139(.a(s_227), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2140(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2141(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2142(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2535(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2536(.a(gate508inter0), .b(s_284), .O(gate508inter1));
  and2  gate2537(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2538(.a(s_284), .O(gate508inter3));
  inv1  gate2539(.a(s_285), .O(gate508inter4));
  nand2 gate2540(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2541(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2542(.a(G1278), .O(gate508inter7));
  inv1  gate2543(.a(G1279), .O(gate508inter8));
  nand2 gate2544(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2545(.a(s_285), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2546(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2547(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2548(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1849(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1850(.a(gate514inter0), .b(s_186), .O(gate514inter1));
  and2  gate1851(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1852(.a(s_186), .O(gate514inter3));
  inv1  gate1853(.a(s_187), .O(gate514inter4));
  nand2 gate1854(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1855(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1856(.a(G1290), .O(gate514inter7));
  inv1  gate1857(.a(G1291), .O(gate514inter8));
  nand2 gate1858(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1859(.a(s_187), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1860(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1861(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1862(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule