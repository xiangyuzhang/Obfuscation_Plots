module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate673(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate674(.a(gate9inter0), .b(s_18), .O(gate9inter1));
  and2  gate675(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate676(.a(s_18), .O(gate9inter3));
  inv1  gate677(.a(s_19), .O(gate9inter4));
  nand2 gate678(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate679(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate680(.a(G1), .O(gate9inter7));
  inv1  gate681(.a(G2), .O(gate9inter8));
  nand2 gate682(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate683(.a(s_19), .b(gate9inter3), .O(gate9inter10));
  nor2  gate684(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate685(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate686(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1667(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1668(.a(gate13inter0), .b(s_160), .O(gate13inter1));
  and2  gate1669(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1670(.a(s_160), .O(gate13inter3));
  inv1  gate1671(.a(s_161), .O(gate13inter4));
  nand2 gate1672(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1673(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1674(.a(G9), .O(gate13inter7));
  inv1  gate1675(.a(G10), .O(gate13inter8));
  nand2 gate1676(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1677(.a(s_161), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1678(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1679(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1680(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1555(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1556(.a(gate19inter0), .b(s_144), .O(gate19inter1));
  and2  gate1557(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1558(.a(s_144), .O(gate19inter3));
  inv1  gate1559(.a(s_145), .O(gate19inter4));
  nand2 gate1560(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1561(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1562(.a(G21), .O(gate19inter7));
  inv1  gate1563(.a(G22), .O(gate19inter8));
  nand2 gate1564(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1565(.a(s_145), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1566(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1567(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1568(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate897(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate898(.a(gate24inter0), .b(s_50), .O(gate24inter1));
  and2  gate899(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate900(.a(s_50), .O(gate24inter3));
  inv1  gate901(.a(s_51), .O(gate24inter4));
  nand2 gate902(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate903(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate904(.a(G31), .O(gate24inter7));
  inv1  gate905(.a(G32), .O(gate24inter8));
  nand2 gate906(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate907(.a(s_51), .b(gate24inter3), .O(gate24inter10));
  nor2  gate908(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate909(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate910(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1261(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1262(.a(gate29inter0), .b(s_102), .O(gate29inter1));
  and2  gate1263(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1264(.a(s_102), .O(gate29inter3));
  inv1  gate1265(.a(s_103), .O(gate29inter4));
  nand2 gate1266(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1267(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1268(.a(G3), .O(gate29inter7));
  inv1  gate1269(.a(G7), .O(gate29inter8));
  nand2 gate1270(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1271(.a(s_103), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1272(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1273(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1274(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1093(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1094(.a(gate37inter0), .b(s_78), .O(gate37inter1));
  and2  gate1095(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1096(.a(s_78), .O(gate37inter3));
  inv1  gate1097(.a(s_79), .O(gate37inter4));
  nand2 gate1098(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1099(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1100(.a(G19), .O(gate37inter7));
  inv1  gate1101(.a(G23), .O(gate37inter8));
  nand2 gate1102(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1103(.a(s_79), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1104(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1105(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1106(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1485(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1486(.a(gate40inter0), .b(s_134), .O(gate40inter1));
  and2  gate1487(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1488(.a(s_134), .O(gate40inter3));
  inv1  gate1489(.a(s_135), .O(gate40inter4));
  nand2 gate1490(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1491(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1492(.a(G28), .O(gate40inter7));
  inv1  gate1493(.a(G32), .O(gate40inter8));
  nand2 gate1494(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1495(.a(s_135), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1496(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1497(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1498(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1793(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1794(.a(gate41inter0), .b(s_178), .O(gate41inter1));
  and2  gate1795(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1796(.a(s_178), .O(gate41inter3));
  inv1  gate1797(.a(s_179), .O(gate41inter4));
  nand2 gate1798(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1799(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1800(.a(G1), .O(gate41inter7));
  inv1  gate1801(.a(G266), .O(gate41inter8));
  nand2 gate1802(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1803(.a(s_179), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1804(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1805(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1806(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1065(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1066(.a(gate46inter0), .b(s_74), .O(gate46inter1));
  and2  gate1067(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1068(.a(s_74), .O(gate46inter3));
  inv1  gate1069(.a(s_75), .O(gate46inter4));
  nand2 gate1070(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1071(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1072(.a(G6), .O(gate46inter7));
  inv1  gate1073(.a(G272), .O(gate46inter8));
  nand2 gate1074(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1075(.a(s_75), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1076(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1077(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1078(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1681(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1682(.a(gate51inter0), .b(s_162), .O(gate51inter1));
  and2  gate1683(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1684(.a(s_162), .O(gate51inter3));
  inv1  gate1685(.a(s_163), .O(gate51inter4));
  nand2 gate1686(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1687(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1688(.a(G11), .O(gate51inter7));
  inv1  gate1689(.a(G281), .O(gate51inter8));
  nand2 gate1690(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1691(.a(s_163), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1692(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1693(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1694(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate603(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate604(.a(gate56inter0), .b(s_8), .O(gate56inter1));
  and2  gate605(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate606(.a(s_8), .O(gate56inter3));
  inv1  gate607(.a(s_9), .O(gate56inter4));
  nand2 gate608(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate609(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate610(.a(G16), .O(gate56inter7));
  inv1  gate611(.a(G287), .O(gate56inter8));
  nand2 gate612(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate613(.a(s_9), .b(gate56inter3), .O(gate56inter10));
  nor2  gate614(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate615(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate616(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1331(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1332(.a(gate60inter0), .b(s_112), .O(gate60inter1));
  and2  gate1333(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1334(.a(s_112), .O(gate60inter3));
  inv1  gate1335(.a(s_113), .O(gate60inter4));
  nand2 gate1336(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1337(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1338(.a(G20), .O(gate60inter7));
  inv1  gate1339(.a(G293), .O(gate60inter8));
  nand2 gate1340(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1341(.a(s_113), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1342(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1343(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1344(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate911(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate912(.a(gate64inter0), .b(s_52), .O(gate64inter1));
  and2  gate913(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate914(.a(s_52), .O(gate64inter3));
  inv1  gate915(.a(s_53), .O(gate64inter4));
  nand2 gate916(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate917(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate918(.a(G24), .O(gate64inter7));
  inv1  gate919(.a(G299), .O(gate64inter8));
  nand2 gate920(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate921(.a(s_53), .b(gate64inter3), .O(gate64inter10));
  nor2  gate922(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate923(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate924(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1597(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1598(.a(gate81inter0), .b(s_150), .O(gate81inter1));
  and2  gate1599(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1600(.a(s_150), .O(gate81inter3));
  inv1  gate1601(.a(s_151), .O(gate81inter4));
  nand2 gate1602(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1603(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1604(.a(G3), .O(gate81inter7));
  inv1  gate1605(.a(G326), .O(gate81inter8));
  nand2 gate1606(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1607(.a(s_151), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1608(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1609(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1610(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1359(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1360(.a(gate86inter0), .b(s_116), .O(gate86inter1));
  and2  gate1361(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1362(.a(s_116), .O(gate86inter3));
  inv1  gate1363(.a(s_117), .O(gate86inter4));
  nand2 gate1364(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1365(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1366(.a(G8), .O(gate86inter7));
  inv1  gate1367(.a(G332), .O(gate86inter8));
  nand2 gate1368(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1369(.a(s_117), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1370(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1371(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1372(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate561(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate562(.a(gate90inter0), .b(s_2), .O(gate90inter1));
  and2  gate563(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate564(.a(s_2), .O(gate90inter3));
  inv1  gate565(.a(s_3), .O(gate90inter4));
  nand2 gate566(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate567(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate568(.a(G21), .O(gate90inter7));
  inv1  gate569(.a(G338), .O(gate90inter8));
  nand2 gate570(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate571(.a(s_3), .b(gate90inter3), .O(gate90inter10));
  nor2  gate572(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate573(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate574(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate883(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate884(.a(gate91inter0), .b(s_48), .O(gate91inter1));
  and2  gate885(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate886(.a(s_48), .O(gate91inter3));
  inv1  gate887(.a(s_49), .O(gate91inter4));
  nand2 gate888(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate889(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate890(.a(G25), .O(gate91inter7));
  inv1  gate891(.a(G341), .O(gate91inter8));
  nand2 gate892(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate893(.a(s_49), .b(gate91inter3), .O(gate91inter10));
  nor2  gate894(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate895(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate896(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1149(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1150(.a(gate93inter0), .b(s_86), .O(gate93inter1));
  and2  gate1151(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1152(.a(s_86), .O(gate93inter3));
  inv1  gate1153(.a(s_87), .O(gate93inter4));
  nand2 gate1154(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1155(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1156(.a(G18), .O(gate93inter7));
  inv1  gate1157(.a(G344), .O(gate93inter8));
  nand2 gate1158(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1159(.a(s_87), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1160(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1161(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1162(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1765(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1766(.a(gate94inter0), .b(s_174), .O(gate94inter1));
  and2  gate1767(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1768(.a(s_174), .O(gate94inter3));
  inv1  gate1769(.a(s_175), .O(gate94inter4));
  nand2 gate1770(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1771(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1772(.a(G22), .O(gate94inter7));
  inv1  gate1773(.a(G344), .O(gate94inter8));
  nand2 gate1774(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1775(.a(s_175), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1776(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1777(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1778(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate827(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate828(.a(gate106inter0), .b(s_40), .O(gate106inter1));
  and2  gate829(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate830(.a(s_40), .O(gate106inter3));
  inv1  gate831(.a(s_41), .O(gate106inter4));
  nand2 gate832(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate833(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate834(.a(G364), .O(gate106inter7));
  inv1  gate835(.a(G365), .O(gate106inter8));
  nand2 gate836(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate837(.a(s_41), .b(gate106inter3), .O(gate106inter10));
  nor2  gate838(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate839(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate840(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1205(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1206(.a(gate108inter0), .b(s_94), .O(gate108inter1));
  and2  gate1207(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1208(.a(s_94), .O(gate108inter3));
  inv1  gate1209(.a(s_95), .O(gate108inter4));
  nand2 gate1210(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1211(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1212(.a(G368), .O(gate108inter7));
  inv1  gate1213(.a(G369), .O(gate108inter8));
  nand2 gate1214(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1215(.a(s_95), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1216(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1217(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1218(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1457(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1458(.a(gate110inter0), .b(s_130), .O(gate110inter1));
  and2  gate1459(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1460(.a(s_130), .O(gate110inter3));
  inv1  gate1461(.a(s_131), .O(gate110inter4));
  nand2 gate1462(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1463(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1464(.a(G372), .O(gate110inter7));
  inv1  gate1465(.a(G373), .O(gate110inter8));
  nand2 gate1466(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1467(.a(s_131), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1468(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1469(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1470(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate575(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate576(.a(gate113inter0), .b(s_4), .O(gate113inter1));
  and2  gate577(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate578(.a(s_4), .O(gate113inter3));
  inv1  gate579(.a(s_5), .O(gate113inter4));
  nand2 gate580(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate581(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate582(.a(G378), .O(gate113inter7));
  inv1  gate583(.a(G379), .O(gate113inter8));
  nand2 gate584(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate585(.a(s_5), .b(gate113inter3), .O(gate113inter10));
  nor2  gate586(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate587(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate588(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate785(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate786(.a(gate114inter0), .b(s_34), .O(gate114inter1));
  and2  gate787(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate788(.a(s_34), .O(gate114inter3));
  inv1  gate789(.a(s_35), .O(gate114inter4));
  nand2 gate790(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate791(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate792(.a(G380), .O(gate114inter7));
  inv1  gate793(.a(G381), .O(gate114inter8));
  nand2 gate794(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate795(.a(s_35), .b(gate114inter3), .O(gate114inter10));
  nor2  gate796(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate797(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate798(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1443(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1444(.a(gate124inter0), .b(s_128), .O(gate124inter1));
  and2  gate1445(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1446(.a(s_128), .O(gate124inter3));
  inv1  gate1447(.a(s_129), .O(gate124inter4));
  nand2 gate1448(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1449(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1450(.a(G400), .O(gate124inter7));
  inv1  gate1451(.a(G401), .O(gate124inter8));
  nand2 gate1452(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1453(.a(s_129), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1454(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1455(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1456(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate589(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate590(.a(gate128inter0), .b(s_6), .O(gate128inter1));
  and2  gate591(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate592(.a(s_6), .O(gate128inter3));
  inv1  gate593(.a(s_7), .O(gate128inter4));
  nand2 gate594(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate595(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate596(.a(G408), .O(gate128inter7));
  inv1  gate597(.a(G409), .O(gate128inter8));
  nand2 gate598(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate599(.a(s_7), .b(gate128inter3), .O(gate128inter10));
  nor2  gate600(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate601(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate602(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate855(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate856(.a(gate129inter0), .b(s_44), .O(gate129inter1));
  and2  gate857(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate858(.a(s_44), .O(gate129inter3));
  inv1  gate859(.a(s_45), .O(gate129inter4));
  nand2 gate860(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate861(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate862(.a(G410), .O(gate129inter7));
  inv1  gate863(.a(G411), .O(gate129inter8));
  nand2 gate864(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate865(.a(s_45), .b(gate129inter3), .O(gate129inter10));
  nor2  gate866(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate867(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate868(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1233(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1234(.a(gate137inter0), .b(s_98), .O(gate137inter1));
  and2  gate1235(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1236(.a(s_98), .O(gate137inter3));
  inv1  gate1237(.a(s_99), .O(gate137inter4));
  nand2 gate1238(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1239(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1240(.a(G426), .O(gate137inter7));
  inv1  gate1241(.a(G429), .O(gate137inter8));
  nand2 gate1242(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1243(.a(s_99), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1244(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1245(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1246(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1779(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1780(.a(gate140inter0), .b(s_176), .O(gate140inter1));
  and2  gate1781(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1782(.a(s_176), .O(gate140inter3));
  inv1  gate1783(.a(s_177), .O(gate140inter4));
  nand2 gate1784(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1785(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1786(.a(G444), .O(gate140inter7));
  inv1  gate1787(.a(G447), .O(gate140inter8));
  nand2 gate1788(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1789(.a(s_177), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1790(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1791(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1792(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1275(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1276(.a(gate141inter0), .b(s_104), .O(gate141inter1));
  and2  gate1277(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1278(.a(s_104), .O(gate141inter3));
  inv1  gate1279(.a(s_105), .O(gate141inter4));
  nand2 gate1280(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1281(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1282(.a(G450), .O(gate141inter7));
  inv1  gate1283(.a(G453), .O(gate141inter8));
  nand2 gate1284(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1285(.a(s_105), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1286(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1287(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1288(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1695(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1696(.a(gate166inter0), .b(s_164), .O(gate166inter1));
  and2  gate1697(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1698(.a(s_164), .O(gate166inter3));
  inv1  gate1699(.a(s_165), .O(gate166inter4));
  nand2 gate1700(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1701(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1702(.a(G465), .O(gate166inter7));
  inv1  gate1703(.a(G540), .O(gate166inter8));
  nand2 gate1704(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1705(.a(s_165), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1706(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1707(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1708(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate939(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate940(.a(gate170inter0), .b(s_56), .O(gate170inter1));
  and2  gate941(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate942(.a(s_56), .O(gate170inter3));
  inv1  gate943(.a(s_57), .O(gate170inter4));
  nand2 gate944(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate945(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate946(.a(G477), .O(gate170inter7));
  inv1  gate947(.a(G546), .O(gate170inter8));
  nand2 gate948(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate949(.a(s_57), .b(gate170inter3), .O(gate170inter10));
  nor2  gate950(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate951(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate952(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1639(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1640(.a(gate180inter0), .b(s_156), .O(gate180inter1));
  and2  gate1641(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1642(.a(s_156), .O(gate180inter3));
  inv1  gate1643(.a(s_157), .O(gate180inter4));
  nand2 gate1644(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1645(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1646(.a(G507), .O(gate180inter7));
  inv1  gate1647(.a(G561), .O(gate180inter8));
  nand2 gate1648(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1649(.a(s_157), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1650(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1651(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1652(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1247(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1248(.a(gate181inter0), .b(s_100), .O(gate181inter1));
  and2  gate1249(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1250(.a(s_100), .O(gate181inter3));
  inv1  gate1251(.a(s_101), .O(gate181inter4));
  nand2 gate1252(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1253(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1254(.a(G510), .O(gate181inter7));
  inv1  gate1255(.a(G564), .O(gate181inter8));
  nand2 gate1256(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1257(.a(s_101), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1258(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1259(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1260(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1569(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1570(.a(gate186inter0), .b(s_146), .O(gate186inter1));
  and2  gate1571(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1572(.a(s_146), .O(gate186inter3));
  inv1  gate1573(.a(s_147), .O(gate186inter4));
  nand2 gate1574(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1575(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1576(.a(G572), .O(gate186inter7));
  inv1  gate1577(.a(G573), .O(gate186inter8));
  nand2 gate1578(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1579(.a(s_147), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1580(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1581(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1582(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate869(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate870(.a(gate187inter0), .b(s_46), .O(gate187inter1));
  and2  gate871(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate872(.a(s_46), .O(gate187inter3));
  inv1  gate873(.a(s_47), .O(gate187inter4));
  nand2 gate874(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate875(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate876(.a(G574), .O(gate187inter7));
  inv1  gate877(.a(G575), .O(gate187inter8));
  nand2 gate878(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate879(.a(s_47), .b(gate187inter3), .O(gate187inter10));
  nor2  gate880(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate881(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate882(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1387(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1388(.a(gate191inter0), .b(s_120), .O(gate191inter1));
  and2  gate1389(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1390(.a(s_120), .O(gate191inter3));
  inv1  gate1391(.a(s_121), .O(gate191inter4));
  nand2 gate1392(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1393(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1394(.a(G582), .O(gate191inter7));
  inv1  gate1395(.a(G583), .O(gate191inter8));
  nand2 gate1396(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1397(.a(s_121), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1398(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1399(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1400(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1471(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1472(.a(gate194inter0), .b(s_132), .O(gate194inter1));
  and2  gate1473(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1474(.a(s_132), .O(gate194inter3));
  inv1  gate1475(.a(s_133), .O(gate194inter4));
  nand2 gate1476(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1477(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1478(.a(G588), .O(gate194inter7));
  inv1  gate1479(.a(G589), .O(gate194inter8));
  nand2 gate1480(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1481(.a(s_133), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1482(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1483(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1484(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate645(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate646(.a(gate197inter0), .b(s_14), .O(gate197inter1));
  and2  gate647(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate648(.a(s_14), .O(gate197inter3));
  inv1  gate649(.a(s_15), .O(gate197inter4));
  nand2 gate650(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate651(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate652(.a(G594), .O(gate197inter7));
  inv1  gate653(.a(G595), .O(gate197inter8));
  nand2 gate654(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate655(.a(s_15), .b(gate197inter3), .O(gate197inter10));
  nor2  gate656(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate657(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate658(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate547(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate548(.a(gate200inter0), .b(s_0), .O(gate200inter1));
  and2  gate549(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate550(.a(s_0), .O(gate200inter3));
  inv1  gate551(.a(s_1), .O(gate200inter4));
  nand2 gate552(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate553(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate554(.a(G600), .O(gate200inter7));
  inv1  gate555(.a(G601), .O(gate200inter8));
  nand2 gate556(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate557(.a(s_1), .b(gate200inter3), .O(gate200inter10));
  nor2  gate558(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate559(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate560(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1163(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1164(.a(gate206inter0), .b(s_88), .O(gate206inter1));
  and2  gate1165(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1166(.a(s_88), .O(gate206inter3));
  inv1  gate1167(.a(s_89), .O(gate206inter4));
  nand2 gate1168(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1169(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1170(.a(G632), .O(gate206inter7));
  inv1  gate1171(.a(G637), .O(gate206inter8));
  nand2 gate1172(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1173(.a(s_89), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1174(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1175(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1176(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate841(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate842(.a(gate208inter0), .b(s_42), .O(gate208inter1));
  and2  gate843(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate844(.a(s_42), .O(gate208inter3));
  inv1  gate845(.a(s_43), .O(gate208inter4));
  nand2 gate846(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate847(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate848(.a(G627), .O(gate208inter7));
  inv1  gate849(.a(G637), .O(gate208inter8));
  nand2 gate850(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate851(.a(s_43), .b(gate208inter3), .O(gate208inter10));
  nor2  gate852(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate853(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate854(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1135(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1136(.a(gate210inter0), .b(s_84), .O(gate210inter1));
  and2  gate1137(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1138(.a(s_84), .O(gate210inter3));
  inv1  gate1139(.a(s_85), .O(gate210inter4));
  nand2 gate1140(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1141(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1142(.a(G607), .O(gate210inter7));
  inv1  gate1143(.a(G666), .O(gate210inter8));
  nand2 gate1144(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1145(.a(s_85), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1146(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1147(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1148(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate687(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate688(.a(gate212inter0), .b(s_20), .O(gate212inter1));
  and2  gate689(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate690(.a(s_20), .O(gate212inter3));
  inv1  gate691(.a(s_21), .O(gate212inter4));
  nand2 gate692(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate693(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate694(.a(G617), .O(gate212inter7));
  inv1  gate695(.a(G669), .O(gate212inter8));
  nand2 gate696(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate697(.a(s_21), .b(gate212inter3), .O(gate212inter10));
  nor2  gate698(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate699(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate700(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate967(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate968(.a(gate213inter0), .b(s_60), .O(gate213inter1));
  and2  gate969(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate970(.a(s_60), .O(gate213inter3));
  inv1  gate971(.a(s_61), .O(gate213inter4));
  nand2 gate972(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate973(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate974(.a(G602), .O(gate213inter7));
  inv1  gate975(.a(G672), .O(gate213inter8));
  nand2 gate976(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate977(.a(s_61), .b(gate213inter3), .O(gate213inter10));
  nor2  gate978(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate979(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate980(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1723(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1724(.a(gate217inter0), .b(s_168), .O(gate217inter1));
  and2  gate1725(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1726(.a(s_168), .O(gate217inter3));
  inv1  gate1727(.a(s_169), .O(gate217inter4));
  nand2 gate1728(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1729(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1730(.a(G622), .O(gate217inter7));
  inv1  gate1731(.a(G678), .O(gate217inter8));
  nand2 gate1732(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1733(.a(s_169), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1734(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1735(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1736(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate953(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate954(.a(gate222inter0), .b(s_58), .O(gate222inter1));
  and2  gate955(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate956(.a(s_58), .O(gate222inter3));
  inv1  gate957(.a(s_59), .O(gate222inter4));
  nand2 gate958(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate959(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate960(.a(G632), .O(gate222inter7));
  inv1  gate961(.a(G684), .O(gate222inter8));
  nand2 gate962(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate963(.a(s_59), .b(gate222inter3), .O(gate222inter10));
  nor2  gate964(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate965(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate966(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate701(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate702(.a(gate230inter0), .b(s_22), .O(gate230inter1));
  and2  gate703(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate704(.a(s_22), .O(gate230inter3));
  inv1  gate705(.a(s_23), .O(gate230inter4));
  nand2 gate706(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate707(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate708(.a(G700), .O(gate230inter7));
  inv1  gate709(.a(G701), .O(gate230inter8));
  nand2 gate710(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate711(.a(s_23), .b(gate230inter3), .O(gate230inter10));
  nor2  gate712(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate713(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate714(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate715(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate716(.a(gate248inter0), .b(s_24), .O(gate248inter1));
  and2  gate717(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate718(.a(s_24), .O(gate248inter3));
  inv1  gate719(.a(s_25), .O(gate248inter4));
  nand2 gate720(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate721(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate722(.a(G727), .O(gate248inter7));
  inv1  gate723(.a(G739), .O(gate248inter8));
  nand2 gate724(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate725(.a(s_25), .b(gate248inter3), .O(gate248inter10));
  nor2  gate726(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate727(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate728(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1373(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1374(.a(gate257inter0), .b(s_118), .O(gate257inter1));
  and2  gate1375(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1376(.a(s_118), .O(gate257inter3));
  inv1  gate1377(.a(s_119), .O(gate257inter4));
  nand2 gate1378(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1379(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1380(.a(G754), .O(gate257inter7));
  inv1  gate1381(.a(G755), .O(gate257inter8));
  nand2 gate1382(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1383(.a(s_119), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1384(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1385(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1386(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1219(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1220(.a(gate259inter0), .b(s_96), .O(gate259inter1));
  and2  gate1221(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1222(.a(s_96), .O(gate259inter3));
  inv1  gate1223(.a(s_97), .O(gate259inter4));
  nand2 gate1224(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1225(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1226(.a(G758), .O(gate259inter7));
  inv1  gate1227(.a(G759), .O(gate259inter8));
  nand2 gate1228(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1229(.a(s_97), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1230(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1231(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1232(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1583(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1584(.a(gate263inter0), .b(s_148), .O(gate263inter1));
  and2  gate1585(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1586(.a(s_148), .O(gate263inter3));
  inv1  gate1587(.a(s_149), .O(gate263inter4));
  nand2 gate1588(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1589(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1590(.a(G766), .O(gate263inter7));
  inv1  gate1591(.a(G767), .O(gate263inter8));
  nand2 gate1592(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1593(.a(s_149), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1594(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1595(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1596(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1611(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1612(.a(gate270inter0), .b(s_152), .O(gate270inter1));
  and2  gate1613(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1614(.a(s_152), .O(gate270inter3));
  inv1  gate1615(.a(s_153), .O(gate270inter4));
  nand2 gate1616(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1617(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1618(.a(G657), .O(gate270inter7));
  inv1  gate1619(.a(G785), .O(gate270inter8));
  nand2 gate1620(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1621(.a(s_153), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1622(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1623(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1624(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate995(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate996(.a(gate271inter0), .b(s_64), .O(gate271inter1));
  and2  gate997(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate998(.a(s_64), .O(gate271inter3));
  inv1  gate999(.a(s_65), .O(gate271inter4));
  nand2 gate1000(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1001(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1002(.a(G660), .O(gate271inter7));
  inv1  gate1003(.a(G788), .O(gate271inter8));
  nand2 gate1004(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1005(.a(s_65), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1006(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1007(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1008(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate757(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate758(.a(gate273inter0), .b(s_30), .O(gate273inter1));
  and2  gate759(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate760(.a(s_30), .O(gate273inter3));
  inv1  gate761(.a(s_31), .O(gate273inter4));
  nand2 gate762(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate763(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate764(.a(G642), .O(gate273inter7));
  inv1  gate765(.a(G794), .O(gate273inter8));
  nand2 gate766(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate767(.a(s_31), .b(gate273inter3), .O(gate273inter10));
  nor2  gate768(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate769(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate770(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate659(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate660(.a(gate274inter0), .b(s_16), .O(gate274inter1));
  and2  gate661(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate662(.a(s_16), .O(gate274inter3));
  inv1  gate663(.a(s_17), .O(gate274inter4));
  nand2 gate664(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate665(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate666(.a(G770), .O(gate274inter7));
  inv1  gate667(.a(G794), .O(gate274inter8));
  nand2 gate668(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate669(.a(s_17), .b(gate274inter3), .O(gate274inter10));
  nor2  gate670(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate671(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate672(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1737(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1738(.a(gate282inter0), .b(s_170), .O(gate282inter1));
  and2  gate1739(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1740(.a(s_170), .O(gate282inter3));
  inv1  gate1741(.a(s_171), .O(gate282inter4));
  nand2 gate1742(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1743(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1744(.a(G782), .O(gate282inter7));
  inv1  gate1745(.a(G806), .O(gate282inter8));
  nand2 gate1746(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1747(.a(s_171), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1748(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1749(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1750(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1415(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1416(.a(gate283inter0), .b(s_124), .O(gate283inter1));
  and2  gate1417(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1418(.a(s_124), .O(gate283inter3));
  inv1  gate1419(.a(s_125), .O(gate283inter4));
  nand2 gate1420(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1421(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1422(.a(G657), .O(gate283inter7));
  inv1  gate1423(.a(G809), .O(gate283inter8));
  nand2 gate1424(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1425(.a(s_125), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1426(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1427(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1428(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate981(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate982(.a(gate285inter0), .b(s_62), .O(gate285inter1));
  and2  gate983(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate984(.a(s_62), .O(gate285inter3));
  inv1  gate985(.a(s_63), .O(gate285inter4));
  nand2 gate986(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate987(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate988(.a(G660), .O(gate285inter7));
  inv1  gate989(.a(G812), .O(gate285inter8));
  nand2 gate990(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate991(.a(s_63), .b(gate285inter3), .O(gate285inter10));
  nor2  gate992(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate993(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate994(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1401(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1402(.a(gate289inter0), .b(s_122), .O(gate289inter1));
  and2  gate1403(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1404(.a(s_122), .O(gate289inter3));
  inv1  gate1405(.a(s_123), .O(gate289inter4));
  nand2 gate1406(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1407(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1408(.a(G818), .O(gate289inter7));
  inv1  gate1409(.a(G819), .O(gate289inter8));
  nand2 gate1410(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1411(.a(s_123), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1412(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1413(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1414(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1345(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1346(.a(gate291inter0), .b(s_114), .O(gate291inter1));
  and2  gate1347(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1348(.a(s_114), .O(gate291inter3));
  inv1  gate1349(.a(s_115), .O(gate291inter4));
  nand2 gate1350(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1351(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1352(.a(G822), .O(gate291inter7));
  inv1  gate1353(.a(G823), .O(gate291inter8));
  nand2 gate1354(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1355(.a(s_115), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1356(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1357(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1358(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1009(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1010(.a(gate294inter0), .b(s_66), .O(gate294inter1));
  and2  gate1011(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1012(.a(s_66), .O(gate294inter3));
  inv1  gate1013(.a(s_67), .O(gate294inter4));
  nand2 gate1014(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1015(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1016(.a(G832), .O(gate294inter7));
  inv1  gate1017(.a(G833), .O(gate294inter8));
  nand2 gate1018(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1019(.a(s_67), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1020(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1021(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1022(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate743(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate744(.a(gate295inter0), .b(s_28), .O(gate295inter1));
  and2  gate745(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate746(.a(s_28), .O(gate295inter3));
  inv1  gate747(.a(s_29), .O(gate295inter4));
  nand2 gate748(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate749(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate750(.a(G830), .O(gate295inter7));
  inv1  gate751(.a(G831), .O(gate295inter8));
  nand2 gate752(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate753(.a(s_29), .b(gate295inter3), .O(gate295inter10));
  nor2  gate754(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate755(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate756(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate771(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate772(.a(gate389inter0), .b(s_32), .O(gate389inter1));
  and2  gate773(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate774(.a(s_32), .O(gate389inter3));
  inv1  gate775(.a(s_33), .O(gate389inter4));
  nand2 gate776(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate777(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate778(.a(G3), .O(gate389inter7));
  inv1  gate779(.a(G1042), .O(gate389inter8));
  nand2 gate780(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate781(.a(s_33), .b(gate389inter3), .O(gate389inter10));
  nor2  gate782(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate783(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate784(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1513(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1514(.a(gate397inter0), .b(s_138), .O(gate397inter1));
  and2  gate1515(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1516(.a(s_138), .O(gate397inter3));
  inv1  gate1517(.a(s_139), .O(gate397inter4));
  nand2 gate1518(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1519(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1520(.a(G11), .O(gate397inter7));
  inv1  gate1521(.a(G1066), .O(gate397inter8));
  nand2 gate1522(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1523(.a(s_139), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1524(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1525(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1526(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1079(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1080(.a(gate406inter0), .b(s_76), .O(gate406inter1));
  and2  gate1081(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1082(.a(s_76), .O(gate406inter3));
  inv1  gate1083(.a(s_77), .O(gate406inter4));
  nand2 gate1084(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1085(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1086(.a(G20), .O(gate406inter7));
  inv1  gate1087(.a(G1093), .O(gate406inter8));
  nand2 gate1088(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1089(.a(s_77), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1090(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1091(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1092(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate631(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate632(.a(gate409inter0), .b(s_12), .O(gate409inter1));
  and2  gate633(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate634(.a(s_12), .O(gate409inter3));
  inv1  gate635(.a(s_13), .O(gate409inter4));
  nand2 gate636(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate637(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate638(.a(G23), .O(gate409inter7));
  inv1  gate639(.a(G1102), .O(gate409inter8));
  nand2 gate640(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate641(.a(s_13), .b(gate409inter3), .O(gate409inter10));
  nor2  gate642(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate643(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate644(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1527(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1528(.a(gate413inter0), .b(s_140), .O(gate413inter1));
  and2  gate1529(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1530(.a(s_140), .O(gate413inter3));
  inv1  gate1531(.a(s_141), .O(gate413inter4));
  nand2 gate1532(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1533(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1534(.a(G27), .O(gate413inter7));
  inv1  gate1535(.a(G1114), .O(gate413inter8));
  nand2 gate1536(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1537(.a(s_141), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1538(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1539(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1540(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate799(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate800(.a(gate416inter0), .b(s_36), .O(gate416inter1));
  and2  gate801(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate802(.a(s_36), .O(gate416inter3));
  inv1  gate803(.a(s_37), .O(gate416inter4));
  nand2 gate804(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate805(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate806(.a(G30), .O(gate416inter7));
  inv1  gate807(.a(G1123), .O(gate416inter8));
  nand2 gate808(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate809(.a(s_37), .b(gate416inter3), .O(gate416inter10));
  nor2  gate810(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate811(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate812(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1751(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1752(.a(gate417inter0), .b(s_172), .O(gate417inter1));
  and2  gate1753(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1754(.a(s_172), .O(gate417inter3));
  inv1  gate1755(.a(s_173), .O(gate417inter4));
  nand2 gate1756(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1757(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1758(.a(G31), .O(gate417inter7));
  inv1  gate1759(.a(G1126), .O(gate417inter8));
  nand2 gate1760(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1761(.a(s_173), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1762(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1763(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1764(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1107(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1108(.a(gate421inter0), .b(s_80), .O(gate421inter1));
  and2  gate1109(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1110(.a(s_80), .O(gate421inter3));
  inv1  gate1111(.a(s_81), .O(gate421inter4));
  nand2 gate1112(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1113(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1114(.a(G2), .O(gate421inter7));
  inv1  gate1115(.a(G1135), .O(gate421inter8));
  nand2 gate1116(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1117(.a(s_81), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1118(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1119(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1120(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1653(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1654(.a(gate425inter0), .b(s_158), .O(gate425inter1));
  and2  gate1655(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1656(.a(s_158), .O(gate425inter3));
  inv1  gate1657(.a(s_159), .O(gate425inter4));
  nand2 gate1658(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1659(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1660(.a(G4), .O(gate425inter7));
  inv1  gate1661(.a(G1141), .O(gate425inter8));
  nand2 gate1662(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1663(.a(s_159), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1664(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1665(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1666(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1023(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1024(.a(gate426inter0), .b(s_68), .O(gate426inter1));
  and2  gate1025(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1026(.a(s_68), .O(gate426inter3));
  inv1  gate1027(.a(s_69), .O(gate426inter4));
  nand2 gate1028(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1029(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1030(.a(G1045), .O(gate426inter7));
  inv1  gate1031(.a(G1141), .O(gate426inter8));
  nand2 gate1032(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1033(.a(s_69), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1034(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1035(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1036(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate925(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate926(.a(gate430inter0), .b(s_54), .O(gate430inter1));
  and2  gate927(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate928(.a(s_54), .O(gate430inter3));
  inv1  gate929(.a(s_55), .O(gate430inter4));
  nand2 gate930(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate931(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate932(.a(G1051), .O(gate430inter7));
  inv1  gate933(.a(G1147), .O(gate430inter8));
  nand2 gate934(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate935(.a(s_55), .b(gate430inter3), .O(gate430inter10));
  nor2  gate936(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate937(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate938(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1121(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1122(.a(gate432inter0), .b(s_82), .O(gate432inter1));
  and2  gate1123(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1124(.a(s_82), .O(gate432inter3));
  inv1  gate1125(.a(s_83), .O(gate432inter4));
  nand2 gate1126(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1127(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1128(.a(G1054), .O(gate432inter7));
  inv1  gate1129(.a(G1150), .O(gate432inter8));
  nand2 gate1130(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1131(.a(s_83), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1132(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1133(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1134(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate729(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate730(.a(gate437inter0), .b(s_26), .O(gate437inter1));
  and2  gate731(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate732(.a(s_26), .O(gate437inter3));
  inv1  gate733(.a(s_27), .O(gate437inter4));
  nand2 gate734(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate735(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate736(.a(G10), .O(gate437inter7));
  inv1  gate737(.a(G1159), .O(gate437inter8));
  nand2 gate738(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate739(.a(s_27), .b(gate437inter3), .O(gate437inter10));
  nor2  gate740(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate741(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate742(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1303(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1304(.a(gate438inter0), .b(s_108), .O(gate438inter1));
  and2  gate1305(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1306(.a(s_108), .O(gate438inter3));
  inv1  gate1307(.a(s_109), .O(gate438inter4));
  nand2 gate1308(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1309(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1310(.a(G1063), .O(gate438inter7));
  inv1  gate1311(.a(G1159), .O(gate438inter8));
  nand2 gate1312(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1313(.a(s_109), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1314(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1315(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1316(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1709(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1710(.a(gate448inter0), .b(s_166), .O(gate448inter1));
  and2  gate1711(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1712(.a(s_166), .O(gate448inter3));
  inv1  gate1713(.a(s_167), .O(gate448inter4));
  nand2 gate1714(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1715(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1716(.a(G1078), .O(gate448inter7));
  inv1  gate1717(.a(G1174), .O(gate448inter8));
  nand2 gate1718(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1719(.a(s_167), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1720(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1721(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1722(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1807(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1808(.a(gate450inter0), .b(s_180), .O(gate450inter1));
  and2  gate1809(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1810(.a(s_180), .O(gate450inter3));
  inv1  gate1811(.a(s_181), .O(gate450inter4));
  nand2 gate1812(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1813(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1814(.a(G1081), .O(gate450inter7));
  inv1  gate1815(.a(G1177), .O(gate450inter8));
  nand2 gate1816(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1817(.a(s_181), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1818(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1819(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1820(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate813(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate814(.a(gate453inter0), .b(s_38), .O(gate453inter1));
  and2  gate815(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate816(.a(s_38), .O(gate453inter3));
  inv1  gate817(.a(s_39), .O(gate453inter4));
  nand2 gate818(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate819(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate820(.a(G18), .O(gate453inter7));
  inv1  gate821(.a(G1183), .O(gate453inter8));
  nand2 gate822(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate823(.a(s_39), .b(gate453inter3), .O(gate453inter10));
  nor2  gate824(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate825(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate826(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate617(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate618(.a(gate454inter0), .b(s_10), .O(gate454inter1));
  and2  gate619(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate620(.a(s_10), .O(gate454inter3));
  inv1  gate621(.a(s_11), .O(gate454inter4));
  nand2 gate622(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate623(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate624(.a(G1087), .O(gate454inter7));
  inv1  gate625(.a(G1183), .O(gate454inter8));
  nand2 gate626(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate627(.a(s_11), .b(gate454inter3), .O(gate454inter10));
  nor2  gate628(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate629(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate630(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1625(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1626(.a(gate460inter0), .b(s_154), .O(gate460inter1));
  and2  gate1627(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1628(.a(s_154), .O(gate460inter3));
  inv1  gate1629(.a(s_155), .O(gate460inter4));
  nand2 gate1630(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1631(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1632(.a(G1096), .O(gate460inter7));
  inv1  gate1633(.a(G1192), .O(gate460inter8));
  nand2 gate1634(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1635(.a(s_155), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1636(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1637(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1638(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate1541(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1542(.a(gate461inter0), .b(s_142), .O(gate461inter1));
  and2  gate1543(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1544(.a(s_142), .O(gate461inter3));
  inv1  gate1545(.a(s_143), .O(gate461inter4));
  nand2 gate1546(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1547(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1548(.a(G22), .O(gate461inter7));
  inv1  gate1549(.a(G1195), .O(gate461inter8));
  nand2 gate1550(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1551(.a(s_143), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1552(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1553(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1554(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1289(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1290(.a(gate481inter0), .b(s_106), .O(gate481inter1));
  and2  gate1291(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1292(.a(s_106), .O(gate481inter3));
  inv1  gate1293(.a(s_107), .O(gate481inter4));
  nand2 gate1294(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1295(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1296(.a(G32), .O(gate481inter7));
  inv1  gate1297(.a(G1225), .O(gate481inter8));
  nand2 gate1298(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1299(.a(s_107), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1300(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1301(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1302(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1317(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1318(.a(gate482inter0), .b(s_110), .O(gate482inter1));
  and2  gate1319(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1320(.a(s_110), .O(gate482inter3));
  inv1  gate1321(.a(s_111), .O(gate482inter4));
  nand2 gate1322(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1323(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1324(.a(G1129), .O(gate482inter7));
  inv1  gate1325(.a(G1225), .O(gate482inter8));
  nand2 gate1326(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1327(.a(s_111), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1328(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1329(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1330(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1499(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1500(.a(gate490inter0), .b(s_136), .O(gate490inter1));
  and2  gate1501(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1502(.a(s_136), .O(gate490inter3));
  inv1  gate1503(.a(s_137), .O(gate490inter4));
  nand2 gate1504(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1505(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1506(.a(G1242), .O(gate490inter7));
  inv1  gate1507(.a(G1243), .O(gate490inter8));
  nand2 gate1508(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1509(.a(s_137), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1510(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1511(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1512(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1191(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1192(.a(gate501inter0), .b(s_92), .O(gate501inter1));
  and2  gate1193(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1194(.a(s_92), .O(gate501inter3));
  inv1  gate1195(.a(s_93), .O(gate501inter4));
  nand2 gate1196(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1197(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1198(.a(G1264), .O(gate501inter7));
  inv1  gate1199(.a(G1265), .O(gate501inter8));
  nand2 gate1200(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1201(.a(s_93), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1202(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1203(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1204(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1037(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1038(.a(gate502inter0), .b(s_70), .O(gate502inter1));
  and2  gate1039(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1040(.a(s_70), .O(gate502inter3));
  inv1  gate1041(.a(s_71), .O(gate502inter4));
  nand2 gate1042(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1043(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1044(.a(G1266), .O(gate502inter7));
  inv1  gate1045(.a(G1267), .O(gate502inter8));
  nand2 gate1046(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1047(.a(s_71), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1048(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1049(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1050(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1429(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1430(.a(gate504inter0), .b(s_126), .O(gate504inter1));
  and2  gate1431(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1432(.a(s_126), .O(gate504inter3));
  inv1  gate1433(.a(s_127), .O(gate504inter4));
  nand2 gate1434(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1435(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1436(.a(G1270), .O(gate504inter7));
  inv1  gate1437(.a(G1271), .O(gate504inter8));
  nand2 gate1438(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1439(.a(s_127), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1440(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1441(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1442(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1051(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1052(.a(gate510inter0), .b(s_72), .O(gate510inter1));
  and2  gate1053(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1054(.a(s_72), .O(gate510inter3));
  inv1  gate1055(.a(s_73), .O(gate510inter4));
  nand2 gate1056(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1057(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1058(.a(G1282), .O(gate510inter7));
  inv1  gate1059(.a(G1283), .O(gate510inter8));
  nand2 gate1060(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1061(.a(s_73), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1062(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1063(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1064(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1177(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1178(.a(gate514inter0), .b(s_90), .O(gate514inter1));
  and2  gate1179(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1180(.a(s_90), .O(gate514inter3));
  inv1  gate1181(.a(s_91), .O(gate514inter4));
  nand2 gate1182(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1183(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1184(.a(G1290), .O(gate514inter7));
  inv1  gate1185(.a(G1291), .O(gate514inter8));
  nand2 gate1186(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1187(.a(s_91), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1188(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1189(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1190(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule