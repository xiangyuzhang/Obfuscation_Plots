module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2199(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2200(.a(gate9inter0), .b(s_236), .O(gate9inter1));
  and2  gate2201(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2202(.a(s_236), .O(gate9inter3));
  inv1  gate2203(.a(s_237), .O(gate9inter4));
  nand2 gate2204(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2205(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2206(.a(G1), .O(gate9inter7));
  inv1  gate2207(.a(G2), .O(gate9inter8));
  nand2 gate2208(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2209(.a(s_237), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2210(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2211(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2212(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2647(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2648(.a(gate13inter0), .b(s_300), .O(gate13inter1));
  and2  gate2649(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2650(.a(s_300), .O(gate13inter3));
  inv1  gate2651(.a(s_301), .O(gate13inter4));
  nand2 gate2652(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2653(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2654(.a(G9), .O(gate13inter7));
  inv1  gate2655(.a(G10), .O(gate13inter8));
  nand2 gate2656(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2657(.a(s_301), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2658(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2659(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2660(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate729(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate730(.a(gate14inter0), .b(s_26), .O(gate14inter1));
  and2  gate731(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate732(.a(s_26), .O(gate14inter3));
  inv1  gate733(.a(s_27), .O(gate14inter4));
  nand2 gate734(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate735(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate736(.a(G11), .O(gate14inter7));
  inv1  gate737(.a(G12), .O(gate14inter8));
  nand2 gate738(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate739(.a(s_27), .b(gate14inter3), .O(gate14inter10));
  nor2  gate740(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate741(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate742(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1037(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1038(.a(gate17inter0), .b(s_70), .O(gate17inter1));
  and2  gate1039(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1040(.a(s_70), .O(gate17inter3));
  inv1  gate1041(.a(s_71), .O(gate17inter4));
  nand2 gate1042(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1043(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1044(.a(G17), .O(gate17inter7));
  inv1  gate1045(.a(G18), .O(gate17inter8));
  nand2 gate1046(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1047(.a(s_71), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1048(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1049(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1050(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1457(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1458(.a(gate20inter0), .b(s_130), .O(gate20inter1));
  and2  gate1459(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1460(.a(s_130), .O(gate20inter3));
  inv1  gate1461(.a(s_131), .O(gate20inter4));
  nand2 gate1462(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1463(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1464(.a(G23), .O(gate20inter7));
  inv1  gate1465(.a(G24), .O(gate20inter8));
  nand2 gate1466(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1467(.a(s_131), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1468(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1469(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1470(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2017(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2018(.a(gate24inter0), .b(s_210), .O(gate24inter1));
  and2  gate2019(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2020(.a(s_210), .O(gate24inter3));
  inv1  gate2021(.a(s_211), .O(gate24inter4));
  nand2 gate2022(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2023(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2024(.a(G31), .O(gate24inter7));
  inv1  gate2025(.a(G32), .O(gate24inter8));
  nand2 gate2026(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2027(.a(s_211), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2028(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2029(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2030(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2437(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2438(.a(gate28inter0), .b(s_270), .O(gate28inter1));
  and2  gate2439(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2440(.a(s_270), .O(gate28inter3));
  inv1  gate2441(.a(s_271), .O(gate28inter4));
  nand2 gate2442(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2443(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2444(.a(G10), .O(gate28inter7));
  inv1  gate2445(.a(G14), .O(gate28inter8));
  nand2 gate2446(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2447(.a(s_271), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2448(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2449(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2450(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1793(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1794(.a(gate30inter0), .b(s_178), .O(gate30inter1));
  and2  gate1795(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1796(.a(s_178), .O(gate30inter3));
  inv1  gate1797(.a(s_179), .O(gate30inter4));
  nand2 gate1798(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1799(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1800(.a(G11), .O(gate30inter7));
  inv1  gate1801(.a(G15), .O(gate30inter8));
  nand2 gate1802(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1803(.a(s_179), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1804(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1805(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1806(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1471(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1472(.a(gate31inter0), .b(s_132), .O(gate31inter1));
  and2  gate1473(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1474(.a(s_132), .O(gate31inter3));
  inv1  gate1475(.a(s_133), .O(gate31inter4));
  nand2 gate1476(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1477(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1478(.a(G4), .O(gate31inter7));
  inv1  gate1479(.a(G8), .O(gate31inter8));
  nand2 gate1480(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1481(.a(s_133), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1482(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1483(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1484(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate561(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate562(.a(gate33inter0), .b(s_2), .O(gate33inter1));
  and2  gate563(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate564(.a(s_2), .O(gate33inter3));
  inv1  gate565(.a(s_3), .O(gate33inter4));
  nand2 gate566(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate567(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate568(.a(G17), .O(gate33inter7));
  inv1  gate569(.a(G21), .O(gate33inter8));
  nand2 gate570(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate571(.a(s_3), .b(gate33inter3), .O(gate33inter10));
  nor2  gate572(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate573(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate574(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2759(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2760(.a(gate34inter0), .b(s_316), .O(gate34inter1));
  and2  gate2761(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2762(.a(s_316), .O(gate34inter3));
  inv1  gate2763(.a(s_317), .O(gate34inter4));
  nand2 gate2764(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2765(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2766(.a(G25), .O(gate34inter7));
  inv1  gate2767(.a(G29), .O(gate34inter8));
  nand2 gate2768(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2769(.a(s_317), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2770(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2771(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2772(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1373(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1374(.a(gate35inter0), .b(s_118), .O(gate35inter1));
  and2  gate1375(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1376(.a(s_118), .O(gate35inter3));
  inv1  gate1377(.a(s_119), .O(gate35inter4));
  nand2 gate1378(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1379(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1380(.a(G18), .O(gate35inter7));
  inv1  gate1381(.a(G22), .O(gate35inter8));
  nand2 gate1382(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1383(.a(s_119), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1384(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1385(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1386(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate981(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate982(.a(gate37inter0), .b(s_62), .O(gate37inter1));
  and2  gate983(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate984(.a(s_62), .O(gate37inter3));
  inv1  gate985(.a(s_63), .O(gate37inter4));
  nand2 gate986(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate987(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate988(.a(G19), .O(gate37inter7));
  inv1  gate989(.a(G23), .O(gate37inter8));
  nand2 gate990(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate991(.a(s_63), .b(gate37inter3), .O(gate37inter10));
  nor2  gate992(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate993(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate994(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1639(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1640(.a(gate38inter0), .b(s_156), .O(gate38inter1));
  and2  gate1641(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1642(.a(s_156), .O(gate38inter3));
  inv1  gate1643(.a(s_157), .O(gate38inter4));
  nand2 gate1644(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1645(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1646(.a(G27), .O(gate38inter7));
  inv1  gate1647(.a(G31), .O(gate38inter8));
  nand2 gate1648(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1649(.a(s_157), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1650(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1651(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1652(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1569(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1570(.a(gate39inter0), .b(s_146), .O(gate39inter1));
  and2  gate1571(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1572(.a(s_146), .O(gate39inter3));
  inv1  gate1573(.a(s_147), .O(gate39inter4));
  nand2 gate1574(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1575(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1576(.a(G20), .O(gate39inter7));
  inv1  gate1577(.a(G24), .O(gate39inter8));
  nand2 gate1578(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1579(.a(s_147), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1580(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1581(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1582(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1317(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1318(.a(gate41inter0), .b(s_110), .O(gate41inter1));
  and2  gate1319(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1320(.a(s_110), .O(gate41inter3));
  inv1  gate1321(.a(s_111), .O(gate41inter4));
  nand2 gate1322(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1323(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1324(.a(G1), .O(gate41inter7));
  inv1  gate1325(.a(G266), .O(gate41inter8));
  nand2 gate1326(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1327(.a(s_111), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1328(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1329(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1330(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2479(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2480(.a(gate46inter0), .b(s_276), .O(gate46inter1));
  and2  gate2481(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2482(.a(s_276), .O(gate46inter3));
  inv1  gate2483(.a(s_277), .O(gate46inter4));
  nand2 gate2484(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2485(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2486(.a(G6), .O(gate46inter7));
  inv1  gate2487(.a(G272), .O(gate46inter8));
  nand2 gate2488(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2489(.a(s_277), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2490(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2491(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2492(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2927(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2928(.a(gate47inter0), .b(s_340), .O(gate47inter1));
  and2  gate2929(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2930(.a(s_340), .O(gate47inter3));
  inv1  gate2931(.a(s_341), .O(gate47inter4));
  nand2 gate2932(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2933(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2934(.a(G7), .O(gate47inter7));
  inv1  gate2935(.a(G275), .O(gate47inter8));
  nand2 gate2936(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2937(.a(s_341), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2938(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2939(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2940(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1625(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1626(.a(gate48inter0), .b(s_154), .O(gate48inter1));
  and2  gate1627(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1628(.a(s_154), .O(gate48inter3));
  inv1  gate1629(.a(s_155), .O(gate48inter4));
  nand2 gate1630(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1631(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1632(.a(G8), .O(gate48inter7));
  inv1  gate1633(.a(G275), .O(gate48inter8));
  nand2 gate1634(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1635(.a(s_155), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1636(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1637(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1638(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1051(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1052(.a(gate49inter0), .b(s_72), .O(gate49inter1));
  and2  gate1053(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1054(.a(s_72), .O(gate49inter3));
  inv1  gate1055(.a(s_73), .O(gate49inter4));
  nand2 gate1056(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1057(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1058(.a(G9), .O(gate49inter7));
  inv1  gate1059(.a(G278), .O(gate49inter8));
  nand2 gate1060(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1061(.a(s_73), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1062(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1063(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1064(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate575(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate576(.a(gate52inter0), .b(s_4), .O(gate52inter1));
  and2  gate577(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate578(.a(s_4), .O(gate52inter3));
  inv1  gate579(.a(s_5), .O(gate52inter4));
  nand2 gate580(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate581(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate582(.a(G12), .O(gate52inter7));
  inv1  gate583(.a(G281), .O(gate52inter8));
  nand2 gate584(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate585(.a(s_5), .b(gate52inter3), .O(gate52inter10));
  nor2  gate586(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate587(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate588(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2731(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2732(.a(gate54inter0), .b(s_312), .O(gate54inter1));
  and2  gate2733(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2734(.a(s_312), .O(gate54inter3));
  inv1  gate2735(.a(s_313), .O(gate54inter4));
  nand2 gate2736(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2737(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2738(.a(G14), .O(gate54inter7));
  inv1  gate2739(.a(G284), .O(gate54inter8));
  nand2 gate2740(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2741(.a(s_313), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2742(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2743(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2744(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate883(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate884(.a(gate57inter0), .b(s_48), .O(gate57inter1));
  and2  gate885(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate886(.a(s_48), .O(gate57inter3));
  inv1  gate887(.a(s_49), .O(gate57inter4));
  nand2 gate888(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate889(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate890(.a(G17), .O(gate57inter7));
  inv1  gate891(.a(G290), .O(gate57inter8));
  nand2 gate892(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate893(.a(s_49), .b(gate57inter3), .O(gate57inter10));
  nor2  gate894(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate895(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate896(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate939(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate940(.a(gate58inter0), .b(s_56), .O(gate58inter1));
  and2  gate941(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate942(.a(s_56), .O(gate58inter3));
  inv1  gate943(.a(s_57), .O(gate58inter4));
  nand2 gate944(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate945(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate946(.a(G18), .O(gate58inter7));
  inv1  gate947(.a(G290), .O(gate58inter8));
  nand2 gate948(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate949(.a(s_57), .b(gate58inter3), .O(gate58inter10));
  nor2  gate950(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate951(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate952(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate645(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate646(.a(gate62inter0), .b(s_14), .O(gate62inter1));
  and2  gate647(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate648(.a(s_14), .O(gate62inter3));
  inv1  gate649(.a(s_15), .O(gate62inter4));
  nand2 gate650(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate651(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate652(.a(G22), .O(gate62inter7));
  inv1  gate653(.a(G296), .O(gate62inter8));
  nand2 gate654(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate655(.a(s_15), .b(gate62inter3), .O(gate62inter10));
  nor2  gate656(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate657(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate658(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2913(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2914(.a(gate66inter0), .b(s_338), .O(gate66inter1));
  and2  gate2915(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2916(.a(s_338), .O(gate66inter3));
  inv1  gate2917(.a(s_339), .O(gate66inter4));
  nand2 gate2918(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2919(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2920(.a(G26), .O(gate66inter7));
  inv1  gate2921(.a(G302), .O(gate66inter8));
  nand2 gate2922(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2923(.a(s_339), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2924(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2925(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2926(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1555(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1556(.a(gate68inter0), .b(s_144), .O(gate68inter1));
  and2  gate1557(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1558(.a(s_144), .O(gate68inter3));
  inv1  gate1559(.a(s_145), .O(gate68inter4));
  nand2 gate1560(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1561(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1562(.a(G28), .O(gate68inter7));
  inv1  gate1563(.a(G305), .O(gate68inter8));
  nand2 gate1564(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1565(.a(s_145), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1566(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1567(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1568(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate631(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate632(.a(gate69inter0), .b(s_12), .O(gate69inter1));
  and2  gate633(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate634(.a(s_12), .O(gate69inter3));
  inv1  gate635(.a(s_13), .O(gate69inter4));
  nand2 gate636(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate637(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate638(.a(G29), .O(gate69inter7));
  inv1  gate639(.a(G308), .O(gate69inter8));
  nand2 gate640(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate641(.a(s_13), .b(gate69inter3), .O(gate69inter10));
  nor2  gate642(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate643(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate644(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1303(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1304(.a(gate70inter0), .b(s_108), .O(gate70inter1));
  and2  gate1305(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1306(.a(s_108), .O(gate70inter3));
  inv1  gate1307(.a(s_109), .O(gate70inter4));
  nand2 gate1308(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1309(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1310(.a(G30), .O(gate70inter7));
  inv1  gate1311(.a(G308), .O(gate70inter8));
  nand2 gate1312(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1313(.a(s_109), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1314(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1315(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1316(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1079(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1080(.a(gate71inter0), .b(s_76), .O(gate71inter1));
  and2  gate1081(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1082(.a(s_76), .O(gate71inter3));
  inv1  gate1083(.a(s_77), .O(gate71inter4));
  nand2 gate1084(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1085(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1086(.a(G31), .O(gate71inter7));
  inv1  gate1087(.a(G311), .O(gate71inter8));
  nand2 gate1088(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1089(.a(s_77), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1090(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1091(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1092(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1891(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1892(.a(gate72inter0), .b(s_192), .O(gate72inter1));
  and2  gate1893(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1894(.a(s_192), .O(gate72inter3));
  inv1  gate1895(.a(s_193), .O(gate72inter4));
  nand2 gate1896(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1897(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1898(.a(G32), .O(gate72inter7));
  inv1  gate1899(.a(G311), .O(gate72inter8));
  nand2 gate1900(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1901(.a(s_193), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1902(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1903(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1904(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate2899(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2900(.a(gate73inter0), .b(s_336), .O(gate73inter1));
  and2  gate2901(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2902(.a(s_336), .O(gate73inter3));
  inv1  gate2903(.a(s_337), .O(gate73inter4));
  nand2 gate2904(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2905(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2906(.a(G1), .O(gate73inter7));
  inv1  gate2907(.a(G314), .O(gate73inter8));
  nand2 gate2908(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2909(.a(s_337), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2910(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2911(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2912(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1415(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1416(.a(gate75inter0), .b(s_124), .O(gate75inter1));
  and2  gate1417(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1418(.a(s_124), .O(gate75inter3));
  inv1  gate1419(.a(s_125), .O(gate75inter4));
  nand2 gate1420(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1421(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1422(.a(G9), .O(gate75inter7));
  inv1  gate1423(.a(G317), .O(gate75inter8));
  nand2 gate1424(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1425(.a(s_125), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1426(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1427(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1428(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1709(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1710(.a(gate78inter0), .b(s_166), .O(gate78inter1));
  and2  gate1711(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1712(.a(s_166), .O(gate78inter3));
  inv1  gate1713(.a(s_167), .O(gate78inter4));
  nand2 gate1714(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1715(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1716(.a(G6), .O(gate78inter7));
  inv1  gate1717(.a(G320), .O(gate78inter8));
  nand2 gate1718(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1719(.a(s_167), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1720(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1721(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1722(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2871(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2872(.a(gate82inter0), .b(s_332), .O(gate82inter1));
  and2  gate2873(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2874(.a(s_332), .O(gate82inter3));
  inv1  gate2875(.a(s_333), .O(gate82inter4));
  nand2 gate2876(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2877(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2878(.a(G7), .O(gate82inter7));
  inv1  gate2879(.a(G326), .O(gate82inter8));
  nand2 gate2880(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2881(.a(s_333), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2882(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2883(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2884(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1093(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1094(.a(gate88inter0), .b(s_78), .O(gate88inter1));
  and2  gate1095(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1096(.a(s_78), .O(gate88inter3));
  inv1  gate1097(.a(s_79), .O(gate88inter4));
  nand2 gate1098(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1099(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1100(.a(G16), .O(gate88inter7));
  inv1  gate1101(.a(G335), .O(gate88inter8));
  nand2 gate1102(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1103(.a(s_79), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1104(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1105(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1106(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate995(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate996(.a(gate89inter0), .b(s_64), .O(gate89inter1));
  and2  gate997(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate998(.a(s_64), .O(gate89inter3));
  inv1  gate999(.a(s_65), .O(gate89inter4));
  nand2 gate1000(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1001(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1002(.a(G17), .O(gate89inter7));
  inv1  gate1003(.a(G338), .O(gate89inter8));
  nand2 gate1004(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1005(.a(s_65), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1006(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1007(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1008(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1247(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1248(.a(gate91inter0), .b(s_100), .O(gate91inter1));
  and2  gate1249(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1250(.a(s_100), .O(gate91inter3));
  inv1  gate1251(.a(s_101), .O(gate91inter4));
  nand2 gate1252(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1253(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1254(.a(G25), .O(gate91inter7));
  inv1  gate1255(.a(G341), .O(gate91inter8));
  nand2 gate1256(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1257(.a(s_101), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1258(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1259(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1260(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate925(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate926(.a(gate95inter0), .b(s_54), .O(gate95inter1));
  and2  gate927(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate928(.a(s_54), .O(gate95inter3));
  inv1  gate929(.a(s_55), .O(gate95inter4));
  nand2 gate930(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate931(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate932(.a(G26), .O(gate95inter7));
  inv1  gate933(.a(G347), .O(gate95inter8));
  nand2 gate934(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate935(.a(s_55), .b(gate95inter3), .O(gate95inter10));
  nor2  gate936(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate937(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate938(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2059(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2060(.a(gate96inter0), .b(s_216), .O(gate96inter1));
  and2  gate2061(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2062(.a(s_216), .O(gate96inter3));
  inv1  gate2063(.a(s_217), .O(gate96inter4));
  nand2 gate2064(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2065(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2066(.a(G30), .O(gate96inter7));
  inv1  gate2067(.a(G347), .O(gate96inter8));
  nand2 gate2068(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2069(.a(s_217), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2070(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2071(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2072(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1205(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1206(.a(gate97inter0), .b(s_94), .O(gate97inter1));
  and2  gate1207(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1208(.a(s_94), .O(gate97inter3));
  inv1  gate1209(.a(s_95), .O(gate97inter4));
  nand2 gate1210(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1211(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1212(.a(G19), .O(gate97inter7));
  inv1  gate1213(.a(G350), .O(gate97inter8));
  nand2 gate1214(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1215(.a(s_95), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1216(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1217(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1218(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate869(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate870(.a(gate100inter0), .b(s_46), .O(gate100inter1));
  and2  gate871(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate872(.a(s_46), .O(gate100inter3));
  inv1  gate873(.a(s_47), .O(gate100inter4));
  nand2 gate874(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate875(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate876(.a(G31), .O(gate100inter7));
  inv1  gate877(.a(G353), .O(gate100inter8));
  nand2 gate878(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate879(.a(s_47), .b(gate100inter3), .O(gate100inter10));
  nor2  gate880(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate881(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate882(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate911(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate912(.a(gate110inter0), .b(s_52), .O(gate110inter1));
  and2  gate913(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate914(.a(s_52), .O(gate110inter3));
  inv1  gate915(.a(s_53), .O(gate110inter4));
  nand2 gate916(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate917(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate918(.a(G372), .O(gate110inter7));
  inv1  gate919(.a(G373), .O(gate110inter8));
  nand2 gate920(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate921(.a(s_53), .b(gate110inter3), .O(gate110inter10));
  nor2  gate922(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate923(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate924(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2661(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2662(.a(gate111inter0), .b(s_302), .O(gate111inter1));
  and2  gate2663(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2664(.a(s_302), .O(gate111inter3));
  inv1  gate2665(.a(s_303), .O(gate111inter4));
  nand2 gate2666(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2667(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2668(.a(G374), .O(gate111inter7));
  inv1  gate2669(.a(G375), .O(gate111inter8));
  nand2 gate2670(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2671(.a(s_303), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2672(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2673(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2674(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2619(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2620(.a(gate112inter0), .b(s_296), .O(gate112inter1));
  and2  gate2621(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2622(.a(s_296), .O(gate112inter3));
  inv1  gate2623(.a(s_297), .O(gate112inter4));
  nand2 gate2624(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2625(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2626(.a(G376), .O(gate112inter7));
  inv1  gate2627(.a(G377), .O(gate112inter8));
  nand2 gate2628(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2629(.a(s_297), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2630(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2631(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2632(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1065(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1066(.a(gate116inter0), .b(s_74), .O(gate116inter1));
  and2  gate1067(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1068(.a(s_74), .O(gate116inter3));
  inv1  gate1069(.a(s_75), .O(gate116inter4));
  nand2 gate1070(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1071(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1072(.a(G384), .O(gate116inter7));
  inv1  gate1073(.a(G385), .O(gate116inter8));
  nand2 gate1074(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1075(.a(s_75), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1076(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1077(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1078(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate603(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate604(.a(gate124inter0), .b(s_8), .O(gate124inter1));
  and2  gate605(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate606(.a(s_8), .O(gate124inter3));
  inv1  gate607(.a(s_9), .O(gate124inter4));
  nand2 gate608(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate609(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate610(.a(G400), .O(gate124inter7));
  inv1  gate611(.a(G401), .O(gate124inter8));
  nand2 gate612(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate613(.a(s_9), .b(gate124inter3), .O(gate124inter10));
  nor2  gate614(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate615(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate616(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate897(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate898(.a(gate126inter0), .b(s_50), .O(gate126inter1));
  and2  gate899(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate900(.a(s_50), .O(gate126inter3));
  inv1  gate901(.a(s_51), .O(gate126inter4));
  nand2 gate902(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate903(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate904(.a(G404), .O(gate126inter7));
  inv1  gate905(.a(G405), .O(gate126inter8));
  nand2 gate906(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate907(.a(s_51), .b(gate126inter3), .O(gate126inter10));
  nor2  gate908(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate909(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate910(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2605(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2606(.a(gate131inter0), .b(s_294), .O(gate131inter1));
  and2  gate2607(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2608(.a(s_294), .O(gate131inter3));
  inv1  gate2609(.a(s_295), .O(gate131inter4));
  nand2 gate2610(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2611(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2612(.a(G414), .O(gate131inter7));
  inv1  gate2613(.a(G415), .O(gate131inter8));
  nand2 gate2614(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2615(.a(s_295), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2616(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2617(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2618(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1401(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1402(.a(gate132inter0), .b(s_122), .O(gate132inter1));
  and2  gate1403(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1404(.a(s_122), .O(gate132inter3));
  inv1  gate1405(.a(s_123), .O(gate132inter4));
  nand2 gate1406(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1407(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1408(.a(G416), .O(gate132inter7));
  inv1  gate1409(.a(G417), .O(gate132inter8));
  nand2 gate1410(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1411(.a(s_123), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1412(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1413(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1414(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1947(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1948(.a(gate133inter0), .b(s_200), .O(gate133inter1));
  and2  gate1949(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1950(.a(s_200), .O(gate133inter3));
  inv1  gate1951(.a(s_201), .O(gate133inter4));
  nand2 gate1952(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1953(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1954(.a(G418), .O(gate133inter7));
  inv1  gate1955(.a(G419), .O(gate133inter8));
  nand2 gate1956(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1957(.a(s_201), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1958(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1959(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1960(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate2717(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2718(.a(gate134inter0), .b(s_310), .O(gate134inter1));
  and2  gate2719(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2720(.a(s_310), .O(gate134inter3));
  inv1  gate2721(.a(s_311), .O(gate134inter4));
  nand2 gate2722(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2723(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2724(.a(G420), .O(gate134inter7));
  inv1  gate2725(.a(G421), .O(gate134inter8));
  nand2 gate2726(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2727(.a(s_311), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2728(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2729(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2730(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2045(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2046(.a(gate137inter0), .b(s_214), .O(gate137inter1));
  and2  gate2047(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2048(.a(s_214), .O(gate137inter3));
  inv1  gate2049(.a(s_215), .O(gate137inter4));
  nand2 gate2050(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2051(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2052(.a(G426), .O(gate137inter7));
  inv1  gate2053(.a(G429), .O(gate137inter8));
  nand2 gate2054(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2055(.a(s_215), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2056(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2057(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2058(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2311(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2312(.a(gate140inter0), .b(s_252), .O(gate140inter1));
  and2  gate2313(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2314(.a(s_252), .O(gate140inter3));
  inv1  gate2315(.a(s_253), .O(gate140inter4));
  nand2 gate2316(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2317(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2318(.a(G444), .O(gate140inter7));
  inv1  gate2319(.a(G447), .O(gate140inter8));
  nand2 gate2320(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2321(.a(s_253), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2322(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2323(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2324(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1289(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1290(.a(gate144inter0), .b(s_106), .O(gate144inter1));
  and2  gate1291(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1292(.a(s_106), .O(gate144inter3));
  inv1  gate1293(.a(s_107), .O(gate144inter4));
  nand2 gate1294(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1295(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1296(.a(G468), .O(gate144inter7));
  inv1  gate1297(.a(G471), .O(gate144inter8));
  nand2 gate1298(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1299(.a(s_107), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1300(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1301(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1302(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2087(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2088(.a(gate146inter0), .b(s_220), .O(gate146inter1));
  and2  gate2089(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2090(.a(s_220), .O(gate146inter3));
  inv1  gate2091(.a(s_221), .O(gate146inter4));
  nand2 gate2092(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2093(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2094(.a(G480), .O(gate146inter7));
  inv1  gate2095(.a(G483), .O(gate146inter8));
  nand2 gate2096(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2097(.a(s_221), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2098(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2099(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2100(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2521(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2522(.a(gate147inter0), .b(s_282), .O(gate147inter1));
  and2  gate2523(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2524(.a(s_282), .O(gate147inter3));
  inv1  gate2525(.a(s_283), .O(gate147inter4));
  nand2 gate2526(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2527(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2528(.a(G486), .O(gate147inter7));
  inv1  gate2529(.a(G489), .O(gate147inter8));
  nand2 gate2530(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2531(.a(s_283), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2532(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2533(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2534(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2031(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2032(.a(gate153inter0), .b(s_212), .O(gate153inter1));
  and2  gate2033(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2034(.a(s_212), .O(gate153inter3));
  inv1  gate2035(.a(s_213), .O(gate153inter4));
  nand2 gate2036(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2037(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2038(.a(G426), .O(gate153inter7));
  inv1  gate2039(.a(G522), .O(gate153inter8));
  nand2 gate2040(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2041(.a(s_213), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2042(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2043(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2044(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1513(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1514(.a(gate155inter0), .b(s_138), .O(gate155inter1));
  and2  gate1515(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1516(.a(s_138), .O(gate155inter3));
  inv1  gate1517(.a(s_139), .O(gate155inter4));
  nand2 gate1518(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1519(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1520(.a(G432), .O(gate155inter7));
  inv1  gate1521(.a(G525), .O(gate155inter8));
  nand2 gate1522(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1523(.a(s_139), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1524(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1525(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1526(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2227(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2228(.a(gate157inter0), .b(s_240), .O(gate157inter1));
  and2  gate2229(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2230(.a(s_240), .O(gate157inter3));
  inv1  gate2231(.a(s_241), .O(gate157inter4));
  nand2 gate2232(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2233(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2234(.a(G438), .O(gate157inter7));
  inv1  gate2235(.a(G528), .O(gate157inter8));
  nand2 gate2236(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2237(.a(s_241), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2238(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2239(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2240(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2157(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2158(.a(gate162inter0), .b(s_230), .O(gate162inter1));
  and2  gate2159(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2160(.a(s_230), .O(gate162inter3));
  inv1  gate2161(.a(s_231), .O(gate162inter4));
  nand2 gate2162(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2163(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2164(.a(G453), .O(gate162inter7));
  inv1  gate2165(.a(G534), .O(gate162inter8));
  nand2 gate2166(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2167(.a(s_231), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2168(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2169(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2170(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2185(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2186(.a(gate163inter0), .b(s_234), .O(gate163inter1));
  and2  gate2187(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2188(.a(s_234), .O(gate163inter3));
  inv1  gate2189(.a(s_235), .O(gate163inter4));
  nand2 gate2190(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2191(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2192(.a(G456), .O(gate163inter7));
  inv1  gate2193(.a(G537), .O(gate163inter8));
  nand2 gate2194(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2195(.a(s_235), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2196(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2197(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2198(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2829(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2830(.a(gate167inter0), .b(s_326), .O(gate167inter1));
  and2  gate2831(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2832(.a(s_326), .O(gate167inter3));
  inv1  gate2833(.a(s_327), .O(gate167inter4));
  nand2 gate2834(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2835(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2836(.a(G468), .O(gate167inter7));
  inv1  gate2837(.a(G543), .O(gate167inter8));
  nand2 gate2838(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2839(.a(s_327), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2840(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2841(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2842(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate2633(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2634(.a(gate168inter0), .b(s_298), .O(gate168inter1));
  and2  gate2635(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2636(.a(s_298), .O(gate168inter3));
  inv1  gate2637(.a(s_299), .O(gate168inter4));
  nand2 gate2638(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2639(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2640(.a(G471), .O(gate168inter7));
  inv1  gate2641(.a(G543), .O(gate168inter8));
  nand2 gate2642(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2643(.a(s_299), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2644(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2645(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2646(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2353(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2354(.a(gate174inter0), .b(s_258), .O(gate174inter1));
  and2  gate2355(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2356(.a(s_258), .O(gate174inter3));
  inv1  gate2357(.a(s_259), .O(gate174inter4));
  nand2 gate2358(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2359(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2360(.a(G489), .O(gate174inter7));
  inv1  gate2361(.a(G552), .O(gate174inter8));
  nand2 gate2362(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2363(.a(s_259), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2364(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2365(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2366(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2073(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2074(.a(gate175inter0), .b(s_218), .O(gate175inter1));
  and2  gate2075(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2076(.a(s_218), .O(gate175inter3));
  inv1  gate2077(.a(s_219), .O(gate175inter4));
  nand2 gate2078(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2079(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2080(.a(G492), .O(gate175inter7));
  inv1  gate2081(.a(G555), .O(gate175inter8));
  nand2 gate2082(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2083(.a(s_219), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2084(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2085(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2086(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate967(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate968(.a(gate180inter0), .b(s_60), .O(gate180inter1));
  and2  gate969(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate970(.a(s_60), .O(gate180inter3));
  inv1  gate971(.a(s_61), .O(gate180inter4));
  nand2 gate972(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate973(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate974(.a(G507), .O(gate180inter7));
  inv1  gate975(.a(G561), .O(gate180inter8));
  nand2 gate976(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate977(.a(s_61), .b(gate180inter3), .O(gate180inter10));
  nor2  gate978(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate979(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate980(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1233(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1234(.a(gate181inter0), .b(s_98), .O(gate181inter1));
  and2  gate1235(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1236(.a(s_98), .O(gate181inter3));
  inv1  gate1237(.a(s_99), .O(gate181inter4));
  nand2 gate1238(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1239(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1240(.a(G510), .O(gate181inter7));
  inv1  gate1241(.a(G564), .O(gate181inter8));
  nand2 gate1242(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1243(.a(s_99), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1244(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1245(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1246(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1191(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1192(.a(gate182inter0), .b(s_92), .O(gate182inter1));
  and2  gate1193(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1194(.a(s_92), .O(gate182inter3));
  inv1  gate1195(.a(s_93), .O(gate182inter4));
  nand2 gate1196(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1197(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1198(.a(G513), .O(gate182inter7));
  inv1  gate1199(.a(G564), .O(gate182inter8));
  nand2 gate1200(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1201(.a(s_93), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1202(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1203(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1204(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1751(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1752(.a(gate183inter0), .b(s_172), .O(gate183inter1));
  and2  gate1753(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1754(.a(s_172), .O(gate183inter3));
  inv1  gate1755(.a(s_173), .O(gate183inter4));
  nand2 gate1756(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1757(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1758(.a(G516), .O(gate183inter7));
  inv1  gate1759(.a(G567), .O(gate183inter8));
  nand2 gate1760(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1761(.a(s_173), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1762(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1763(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1764(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1961(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1962(.a(gate185inter0), .b(s_202), .O(gate185inter1));
  and2  gate1963(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1964(.a(s_202), .O(gate185inter3));
  inv1  gate1965(.a(s_203), .O(gate185inter4));
  nand2 gate1966(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1967(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1968(.a(G570), .O(gate185inter7));
  inv1  gate1969(.a(G571), .O(gate185inter8));
  nand2 gate1970(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1971(.a(s_203), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1972(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1973(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1974(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate715(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate716(.a(gate187inter0), .b(s_24), .O(gate187inter1));
  and2  gate717(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate718(.a(s_24), .O(gate187inter3));
  inv1  gate719(.a(s_25), .O(gate187inter4));
  nand2 gate720(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate721(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate722(.a(G574), .O(gate187inter7));
  inv1  gate723(.a(G575), .O(gate187inter8));
  nand2 gate724(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate725(.a(s_25), .b(gate187inter3), .O(gate187inter10));
  nor2  gate726(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate727(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate728(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1695(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1696(.a(gate191inter0), .b(s_164), .O(gate191inter1));
  and2  gate1697(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1698(.a(s_164), .O(gate191inter3));
  inv1  gate1699(.a(s_165), .O(gate191inter4));
  nand2 gate1700(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1701(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1702(.a(G582), .O(gate191inter7));
  inv1  gate1703(.a(G583), .O(gate191inter8));
  nand2 gate1704(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1705(.a(s_165), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1706(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1707(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1708(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2535(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2536(.a(gate192inter0), .b(s_284), .O(gate192inter1));
  and2  gate2537(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2538(.a(s_284), .O(gate192inter3));
  inv1  gate2539(.a(s_285), .O(gate192inter4));
  nand2 gate2540(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2541(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2542(.a(G584), .O(gate192inter7));
  inv1  gate2543(.a(G585), .O(gate192inter8));
  nand2 gate2544(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2545(.a(s_285), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2546(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2547(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2548(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1485(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1486(.a(gate195inter0), .b(s_134), .O(gate195inter1));
  and2  gate1487(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1488(.a(s_134), .O(gate195inter3));
  inv1  gate1489(.a(s_135), .O(gate195inter4));
  nand2 gate1490(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1491(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1492(.a(G590), .O(gate195inter7));
  inv1  gate1493(.a(G591), .O(gate195inter8));
  nand2 gate1494(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1495(.a(s_135), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1496(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1497(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1498(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2339(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2340(.a(gate196inter0), .b(s_256), .O(gate196inter1));
  and2  gate2341(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2342(.a(s_256), .O(gate196inter3));
  inv1  gate2343(.a(s_257), .O(gate196inter4));
  nand2 gate2344(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2345(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2346(.a(G592), .O(gate196inter7));
  inv1  gate2347(.a(G593), .O(gate196inter8));
  nand2 gate2348(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2349(.a(s_257), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2350(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2351(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2352(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1849(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1850(.a(gate198inter0), .b(s_186), .O(gate198inter1));
  and2  gate1851(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1852(.a(s_186), .O(gate198inter3));
  inv1  gate1853(.a(s_187), .O(gate198inter4));
  nand2 gate1854(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1855(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1856(.a(G596), .O(gate198inter7));
  inv1  gate1857(.a(G597), .O(gate198inter8));
  nand2 gate1858(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1859(.a(s_187), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1860(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1861(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1862(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2423(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2424(.a(gate199inter0), .b(s_268), .O(gate199inter1));
  and2  gate2425(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2426(.a(s_268), .O(gate199inter3));
  inv1  gate2427(.a(s_269), .O(gate199inter4));
  nand2 gate2428(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2429(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2430(.a(G598), .O(gate199inter7));
  inv1  gate2431(.a(G599), .O(gate199inter8));
  nand2 gate2432(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2433(.a(s_269), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2434(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2435(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2436(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2451(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2452(.a(gate204inter0), .b(s_272), .O(gate204inter1));
  and2  gate2453(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2454(.a(s_272), .O(gate204inter3));
  inv1  gate2455(.a(s_273), .O(gate204inter4));
  nand2 gate2456(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2457(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2458(.a(G607), .O(gate204inter7));
  inv1  gate2459(.a(G617), .O(gate204inter8));
  nand2 gate2460(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2461(.a(s_273), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2462(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2463(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2464(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1163(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1164(.a(gate206inter0), .b(s_88), .O(gate206inter1));
  and2  gate1165(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1166(.a(s_88), .O(gate206inter3));
  inv1  gate1167(.a(s_89), .O(gate206inter4));
  nand2 gate1168(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1169(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1170(.a(G632), .O(gate206inter7));
  inv1  gate1171(.a(G637), .O(gate206inter8));
  nand2 gate1172(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1173(.a(s_89), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1174(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1175(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1176(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2773(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2774(.a(gate208inter0), .b(s_318), .O(gate208inter1));
  and2  gate2775(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2776(.a(s_318), .O(gate208inter3));
  inv1  gate2777(.a(s_319), .O(gate208inter4));
  nand2 gate2778(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2779(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2780(.a(G627), .O(gate208inter7));
  inv1  gate2781(.a(G637), .O(gate208inter8));
  nand2 gate2782(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2783(.a(s_319), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2784(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2785(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2786(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1135(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1136(.a(gate210inter0), .b(s_84), .O(gate210inter1));
  and2  gate1137(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1138(.a(s_84), .O(gate210inter3));
  inv1  gate1139(.a(s_85), .O(gate210inter4));
  nand2 gate1140(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1141(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1142(.a(G607), .O(gate210inter7));
  inv1  gate1143(.a(G666), .O(gate210inter8));
  nand2 gate1144(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1145(.a(s_85), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1146(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1147(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1148(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1597(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1598(.a(gate211inter0), .b(s_150), .O(gate211inter1));
  and2  gate1599(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1600(.a(s_150), .O(gate211inter3));
  inv1  gate1601(.a(s_151), .O(gate211inter4));
  nand2 gate1602(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1603(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1604(.a(G612), .O(gate211inter7));
  inv1  gate1605(.a(G669), .O(gate211inter8));
  nand2 gate1606(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1607(.a(s_151), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1608(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1609(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1610(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1009(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1010(.a(gate214inter0), .b(s_66), .O(gate214inter1));
  and2  gate1011(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1012(.a(s_66), .O(gate214inter3));
  inv1  gate1013(.a(s_67), .O(gate214inter4));
  nand2 gate1014(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1015(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1016(.a(G612), .O(gate214inter7));
  inv1  gate1017(.a(G672), .O(gate214inter8));
  nand2 gate1018(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1019(.a(s_67), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1020(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1021(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1022(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1443(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1444(.a(gate215inter0), .b(s_128), .O(gate215inter1));
  and2  gate1445(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1446(.a(s_128), .O(gate215inter3));
  inv1  gate1447(.a(s_129), .O(gate215inter4));
  nand2 gate1448(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1449(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1450(.a(G607), .O(gate215inter7));
  inv1  gate1451(.a(G675), .O(gate215inter8));
  nand2 gate1452(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1453(.a(s_129), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1454(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1455(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1456(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2367(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2368(.a(gate218inter0), .b(s_260), .O(gate218inter1));
  and2  gate2369(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2370(.a(s_260), .O(gate218inter3));
  inv1  gate2371(.a(s_261), .O(gate218inter4));
  nand2 gate2372(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2373(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2374(.a(G627), .O(gate218inter7));
  inv1  gate2375(.a(G678), .O(gate218inter8));
  nand2 gate2376(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2377(.a(s_261), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2378(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2379(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2380(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate771(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate772(.a(gate220inter0), .b(s_32), .O(gate220inter1));
  and2  gate773(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate774(.a(s_32), .O(gate220inter3));
  inv1  gate775(.a(s_33), .O(gate220inter4));
  nand2 gate776(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate777(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate778(.a(G637), .O(gate220inter7));
  inv1  gate779(.a(G681), .O(gate220inter8));
  nand2 gate780(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate781(.a(s_33), .b(gate220inter3), .O(gate220inter10));
  nor2  gate782(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate783(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate784(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1765(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1766(.a(gate223inter0), .b(s_174), .O(gate223inter1));
  and2  gate1767(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1768(.a(s_174), .O(gate223inter3));
  inv1  gate1769(.a(s_175), .O(gate223inter4));
  nand2 gate1770(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1771(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1772(.a(G627), .O(gate223inter7));
  inv1  gate1773(.a(G687), .O(gate223inter8));
  nand2 gate1774(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1775(.a(s_175), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1776(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1777(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1778(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate841(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate842(.a(gate224inter0), .b(s_42), .O(gate224inter1));
  and2  gate843(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate844(.a(s_42), .O(gate224inter3));
  inv1  gate845(.a(s_43), .O(gate224inter4));
  nand2 gate846(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate847(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate848(.a(G637), .O(gate224inter7));
  inv1  gate849(.a(G687), .O(gate224inter8));
  nand2 gate850(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate851(.a(s_43), .b(gate224inter3), .O(gate224inter10));
  nor2  gate852(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate853(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate854(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate2563(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate2564(.a(gate226inter0), .b(s_288), .O(gate226inter1));
  and2  gate2565(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate2566(.a(s_288), .O(gate226inter3));
  inv1  gate2567(.a(s_289), .O(gate226inter4));
  nand2 gate2568(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate2569(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate2570(.a(G692), .O(gate226inter7));
  inv1  gate2571(.a(G693), .O(gate226inter8));
  nand2 gate2572(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate2573(.a(s_289), .b(gate226inter3), .O(gate226inter10));
  nor2  gate2574(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate2575(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate2576(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2787(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2788(.a(gate230inter0), .b(s_320), .O(gate230inter1));
  and2  gate2789(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2790(.a(s_320), .O(gate230inter3));
  inv1  gate2791(.a(s_321), .O(gate230inter4));
  nand2 gate2792(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2793(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2794(.a(G700), .O(gate230inter7));
  inv1  gate2795(.a(G701), .O(gate230inter8));
  nand2 gate2796(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2797(.a(s_321), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2798(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2799(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2800(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2325(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2326(.a(gate232inter0), .b(s_254), .O(gate232inter1));
  and2  gate2327(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2328(.a(s_254), .O(gate232inter3));
  inv1  gate2329(.a(s_255), .O(gate232inter4));
  nand2 gate2330(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2331(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2332(.a(G704), .O(gate232inter7));
  inv1  gate2333(.a(G705), .O(gate232inter8));
  nand2 gate2334(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2335(.a(s_255), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2336(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2337(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2338(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1387(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1388(.a(gate236inter0), .b(s_120), .O(gate236inter1));
  and2  gate1389(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1390(.a(s_120), .O(gate236inter3));
  inv1  gate1391(.a(s_121), .O(gate236inter4));
  nand2 gate1392(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1393(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1394(.a(G251), .O(gate236inter7));
  inv1  gate1395(.a(G727), .O(gate236inter8));
  nand2 gate1396(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1397(.a(s_121), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1398(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1399(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1400(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1219(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1220(.a(gate238inter0), .b(s_96), .O(gate238inter1));
  and2  gate1221(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1222(.a(s_96), .O(gate238inter3));
  inv1  gate1223(.a(s_97), .O(gate238inter4));
  nand2 gate1224(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1225(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1226(.a(G257), .O(gate238inter7));
  inv1  gate1227(.a(G709), .O(gate238inter8));
  nand2 gate1228(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1229(.a(s_97), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1230(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1231(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1232(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate953(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate954(.a(gate243inter0), .b(s_58), .O(gate243inter1));
  and2  gate955(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate956(.a(s_58), .O(gate243inter3));
  inv1  gate957(.a(s_59), .O(gate243inter4));
  nand2 gate958(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate959(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate960(.a(G245), .O(gate243inter7));
  inv1  gate961(.a(G733), .O(gate243inter8));
  nand2 gate962(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate963(.a(s_59), .b(gate243inter3), .O(gate243inter10));
  nor2  gate964(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate965(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate966(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1345(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1346(.a(gate244inter0), .b(s_114), .O(gate244inter1));
  and2  gate1347(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1348(.a(s_114), .O(gate244inter3));
  inv1  gate1349(.a(s_115), .O(gate244inter4));
  nand2 gate1350(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1351(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1352(.a(G721), .O(gate244inter7));
  inv1  gate1353(.a(G733), .O(gate244inter8));
  nand2 gate1354(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1355(.a(s_115), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1356(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1357(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1358(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate2115(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2116(.a(gate245inter0), .b(s_224), .O(gate245inter1));
  and2  gate2117(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2118(.a(s_224), .O(gate245inter3));
  inv1  gate2119(.a(s_225), .O(gate245inter4));
  nand2 gate2120(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2121(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2122(.a(G248), .O(gate245inter7));
  inv1  gate2123(.a(G736), .O(gate245inter8));
  nand2 gate2124(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2125(.a(s_225), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2126(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2127(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2128(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1933(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1934(.a(gate248inter0), .b(s_198), .O(gate248inter1));
  and2  gate1935(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1936(.a(s_198), .O(gate248inter3));
  inv1  gate1937(.a(s_199), .O(gate248inter4));
  nand2 gate1938(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1939(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1940(.a(G727), .O(gate248inter7));
  inv1  gate1941(.a(G739), .O(gate248inter8));
  nand2 gate1942(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1943(.a(s_199), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1944(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1945(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1946(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2465(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2466(.a(gate249inter0), .b(s_274), .O(gate249inter1));
  and2  gate2467(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2468(.a(s_274), .O(gate249inter3));
  inv1  gate2469(.a(s_275), .O(gate249inter4));
  nand2 gate2470(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2471(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2472(.a(G254), .O(gate249inter7));
  inv1  gate2473(.a(G742), .O(gate249inter8));
  nand2 gate2474(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2475(.a(s_275), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2476(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2477(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2478(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2885(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2886(.a(gate250inter0), .b(s_334), .O(gate250inter1));
  and2  gate2887(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2888(.a(s_334), .O(gate250inter3));
  inv1  gate2889(.a(s_335), .O(gate250inter4));
  nand2 gate2890(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2891(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2892(.a(G706), .O(gate250inter7));
  inv1  gate2893(.a(G742), .O(gate250inter8));
  nand2 gate2894(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2895(.a(s_335), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2896(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2897(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2898(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2395(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2396(.a(gate252inter0), .b(s_264), .O(gate252inter1));
  and2  gate2397(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2398(.a(s_264), .O(gate252inter3));
  inv1  gate2399(.a(s_265), .O(gate252inter4));
  nand2 gate2400(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2401(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2402(.a(G709), .O(gate252inter7));
  inv1  gate2403(.a(G745), .O(gate252inter8));
  nand2 gate2404(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2405(.a(s_265), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2406(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2407(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2408(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2577(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2578(.a(gate257inter0), .b(s_290), .O(gate257inter1));
  and2  gate2579(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2580(.a(s_290), .O(gate257inter3));
  inv1  gate2581(.a(s_291), .O(gate257inter4));
  nand2 gate2582(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2583(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2584(.a(G754), .O(gate257inter7));
  inv1  gate2585(.a(G755), .O(gate257inter8));
  nand2 gate2586(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2587(.a(s_291), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2588(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2589(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2590(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate617(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate618(.a(gate259inter0), .b(s_10), .O(gate259inter1));
  and2  gate619(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate620(.a(s_10), .O(gate259inter3));
  inv1  gate621(.a(s_11), .O(gate259inter4));
  nand2 gate622(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate623(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate624(.a(G758), .O(gate259inter7));
  inv1  gate625(.a(G759), .O(gate259inter8));
  nand2 gate626(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate627(.a(s_11), .b(gate259inter3), .O(gate259inter10));
  nor2  gate628(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate629(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate630(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2549(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2550(.a(gate261inter0), .b(s_286), .O(gate261inter1));
  and2  gate2551(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2552(.a(s_286), .O(gate261inter3));
  inv1  gate2553(.a(s_287), .O(gate261inter4));
  nand2 gate2554(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2555(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2556(.a(G762), .O(gate261inter7));
  inv1  gate2557(.a(G763), .O(gate261inter8));
  nand2 gate2558(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2559(.a(s_287), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2560(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2561(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2562(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2143(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2144(.a(gate264inter0), .b(s_228), .O(gate264inter1));
  and2  gate2145(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2146(.a(s_228), .O(gate264inter3));
  inv1  gate2147(.a(s_229), .O(gate264inter4));
  nand2 gate2148(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2149(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2150(.a(G768), .O(gate264inter7));
  inv1  gate2151(.a(G769), .O(gate264inter8));
  nand2 gate2152(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2153(.a(s_229), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2154(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2155(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2156(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1149(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1150(.a(gate267inter0), .b(s_86), .O(gate267inter1));
  and2  gate1151(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1152(.a(s_86), .O(gate267inter3));
  inv1  gate1153(.a(s_87), .O(gate267inter4));
  nand2 gate1154(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1155(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1156(.a(G648), .O(gate267inter7));
  inv1  gate1157(.a(G776), .O(gate267inter8));
  nand2 gate1158(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1159(.a(s_87), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1160(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1161(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1162(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate813(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate814(.a(gate269inter0), .b(s_38), .O(gate269inter1));
  and2  gate815(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate816(.a(s_38), .O(gate269inter3));
  inv1  gate817(.a(s_39), .O(gate269inter4));
  nand2 gate818(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate819(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate820(.a(G654), .O(gate269inter7));
  inv1  gate821(.a(G782), .O(gate269inter8));
  nand2 gate822(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate823(.a(s_39), .b(gate269inter3), .O(gate269inter10));
  nor2  gate824(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate825(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate826(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1121(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1122(.a(gate272inter0), .b(s_82), .O(gate272inter1));
  and2  gate1123(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1124(.a(s_82), .O(gate272inter3));
  inv1  gate1125(.a(s_83), .O(gate272inter4));
  nand2 gate1126(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1127(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1128(.a(G663), .O(gate272inter7));
  inv1  gate1129(.a(G791), .O(gate272inter8));
  nand2 gate1130(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1131(.a(s_83), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1132(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1133(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1134(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2689(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2690(.a(gate274inter0), .b(s_306), .O(gate274inter1));
  and2  gate2691(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2692(.a(s_306), .O(gate274inter3));
  inv1  gate2693(.a(s_307), .O(gate274inter4));
  nand2 gate2694(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2695(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2696(.a(G770), .O(gate274inter7));
  inv1  gate2697(.a(G794), .O(gate274inter8));
  nand2 gate2698(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2699(.a(s_307), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2700(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2701(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2702(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1779(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1780(.a(gate275inter0), .b(s_176), .O(gate275inter1));
  and2  gate1781(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1782(.a(s_176), .O(gate275inter3));
  inv1  gate1783(.a(s_177), .O(gate275inter4));
  nand2 gate1784(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1785(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1786(.a(G645), .O(gate275inter7));
  inv1  gate1787(.a(G797), .O(gate275inter8));
  nand2 gate1788(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1789(.a(s_177), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1790(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1791(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1792(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1359(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1360(.a(gate276inter0), .b(s_116), .O(gate276inter1));
  and2  gate1361(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1362(.a(s_116), .O(gate276inter3));
  inv1  gate1363(.a(s_117), .O(gate276inter4));
  nand2 gate1364(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1365(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1366(.a(G773), .O(gate276inter7));
  inv1  gate1367(.a(G797), .O(gate276inter8));
  nand2 gate1368(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1369(.a(s_117), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1370(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1371(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1372(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1331(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1332(.a(gate280inter0), .b(s_112), .O(gate280inter1));
  and2  gate1333(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1334(.a(s_112), .O(gate280inter3));
  inv1  gate1335(.a(s_113), .O(gate280inter4));
  nand2 gate1336(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1337(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1338(.a(G779), .O(gate280inter7));
  inv1  gate1339(.a(G803), .O(gate280inter8));
  nand2 gate1340(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1341(.a(s_113), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1342(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1343(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1344(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1667(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1668(.a(gate281inter0), .b(s_160), .O(gate281inter1));
  and2  gate1669(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1670(.a(s_160), .O(gate281inter3));
  inv1  gate1671(.a(s_161), .O(gate281inter4));
  nand2 gate1672(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1673(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1674(.a(G654), .O(gate281inter7));
  inv1  gate1675(.a(G806), .O(gate281inter8));
  nand2 gate1676(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1677(.a(s_161), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1678(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1679(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1680(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1989(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1990(.a(gate288inter0), .b(s_206), .O(gate288inter1));
  and2  gate1991(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1992(.a(s_206), .O(gate288inter3));
  inv1  gate1993(.a(s_207), .O(gate288inter4));
  nand2 gate1994(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1995(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1996(.a(G791), .O(gate288inter7));
  inv1  gate1997(.a(G815), .O(gate288inter8));
  nand2 gate1998(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1999(.a(s_207), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2000(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2001(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2002(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1863(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1864(.a(gate290inter0), .b(s_188), .O(gate290inter1));
  and2  gate1865(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1866(.a(s_188), .O(gate290inter3));
  inv1  gate1867(.a(s_189), .O(gate290inter4));
  nand2 gate1868(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1869(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1870(.a(G820), .O(gate290inter7));
  inv1  gate1871(.a(G821), .O(gate290inter8));
  nand2 gate1872(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1873(.a(s_189), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1874(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1875(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1876(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2801(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2802(.a(gate291inter0), .b(s_322), .O(gate291inter1));
  and2  gate2803(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2804(.a(s_322), .O(gate291inter3));
  inv1  gate2805(.a(s_323), .O(gate291inter4));
  nand2 gate2806(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2807(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2808(.a(G822), .O(gate291inter7));
  inv1  gate2809(.a(G823), .O(gate291inter8));
  nand2 gate2810(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2811(.a(s_323), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2812(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2813(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2814(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1583(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1584(.a(gate292inter0), .b(s_148), .O(gate292inter1));
  and2  gate1585(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1586(.a(s_148), .O(gate292inter3));
  inv1  gate1587(.a(s_149), .O(gate292inter4));
  nand2 gate1588(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1589(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1590(.a(G824), .O(gate292inter7));
  inv1  gate1591(.a(G825), .O(gate292inter8));
  nand2 gate1592(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1593(.a(s_149), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1594(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1595(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1596(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2297(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2298(.a(gate387inter0), .b(s_250), .O(gate387inter1));
  and2  gate2299(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2300(.a(s_250), .O(gate387inter3));
  inv1  gate2301(.a(s_251), .O(gate387inter4));
  nand2 gate2302(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2303(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2304(.a(G1), .O(gate387inter7));
  inv1  gate2305(.a(G1036), .O(gate387inter8));
  nand2 gate2306(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2307(.a(s_251), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2308(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2309(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2310(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate799(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate800(.a(gate388inter0), .b(s_36), .O(gate388inter1));
  and2  gate801(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate802(.a(s_36), .O(gate388inter3));
  inv1  gate803(.a(s_37), .O(gate388inter4));
  nand2 gate804(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate805(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate806(.a(G2), .O(gate388inter7));
  inv1  gate807(.a(G1039), .O(gate388inter8));
  nand2 gate808(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate809(.a(s_37), .b(gate388inter3), .O(gate388inter10));
  nor2  gate810(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate811(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate812(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2843(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2844(.a(gate392inter0), .b(s_328), .O(gate392inter1));
  and2  gate2845(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2846(.a(s_328), .O(gate392inter3));
  inv1  gate2847(.a(s_329), .O(gate392inter4));
  nand2 gate2848(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2849(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2850(.a(G6), .O(gate392inter7));
  inv1  gate2851(.a(G1051), .O(gate392inter8));
  nand2 gate2852(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2853(.a(s_329), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2854(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2855(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2856(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1821(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1822(.a(gate393inter0), .b(s_182), .O(gate393inter1));
  and2  gate1823(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1824(.a(s_182), .O(gate393inter3));
  inv1  gate1825(.a(s_183), .O(gate393inter4));
  nand2 gate1826(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1827(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1828(.a(G7), .O(gate393inter7));
  inv1  gate1829(.a(G1054), .O(gate393inter8));
  nand2 gate1830(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1831(.a(s_183), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1832(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1833(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1834(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2507(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2508(.a(gate396inter0), .b(s_280), .O(gate396inter1));
  and2  gate2509(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2510(.a(s_280), .O(gate396inter3));
  inv1  gate2511(.a(s_281), .O(gate396inter4));
  nand2 gate2512(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2513(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2514(.a(G10), .O(gate396inter7));
  inv1  gate2515(.a(G1063), .O(gate396inter8));
  nand2 gate2516(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2517(.a(s_281), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2518(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2519(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2520(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate659(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate660(.a(gate398inter0), .b(s_16), .O(gate398inter1));
  and2  gate661(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate662(.a(s_16), .O(gate398inter3));
  inv1  gate663(.a(s_17), .O(gate398inter4));
  nand2 gate664(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate665(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate666(.a(G12), .O(gate398inter7));
  inv1  gate667(.a(G1069), .O(gate398inter8));
  nand2 gate668(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate669(.a(s_17), .b(gate398inter3), .O(gate398inter10));
  nor2  gate670(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate671(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate672(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate2409(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2410(.a(gate399inter0), .b(s_266), .O(gate399inter1));
  and2  gate2411(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2412(.a(s_266), .O(gate399inter3));
  inv1  gate2413(.a(s_267), .O(gate399inter4));
  nand2 gate2414(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2415(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2416(.a(G13), .O(gate399inter7));
  inv1  gate2417(.a(G1072), .O(gate399inter8));
  nand2 gate2418(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2419(.a(s_267), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2420(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2421(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2422(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2255(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2256(.a(gate400inter0), .b(s_244), .O(gate400inter1));
  and2  gate2257(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2258(.a(s_244), .O(gate400inter3));
  inv1  gate2259(.a(s_245), .O(gate400inter4));
  nand2 gate2260(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2261(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2262(.a(G14), .O(gate400inter7));
  inv1  gate2263(.a(G1075), .O(gate400inter8));
  nand2 gate2264(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2265(.a(s_245), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2266(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2267(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2268(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2283(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2284(.a(gate406inter0), .b(s_248), .O(gate406inter1));
  and2  gate2285(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2286(.a(s_248), .O(gate406inter3));
  inv1  gate2287(.a(s_249), .O(gate406inter4));
  nand2 gate2288(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2289(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2290(.a(G20), .O(gate406inter7));
  inv1  gate2291(.a(G1093), .O(gate406inter8));
  nand2 gate2292(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2293(.a(s_249), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2294(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2295(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2296(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate701(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate702(.a(gate407inter0), .b(s_22), .O(gate407inter1));
  and2  gate703(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate704(.a(s_22), .O(gate407inter3));
  inv1  gate705(.a(s_23), .O(gate407inter4));
  nand2 gate706(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate707(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate708(.a(G21), .O(gate407inter7));
  inv1  gate709(.a(G1096), .O(gate407inter8));
  nand2 gate710(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate711(.a(s_23), .b(gate407inter3), .O(gate407inter10));
  nor2  gate712(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate713(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate714(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate827(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate828(.a(gate410inter0), .b(s_40), .O(gate410inter1));
  and2  gate829(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate830(.a(s_40), .O(gate410inter3));
  inv1  gate831(.a(s_41), .O(gate410inter4));
  nand2 gate832(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate833(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate834(.a(G24), .O(gate410inter7));
  inv1  gate835(.a(G1105), .O(gate410inter8));
  nand2 gate836(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate837(.a(s_41), .b(gate410inter3), .O(gate410inter10));
  nor2  gate838(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate839(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate840(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1275(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1276(.a(gate412inter0), .b(s_104), .O(gate412inter1));
  and2  gate1277(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1278(.a(s_104), .O(gate412inter3));
  inv1  gate1279(.a(s_105), .O(gate412inter4));
  nand2 gate1280(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1281(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1282(.a(G26), .O(gate412inter7));
  inv1  gate1283(.a(G1111), .O(gate412inter8));
  nand2 gate1284(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1285(.a(s_105), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1286(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1287(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1288(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate785(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate786(.a(gate419inter0), .b(s_34), .O(gate419inter1));
  and2  gate787(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate788(.a(s_34), .O(gate419inter3));
  inv1  gate789(.a(s_35), .O(gate419inter4));
  nand2 gate790(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate791(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate792(.a(G1), .O(gate419inter7));
  inv1  gate793(.a(G1132), .O(gate419inter8));
  nand2 gate794(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate795(.a(s_35), .b(gate419inter3), .O(gate419inter10));
  nor2  gate796(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate797(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate798(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1723(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1724(.a(gate421inter0), .b(s_168), .O(gate421inter1));
  and2  gate1725(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1726(.a(s_168), .O(gate421inter3));
  inv1  gate1727(.a(s_169), .O(gate421inter4));
  nand2 gate1728(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1729(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1730(.a(G2), .O(gate421inter7));
  inv1  gate1731(.a(G1135), .O(gate421inter8));
  nand2 gate1732(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1733(.a(s_169), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1734(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1735(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1736(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1681(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1682(.a(gate422inter0), .b(s_162), .O(gate422inter1));
  and2  gate1683(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1684(.a(s_162), .O(gate422inter3));
  inv1  gate1685(.a(s_163), .O(gate422inter4));
  nand2 gate1686(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1687(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1688(.a(G1039), .O(gate422inter7));
  inv1  gate1689(.a(G1135), .O(gate422inter8));
  nand2 gate1690(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1691(.a(s_163), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1692(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1693(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1694(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1905(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1906(.a(gate423inter0), .b(s_194), .O(gate423inter1));
  and2  gate1907(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1908(.a(s_194), .O(gate423inter3));
  inv1  gate1909(.a(s_195), .O(gate423inter4));
  nand2 gate1910(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1911(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1912(.a(G3), .O(gate423inter7));
  inv1  gate1913(.a(G1138), .O(gate423inter8));
  nand2 gate1914(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1915(.a(s_195), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1916(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1917(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1918(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2129(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2130(.a(gate427inter0), .b(s_226), .O(gate427inter1));
  and2  gate2131(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2132(.a(s_226), .O(gate427inter3));
  inv1  gate2133(.a(s_227), .O(gate427inter4));
  nand2 gate2134(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2135(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2136(.a(G5), .O(gate427inter7));
  inv1  gate2137(.a(G1144), .O(gate427inter8));
  nand2 gate2138(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2139(.a(s_227), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2140(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2141(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2142(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1835(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1836(.a(gate430inter0), .b(s_184), .O(gate430inter1));
  and2  gate1837(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1838(.a(s_184), .O(gate430inter3));
  inv1  gate1839(.a(s_185), .O(gate430inter4));
  nand2 gate1840(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1841(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1842(.a(G1051), .O(gate430inter7));
  inv1  gate1843(.a(G1147), .O(gate430inter8));
  nand2 gate1844(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1845(.a(s_185), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1846(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1847(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1848(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2381(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2382(.a(gate432inter0), .b(s_262), .O(gate432inter1));
  and2  gate2383(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2384(.a(s_262), .O(gate432inter3));
  inv1  gate2385(.a(s_263), .O(gate432inter4));
  nand2 gate2386(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2387(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2388(.a(G1054), .O(gate432inter7));
  inv1  gate2389(.a(G1150), .O(gate432inter8));
  nand2 gate2390(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2391(.a(s_263), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2392(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2393(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2394(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate2675(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2676(.a(gate437inter0), .b(s_304), .O(gate437inter1));
  and2  gate2677(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2678(.a(s_304), .O(gate437inter3));
  inv1  gate2679(.a(s_305), .O(gate437inter4));
  nand2 gate2680(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2681(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2682(.a(G10), .O(gate437inter7));
  inv1  gate2683(.a(G1159), .O(gate437inter8));
  nand2 gate2684(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2685(.a(s_305), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2686(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2687(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2688(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate757(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate758(.a(gate439inter0), .b(s_30), .O(gate439inter1));
  and2  gate759(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate760(.a(s_30), .O(gate439inter3));
  inv1  gate761(.a(s_31), .O(gate439inter4));
  nand2 gate762(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate763(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate764(.a(G11), .O(gate439inter7));
  inv1  gate765(.a(G1162), .O(gate439inter8));
  nand2 gate766(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate767(.a(s_31), .b(gate439inter3), .O(gate439inter10));
  nor2  gate768(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate769(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate770(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1499(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1500(.a(gate440inter0), .b(s_136), .O(gate440inter1));
  and2  gate1501(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1502(.a(s_136), .O(gate440inter3));
  inv1  gate1503(.a(s_137), .O(gate440inter4));
  nand2 gate1504(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1505(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1506(.a(G1066), .O(gate440inter7));
  inv1  gate1507(.a(G1162), .O(gate440inter8));
  nand2 gate1508(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1509(.a(s_137), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1510(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1511(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1512(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate673(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate674(.a(gate446inter0), .b(s_18), .O(gate446inter1));
  and2  gate675(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate676(.a(s_18), .O(gate446inter3));
  inv1  gate677(.a(s_19), .O(gate446inter4));
  nand2 gate678(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate679(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate680(.a(G1075), .O(gate446inter7));
  inv1  gate681(.a(G1171), .O(gate446inter8));
  nand2 gate682(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate683(.a(s_19), .b(gate446inter3), .O(gate446inter10));
  nor2  gate684(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate685(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate686(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1737(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1738(.a(gate447inter0), .b(s_170), .O(gate447inter1));
  and2  gate1739(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1740(.a(s_170), .O(gate447inter3));
  inv1  gate1741(.a(s_171), .O(gate447inter4));
  nand2 gate1742(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1743(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1744(.a(G15), .O(gate447inter7));
  inv1  gate1745(.a(G1174), .O(gate447inter8));
  nand2 gate1746(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1747(.a(s_171), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1748(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1749(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1750(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1107(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1108(.a(gate449inter0), .b(s_80), .O(gate449inter1));
  and2  gate1109(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1110(.a(s_80), .O(gate449inter3));
  inv1  gate1111(.a(s_81), .O(gate449inter4));
  nand2 gate1112(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1113(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1114(.a(G16), .O(gate449inter7));
  inv1  gate1115(.a(G1177), .O(gate449inter8));
  nand2 gate1116(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1117(.a(s_81), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1118(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1119(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1120(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate743(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate744(.a(gate450inter0), .b(s_28), .O(gate450inter1));
  and2  gate745(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate746(.a(s_28), .O(gate450inter3));
  inv1  gate747(.a(s_29), .O(gate450inter4));
  nand2 gate748(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate749(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate750(.a(G1081), .O(gate450inter7));
  inv1  gate751(.a(G1177), .O(gate450inter8));
  nand2 gate752(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate753(.a(s_29), .b(gate450inter3), .O(gate450inter10));
  nor2  gate754(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate755(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate756(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2591(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2592(.a(gate456inter0), .b(s_292), .O(gate456inter1));
  and2  gate2593(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2594(.a(s_292), .O(gate456inter3));
  inv1  gate2595(.a(s_293), .O(gate456inter4));
  nand2 gate2596(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2597(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2598(.a(G1090), .O(gate456inter7));
  inv1  gate2599(.a(G1186), .O(gate456inter8));
  nand2 gate2600(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2601(.a(s_293), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2602(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2603(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2604(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate2171(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2172(.a(gate457inter0), .b(s_232), .O(gate457inter1));
  and2  gate2173(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2174(.a(s_232), .O(gate457inter3));
  inv1  gate2175(.a(s_233), .O(gate457inter4));
  nand2 gate2176(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2177(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2178(.a(G20), .O(gate457inter7));
  inv1  gate2179(.a(G1189), .O(gate457inter8));
  nand2 gate2180(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2181(.a(s_233), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2182(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2183(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2184(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1975(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1976(.a(gate458inter0), .b(s_204), .O(gate458inter1));
  and2  gate1977(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1978(.a(s_204), .O(gate458inter3));
  inv1  gate1979(.a(s_205), .O(gate458inter4));
  nand2 gate1980(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1981(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1982(.a(G1093), .O(gate458inter7));
  inv1  gate1983(.a(G1189), .O(gate458inter8));
  nand2 gate1984(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1985(.a(s_205), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1986(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1987(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1988(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate2213(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2214(.a(gate459inter0), .b(s_238), .O(gate459inter1));
  and2  gate2215(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2216(.a(s_238), .O(gate459inter3));
  inv1  gate2217(.a(s_239), .O(gate459inter4));
  nand2 gate2218(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2219(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2220(.a(G21), .O(gate459inter7));
  inv1  gate2221(.a(G1192), .O(gate459inter8));
  nand2 gate2222(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2223(.a(s_239), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2224(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2225(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2226(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2857(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2858(.a(gate461inter0), .b(s_330), .O(gate461inter1));
  and2  gate2859(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2860(.a(s_330), .O(gate461inter3));
  inv1  gate2861(.a(s_331), .O(gate461inter4));
  nand2 gate2862(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2863(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2864(.a(G22), .O(gate461inter7));
  inv1  gate2865(.a(G1195), .O(gate461inter8));
  nand2 gate2866(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2867(.a(s_331), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2868(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2869(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2870(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2003(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2004(.a(gate462inter0), .b(s_208), .O(gate462inter1));
  and2  gate2005(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2006(.a(s_208), .O(gate462inter3));
  inv1  gate2007(.a(s_209), .O(gate462inter4));
  nand2 gate2008(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2009(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2010(.a(G1099), .O(gate462inter7));
  inv1  gate2011(.a(G1195), .O(gate462inter8));
  nand2 gate2012(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2013(.a(s_209), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2014(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2015(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2016(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1807(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1808(.a(gate467inter0), .b(s_180), .O(gate467inter1));
  and2  gate1809(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1810(.a(s_180), .O(gate467inter3));
  inv1  gate1811(.a(s_181), .O(gate467inter4));
  nand2 gate1812(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1813(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1814(.a(G25), .O(gate467inter7));
  inv1  gate1815(.a(G1204), .O(gate467inter8));
  nand2 gate1816(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1817(.a(s_181), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1818(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1819(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1820(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1653(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1654(.a(gate468inter0), .b(s_158), .O(gate468inter1));
  and2  gate1655(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1656(.a(s_158), .O(gate468inter3));
  inv1  gate1657(.a(s_159), .O(gate468inter4));
  nand2 gate1658(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1659(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1660(.a(G1108), .O(gate468inter7));
  inv1  gate1661(.a(G1204), .O(gate468inter8));
  nand2 gate1662(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1663(.a(s_159), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1664(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1665(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1666(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1023(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1024(.a(gate470inter0), .b(s_68), .O(gate470inter1));
  and2  gate1025(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1026(.a(s_68), .O(gate470inter3));
  inv1  gate1027(.a(s_69), .O(gate470inter4));
  nand2 gate1028(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1029(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1030(.a(G1111), .O(gate470inter7));
  inv1  gate1031(.a(G1207), .O(gate470inter8));
  nand2 gate1032(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1033(.a(s_69), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1034(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1035(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1036(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1877(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1878(.a(gate471inter0), .b(s_190), .O(gate471inter1));
  and2  gate1879(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1880(.a(s_190), .O(gate471inter3));
  inv1  gate1881(.a(s_191), .O(gate471inter4));
  nand2 gate1882(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1883(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1884(.a(G27), .O(gate471inter7));
  inv1  gate1885(.a(G1210), .O(gate471inter8));
  nand2 gate1886(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1887(.a(s_191), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1888(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1889(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1890(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2493(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2494(.a(gate472inter0), .b(s_278), .O(gate472inter1));
  and2  gate2495(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2496(.a(s_278), .O(gate472inter3));
  inv1  gate2497(.a(s_279), .O(gate472inter4));
  nand2 gate2498(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2499(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2500(.a(G1114), .O(gate472inter7));
  inv1  gate2501(.a(G1210), .O(gate472inter8));
  nand2 gate2502(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2503(.a(s_279), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2504(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2505(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2506(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2101(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2102(.a(gate477inter0), .b(s_222), .O(gate477inter1));
  and2  gate2103(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2104(.a(s_222), .O(gate477inter3));
  inv1  gate2105(.a(s_223), .O(gate477inter4));
  nand2 gate2106(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2107(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2108(.a(G30), .O(gate477inter7));
  inv1  gate2109(.a(G1219), .O(gate477inter8));
  nand2 gate2110(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2111(.a(s_223), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2112(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2113(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2114(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1611(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1612(.a(gate478inter0), .b(s_152), .O(gate478inter1));
  and2  gate1613(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1614(.a(s_152), .O(gate478inter3));
  inv1  gate1615(.a(s_153), .O(gate478inter4));
  nand2 gate1616(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1617(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1618(.a(G1123), .O(gate478inter7));
  inv1  gate1619(.a(G1219), .O(gate478inter8));
  nand2 gate1620(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1621(.a(s_153), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1622(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1623(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1624(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate2815(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2816(.a(gate481inter0), .b(s_324), .O(gate481inter1));
  and2  gate2817(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2818(.a(s_324), .O(gate481inter3));
  inv1  gate2819(.a(s_325), .O(gate481inter4));
  nand2 gate2820(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2821(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2822(.a(G32), .O(gate481inter7));
  inv1  gate2823(.a(G1225), .O(gate481inter8));
  nand2 gate2824(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2825(.a(s_325), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2826(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2827(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2828(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate2703(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2704(.a(gate482inter0), .b(s_308), .O(gate482inter1));
  and2  gate2705(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2706(.a(s_308), .O(gate482inter3));
  inv1  gate2707(.a(s_309), .O(gate482inter4));
  nand2 gate2708(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2709(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2710(.a(G1129), .O(gate482inter7));
  inv1  gate2711(.a(G1225), .O(gate482inter8));
  nand2 gate2712(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2713(.a(s_309), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2714(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2715(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2716(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2241(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2242(.a(gate486inter0), .b(s_242), .O(gate486inter1));
  and2  gate2243(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2244(.a(s_242), .O(gate486inter3));
  inv1  gate2245(.a(s_243), .O(gate486inter4));
  nand2 gate2246(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2247(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2248(.a(G1234), .O(gate486inter7));
  inv1  gate2249(.a(G1235), .O(gate486inter8));
  nand2 gate2250(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2251(.a(s_243), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2252(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2253(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2254(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1919(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1920(.a(gate493inter0), .b(s_196), .O(gate493inter1));
  and2  gate1921(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1922(.a(s_196), .O(gate493inter3));
  inv1  gate1923(.a(s_197), .O(gate493inter4));
  nand2 gate1924(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1925(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1926(.a(G1248), .O(gate493inter7));
  inv1  gate1927(.a(G1249), .O(gate493inter8));
  nand2 gate1928(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1929(.a(s_197), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1930(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1931(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1932(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1429(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1430(.a(gate494inter0), .b(s_126), .O(gate494inter1));
  and2  gate1431(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1432(.a(s_126), .O(gate494inter3));
  inv1  gate1433(.a(s_127), .O(gate494inter4));
  nand2 gate1434(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1435(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1436(.a(G1250), .O(gate494inter7));
  inv1  gate1437(.a(G1251), .O(gate494inter8));
  nand2 gate1438(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1439(.a(s_127), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1440(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1441(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1442(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate589(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate590(.a(gate496inter0), .b(s_6), .O(gate496inter1));
  and2  gate591(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate592(.a(s_6), .O(gate496inter3));
  inv1  gate593(.a(s_7), .O(gate496inter4));
  nand2 gate594(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate595(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate596(.a(G1254), .O(gate496inter7));
  inv1  gate597(.a(G1255), .O(gate496inter8));
  nand2 gate598(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate599(.a(s_7), .b(gate496inter3), .O(gate496inter10));
  nor2  gate600(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate601(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate602(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1261(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1262(.a(gate502inter0), .b(s_102), .O(gate502inter1));
  and2  gate1263(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1264(.a(s_102), .O(gate502inter3));
  inv1  gate1265(.a(s_103), .O(gate502inter4));
  nand2 gate1266(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1267(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1268(.a(G1266), .O(gate502inter7));
  inv1  gate1269(.a(G1267), .O(gate502inter8));
  nand2 gate1270(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1271(.a(s_103), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1272(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1273(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1274(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2269(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2270(.a(gate503inter0), .b(s_246), .O(gate503inter1));
  and2  gate2271(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2272(.a(s_246), .O(gate503inter3));
  inv1  gate2273(.a(s_247), .O(gate503inter4));
  nand2 gate2274(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2275(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2276(.a(G1268), .O(gate503inter7));
  inv1  gate2277(.a(G1269), .O(gate503inter8));
  nand2 gate2278(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2279(.a(s_247), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2280(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2281(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2282(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1527(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1528(.a(gate505inter0), .b(s_140), .O(gate505inter1));
  and2  gate1529(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1530(.a(s_140), .O(gate505inter3));
  inv1  gate1531(.a(s_141), .O(gate505inter4));
  nand2 gate1532(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1533(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1534(.a(G1272), .O(gate505inter7));
  inv1  gate1535(.a(G1273), .O(gate505inter8));
  nand2 gate1536(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1537(.a(s_141), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1538(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1539(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1540(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate2745(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2746(.a(gate506inter0), .b(s_314), .O(gate506inter1));
  and2  gate2747(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2748(.a(s_314), .O(gate506inter3));
  inv1  gate2749(.a(s_315), .O(gate506inter4));
  nand2 gate2750(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2751(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2752(.a(G1274), .O(gate506inter7));
  inv1  gate2753(.a(G1275), .O(gate506inter8));
  nand2 gate2754(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2755(.a(s_315), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2756(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2757(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2758(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1541(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1542(.a(gate508inter0), .b(s_142), .O(gate508inter1));
  and2  gate1543(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1544(.a(s_142), .O(gate508inter3));
  inv1  gate1545(.a(s_143), .O(gate508inter4));
  nand2 gate1546(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1547(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1548(.a(G1278), .O(gate508inter7));
  inv1  gate1549(.a(G1279), .O(gate508inter8));
  nand2 gate1550(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1551(.a(s_143), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1552(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1553(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1554(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate547(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate548(.a(gate509inter0), .b(s_0), .O(gate509inter1));
  and2  gate549(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate550(.a(s_0), .O(gate509inter3));
  inv1  gate551(.a(s_1), .O(gate509inter4));
  nand2 gate552(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate553(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate554(.a(G1280), .O(gate509inter7));
  inv1  gate555(.a(G1281), .O(gate509inter8));
  nand2 gate556(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate557(.a(s_1), .b(gate509inter3), .O(gate509inter10));
  nor2  gate558(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate559(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate560(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate855(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate856(.a(gate510inter0), .b(s_44), .O(gate510inter1));
  and2  gate857(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate858(.a(s_44), .O(gate510inter3));
  inv1  gate859(.a(s_45), .O(gate510inter4));
  nand2 gate860(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate861(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate862(.a(G1282), .O(gate510inter7));
  inv1  gate863(.a(G1283), .O(gate510inter8));
  nand2 gate864(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate865(.a(s_45), .b(gate510inter3), .O(gate510inter10));
  nor2  gate866(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate867(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate868(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1177(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1178(.a(gate511inter0), .b(s_90), .O(gate511inter1));
  and2  gate1179(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1180(.a(s_90), .O(gate511inter3));
  inv1  gate1181(.a(s_91), .O(gate511inter4));
  nand2 gate1182(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1183(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1184(.a(G1284), .O(gate511inter7));
  inv1  gate1185(.a(G1285), .O(gate511inter8));
  nand2 gate1186(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1187(.a(s_91), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1188(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1189(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1190(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate687(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate688(.a(gate513inter0), .b(s_20), .O(gate513inter1));
  and2  gate689(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate690(.a(s_20), .O(gate513inter3));
  inv1  gate691(.a(s_21), .O(gate513inter4));
  nand2 gate692(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate693(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate694(.a(G1288), .O(gate513inter7));
  inv1  gate695(.a(G1289), .O(gate513inter8));
  nand2 gate696(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate697(.a(s_21), .b(gate513inter3), .O(gate513inter10));
  nor2  gate698(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate699(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate700(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule