module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2465(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2466(.a(gate9inter0), .b(s_274), .O(gate9inter1));
  and2  gate2467(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2468(.a(s_274), .O(gate9inter3));
  inv1  gate2469(.a(s_275), .O(gate9inter4));
  nand2 gate2470(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2471(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2472(.a(G1), .O(gate9inter7));
  inv1  gate2473(.a(G2), .O(gate9inter8));
  nand2 gate2474(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2475(.a(s_275), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2476(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2477(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2478(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate659(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate660(.a(gate11inter0), .b(s_16), .O(gate11inter1));
  and2  gate661(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate662(.a(s_16), .O(gate11inter3));
  inv1  gate663(.a(s_17), .O(gate11inter4));
  nand2 gate664(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate665(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate666(.a(G5), .O(gate11inter7));
  inv1  gate667(.a(G6), .O(gate11inter8));
  nand2 gate668(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate669(.a(s_17), .b(gate11inter3), .O(gate11inter10));
  nor2  gate670(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate671(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate672(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2241(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2242(.a(gate15inter0), .b(s_242), .O(gate15inter1));
  and2  gate2243(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2244(.a(s_242), .O(gate15inter3));
  inv1  gate2245(.a(s_243), .O(gate15inter4));
  nand2 gate2246(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2247(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2248(.a(G13), .O(gate15inter7));
  inv1  gate2249(.a(G14), .O(gate15inter8));
  nand2 gate2250(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2251(.a(s_243), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2252(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2253(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2254(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1975(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1976(.a(gate16inter0), .b(s_204), .O(gate16inter1));
  and2  gate1977(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1978(.a(s_204), .O(gate16inter3));
  inv1  gate1979(.a(s_205), .O(gate16inter4));
  nand2 gate1980(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1981(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1982(.a(G15), .O(gate16inter7));
  inv1  gate1983(.a(G16), .O(gate16inter8));
  nand2 gate1984(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1985(.a(s_205), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1986(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1987(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1988(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2059(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2060(.a(gate17inter0), .b(s_216), .O(gate17inter1));
  and2  gate2061(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2062(.a(s_216), .O(gate17inter3));
  inv1  gate2063(.a(s_217), .O(gate17inter4));
  nand2 gate2064(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2065(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2066(.a(G17), .O(gate17inter7));
  inv1  gate2067(.a(G18), .O(gate17inter8));
  nand2 gate2068(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2069(.a(s_217), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2070(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2071(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2072(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate3179(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate3180(.a(gate21inter0), .b(s_376), .O(gate21inter1));
  and2  gate3181(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate3182(.a(s_376), .O(gate21inter3));
  inv1  gate3183(.a(s_377), .O(gate21inter4));
  nand2 gate3184(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate3185(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate3186(.a(G25), .O(gate21inter7));
  inv1  gate3187(.a(G26), .O(gate21inter8));
  nand2 gate3188(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate3189(.a(s_377), .b(gate21inter3), .O(gate21inter10));
  nor2  gate3190(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate3191(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate3192(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate617(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate618(.a(gate22inter0), .b(s_10), .O(gate22inter1));
  and2  gate619(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate620(.a(s_10), .O(gate22inter3));
  inv1  gate621(.a(s_11), .O(gate22inter4));
  nand2 gate622(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate623(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate624(.a(G27), .O(gate22inter7));
  inv1  gate625(.a(G28), .O(gate22inter8));
  nand2 gate626(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate627(.a(s_11), .b(gate22inter3), .O(gate22inter10));
  nor2  gate628(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate629(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate630(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate729(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate730(.a(gate23inter0), .b(s_26), .O(gate23inter1));
  and2  gate731(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate732(.a(s_26), .O(gate23inter3));
  inv1  gate733(.a(s_27), .O(gate23inter4));
  nand2 gate734(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate735(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate736(.a(G29), .O(gate23inter7));
  inv1  gate737(.a(G30), .O(gate23inter8));
  nand2 gate738(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate739(.a(s_27), .b(gate23inter3), .O(gate23inter10));
  nor2  gate740(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate741(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate742(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate575(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate576(.a(gate26inter0), .b(s_4), .O(gate26inter1));
  and2  gate577(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate578(.a(s_4), .O(gate26inter3));
  inv1  gate579(.a(s_5), .O(gate26inter4));
  nand2 gate580(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate581(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate582(.a(G9), .O(gate26inter7));
  inv1  gate583(.a(G13), .O(gate26inter8));
  nand2 gate584(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate585(.a(s_5), .b(gate26inter3), .O(gate26inter10));
  nor2  gate586(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate587(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate588(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate2213(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2214(.a(gate27inter0), .b(s_238), .O(gate27inter1));
  and2  gate2215(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2216(.a(s_238), .O(gate27inter3));
  inv1  gate2217(.a(s_239), .O(gate27inter4));
  nand2 gate2218(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2219(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2220(.a(G2), .O(gate27inter7));
  inv1  gate2221(.a(G6), .O(gate27inter8));
  nand2 gate2222(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2223(.a(s_239), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2224(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2225(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2226(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2577(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2578(.a(gate29inter0), .b(s_290), .O(gate29inter1));
  and2  gate2579(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2580(.a(s_290), .O(gate29inter3));
  inv1  gate2581(.a(s_291), .O(gate29inter4));
  nand2 gate2582(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2583(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2584(.a(G3), .O(gate29inter7));
  inv1  gate2585(.a(G7), .O(gate29inter8));
  nand2 gate2586(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2587(.a(s_291), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2588(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2589(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2590(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate547(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate548(.a(gate31inter0), .b(s_0), .O(gate31inter1));
  and2  gate549(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate550(.a(s_0), .O(gate31inter3));
  inv1  gate551(.a(s_1), .O(gate31inter4));
  nand2 gate552(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate553(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate554(.a(G4), .O(gate31inter7));
  inv1  gate555(.a(G8), .O(gate31inter8));
  nand2 gate556(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate557(.a(s_1), .b(gate31inter3), .O(gate31inter10));
  nor2  gate558(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate559(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate560(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate841(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate842(.a(gate36inter0), .b(s_42), .O(gate36inter1));
  and2  gate843(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate844(.a(s_42), .O(gate36inter3));
  inv1  gate845(.a(s_43), .O(gate36inter4));
  nand2 gate846(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate847(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate848(.a(G26), .O(gate36inter7));
  inv1  gate849(.a(G30), .O(gate36inter8));
  nand2 gate850(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate851(.a(s_43), .b(gate36inter3), .O(gate36inter10));
  nor2  gate852(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate853(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate854(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate995(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate996(.a(gate43inter0), .b(s_64), .O(gate43inter1));
  and2  gate997(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate998(.a(s_64), .O(gate43inter3));
  inv1  gate999(.a(s_65), .O(gate43inter4));
  nand2 gate1000(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1001(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1002(.a(G3), .O(gate43inter7));
  inv1  gate1003(.a(G269), .O(gate43inter8));
  nand2 gate1004(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1005(.a(s_65), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1006(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1007(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1008(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1149(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1150(.a(gate44inter0), .b(s_86), .O(gate44inter1));
  and2  gate1151(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1152(.a(s_86), .O(gate44inter3));
  inv1  gate1153(.a(s_87), .O(gate44inter4));
  nand2 gate1154(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1155(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1156(.a(G4), .O(gate44inter7));
  inv1  gate1157(.a(G269), .O(gate44inter8));
  nand2 gate1158(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1159(.a(s_87), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1160(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1161(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1162(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1611(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1612(.a(gate46inter0), .b(s_152), .O(gate46inter1));
  and2  gate1613(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1614(.a(s_152), .O(gate46inter3));
  inv1  gate1615(.a(s_153), .O(gate46inter4));
  nand2 gate1616(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1617(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1618(.a(G6), .O(gate46inter7));
  inv1  gate1619(.a(G272), .O(gate46inter8));
  nand2 gate1620(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1621(.a(s_153), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1622(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1623(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1624(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1387(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1388(.a(gate47inter0), .b(s_120), .O(gate47inter1));
  and2  gate1389(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1390(.a(s_120), .O(gate47inter3));
  inv1  gate1391(.a(s_121), .O(gate47inter4));
  nand2 gate1392(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1393(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1394(.a(G7), .O(gate47inter7));
  inv1  gate1395(.a(G275), .O(gate47inter8));
  nand2 gate1396(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1397(.a(s_121), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1398(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1399(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1400(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1107(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1108(.a(gate48inter0), .b(s_80), .O(gate48inter1));
  and2  gate1109(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1110(.a(s_80), .O(gate48inter3));
  inv1  gate1111(.a(s_81), .O(gate48inter4));
  nand2 gate1112(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1113(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1114(.a(G8), .O(gate48inter7));
  inv1  gate1115(.a(G275), .O(gate48inter8));
  nand2 gate1116(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1117(.a(s_81), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1118(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1119(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1120(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate3081(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate3082(.a(gate52inter0), .b(s_362), .O(gate52inter1));
  and2  gate3083(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate3084(.a(s_362), .O(gate52inter3));
  inv1  gate3085(.a(s_363), .O(gate52inter4));
  nand2 gate3086(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate3087(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate3088(.a(G12), .O(gate52inter7));
  inv1  gate3089(.a(G281), .O(gate52inter8));
  nand2 gate3090(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate3091(.a(s_363), .b(gate52inter3), .O(gate52inter10));
  nor2  gate3092(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate3093(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate3094(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1779(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1780(.a(gate53inter0), .b(s_176), .O(gate53inter1));
  and2  gate1781(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1782(.a(s_176), .O(gate53inter3));
  inv1  gate1783(.a(s_177), .O(gate53inter4));
  nand2 gate1784(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1785(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1786(.a(G13), .O(gate53inter7));
  inv1  gate1787(.a(G284), .O(gate53inter8));
  nand2 gate1788(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1789(.a(s_177), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1790(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1791(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1792(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1989(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1990(.a(gate55inter0), .b(s_206), .O(gate55inter1));
  and2  gate1991(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1992(.a(s_206), .O(gate55inter3));
  inv1  gate1993(.a(s_207), .O(gate55inter4));
  nand2 gate1994(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1995(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1996(.a(G15), .O(gate55inter7));
  inv1  gate1997(.a(G287), .O(gate55inter8));
  nand2 gate1998(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1999(.a(s_207), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2000(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2001(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2002(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate2913(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2914(.a(gate57inter0), .b(s_338), .O(gate57inter1));
  and2  gate2915(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2916(.a(s_338), .O(gate57inter3));
  inv1  gate2917(.a(s_339), .O(gate57inter4));
  nand2 gate2918(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2919(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2920(.a(G17), .O(gate57inter7));
  inv1  gate2921(.a(G290), .O(gate57inter8));
  nand2 gate2922(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2923(.a(s_339), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2924(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2925(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2926(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1457(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1458(.a(gate59inter0), .b(s_130), .O(gate59inter1));
  and2  gate1459(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1460(.a(s_130), .O(gate59inter3));
  inv1  gate1461(.a(s_131), .O(gate59inter4));
  nand2 gate1462(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1463(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1464(.a(G19), .O(gate59inter7));
  inv1  gate1465(.a(G293), .O(gate59inter8));
  nand2 gate1466(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1467(.a(s_131), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1468(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1469(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1470(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2885(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2886(.a(gate62inter0), .b(s_334), .O(gate62inter1));
  and2  gate2887(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2888(.a(s_334), .O(gate62inter3));
  inv1  gate2889(.a(s_335), .O(gate62inter4));
  nand2 gate2890(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2891(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2892(.a(G22), .O(gate62inter7));
  inv1  gate2893(.a(G296), .O(gate62inter8));
  nand2 gate2894(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2895(.a(s_335), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2896(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2897(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2898(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1051(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1052(.a(gate64inter0), .b(s_72), .O(gate64inter1));
  and2  gate1053(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1054(.a(s_72), .O(gate64inter3));
  inv1  gate1055(.a(s_73), .O(gate64inter4));
  nand2 gate1056(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1057(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1058(.a(G24), .O(gate64inter7));
  inv1  gate1059(.a(G299), .O(gate64inter8));
  nand2 gate1060(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1061(.a(s_73), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1062(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1063(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1064(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1065(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1066(.a(gate75inter0), .b(s_74), .O(gate75inter1));
  and2  gate1067(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1068(.a(s_74), .O(gate75inter3));
  inv1  gate1069(.a(s_75), .O(gate75inter4));
  nand2 gate1070(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1071(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1072(.a(G9), .O(gate75inter7));
  inv1  gate1073(.a(G317), .O(gate75inter8));
  nand2 gate1074(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1075(.a(s_75), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1076(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1077(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1078(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate813(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate814(.a(gate76inter0), .b(s_38), .O(gate76inter1));
  and2  gate815(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate816(.a(s_38), .O(gate76inter3));
  inv1  gate817(.a(s_39), .O(gate76inter4));
  nand2 gate818(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate819(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate820(.a(G13), .O(gate76inter7));
  inv1  gate821(.a(G317), .O(gate76inter8));
  nand2 gate822(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate823(.a(s_39), .b(gate76inter3), .O(gate76inter10));
  nor2  gate824(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate825(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate826(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2269(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2270(.a(gate84inter0), .b(s_246), .O(gate84inter1));
  and2  gate2271(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2272(.a(s_246), .O(gate84inter3));
  inv1  gate2273(.a(s_247), .O(gate84inter4));
  nand2 gate2274(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2275(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2276(.a(G15), .O(gate84inter7));
  inv1  gate2277(.a(G329), .O(gate84inter8));
  nand2 gate2278(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2279(.a(s_247), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2280(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2281(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2282(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2563(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2564(.a(gate87inter0), .b(s_288), .O(gate87inter1));
  and2  gate2565(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2566(.a(s_288), .O(gate87inter3));
  inv1  gate2567(.a(s_289), .O(gate87inter4));
  nand2 gate2568(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2569(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2570(.a(G12), .O(gate87inter7));
  inv1  gate2571(.a(G335), .O(gate87inter8));
  nand2 gate2572(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2573(.a(s_289), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2574(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2575(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2576(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1751(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1752(.a(gate88inter0), .b(s_172), .O(gate88inter1));
  and2  gate1753(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1754(.a(s_172), .O(gate88inter3));
  inv1  gate1755(.a(s_173), .O(gate88inter4));
  nand2 gate1756(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1757(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1758(.a(G16), .O(gate88inter7));
  inv1  gate1759(.a(G335), .O(gate88inter8));
  nand2 gate1760(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1761(.a(s_173), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1762(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1763(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1764(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1723(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1724(.a(gate89inter0), .b(s_168), .O(gate89inter1));
  and2  gate1725(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1726(.a(s_168), .O(gate89inter3));
  inv1  gate1727(.a(s_169), .O(gate89inter4));
  nand2 gate1728(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1729(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1730(.a(G17), .O(gate89inter7));
  inv1  gate1731(.a(G338), .O(gate89inter8));
  nand2 gate1732(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1733(.a(s_169), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1734(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1735(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1736(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2507(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2508(.a(gate91inter0), .b(s_280), .O(gate91inter1));
  and2  gate2509(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2510(.a(s_280), .O(gate91inter3));
  inv1  gate2511(.a(s_281), .O(gate91inter4));
  nand2 gate2512(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2513(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2514(.a(G25), .O(gate91inter7));
  inv1  gate2515(.a(G341), .O(gate91inter8));
  nand2 gate2516(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2517(.a(s_281), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2518(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2519(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2520(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate3207(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate3208(.a(gate95inter0), .b(s_380), .O(gate95inter1));
  and2  gate3209(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate3210(.a(s_380), .O(gate95inter3));
  inv1  gate3211(.a(s_381), .O(gate95inter4));
  nand2 gate3212(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate3213(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate3214(.a(G26), .O(gate95inter7));
  inv1  gate3215(.a(G347), .O(gate95inter8));
  nand2 gate3216(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate3217(.a(s_381), .b(gate95inter3), .O(gate95inter10));
  nor2  gate3218(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate3219(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate3220(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate561(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate562(.a(gate96inter0), .b(s_2), .O(gate96inter1));
  and2  gate563(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate564(.a(s_2), .O(gate96inter3));
  inv1  gate565(.a(s_3), .O(gate96inter4));
  nand2 gate566(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate567(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate568(.a(G30), .O(gate96inter7));
  inv1  gate569(.a(G347), .O(gate96inter8));
  nand2 gate570(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate571(.a(s_3), .b(gate96inter3), .O(gate96inter10));
  nor2  gate572(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate573(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate574(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1849(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1850(.a(gate98inter0), .b(s_186), .O(gate98inter1));
  and2  gate1851(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1852(.a(s_186), .O(gate98inter3));
  inv1  gate1853(.a(s_187), .O(gate98inter4));
  nand2 gate1854(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1855(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1856(.a(G23), .O(gate98inter7));
  inv1  gate1857(.a(G350), .O(gate98inter8));
  nand2 gate1858(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1859(.a(s_187), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1860(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1861(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1862(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate3137(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate3138(.a(gate100inter0), .b(s_370), .O(gate100inter1));
  and2  gate3139(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate3140(.a(s_370), .O(gate100inter3));
  inv1  gate3141(.a(s_371), .O(gate100inter4));
  nand2 gate3142(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate3143(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate3144(.a(G31), .O(gate100inter7));
  inv1  gate3145(.a(G353), .O(gate100inter8));
  nand2 gate3146(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate3147(.a(s_371), .b(gate100inter3), .O(gate100inter10));
  nor2  gate3148(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate3149(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate3150(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1079(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1080(.a(gate104inter0), .b(s_76), .O(gate104inter1));
  and2  gate1081(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1082(.a(s_76), .O(gate104inter3));
  inv1  gate1083(.a(s_77), .O(gate104inter4));
  nand2 gate1084(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1085(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1086(.a(G32), .O(gate104inter7));
  inv1  gate1087(.a(G359), .O(gate104inter8));
  nand2 gate1088(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1089(.a(s_77), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1090(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1091(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1092(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2773(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2774(.a(gate106inter0), .b(s_318), .O(gate106inter1));
  and2  gate2775(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2776(.a(s_318), .O(gate106inter3));
  inv1  gate2777(.a(s_319), .O(gate106inter4));
  nand2 gate2778(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2779(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2780(.a(G364), .O(gate106inter7));
  inv1  gate2781(.a(G365), .O(gate106inter8));
  nand2 gate2782(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2783(.a(s_319), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2784(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2785(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2786(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2199(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2200(.a(gate107inter0), .b(s_236), .O(gate107inter1));
  and2  gate2201(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2202(.a(s_236), .O(gate107inter3));
  inv1  gate2203(.a(s_237), .O(gate107inter4));
  nand2 gate2204(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2205(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2206(.a(G366), .O(gate107inter7));
  inv1  gate2207(.a(G367), .O(gate107inter8));
  nand2 gate2208(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2209(.a(s_237), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2210(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2211(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2212(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate925(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate926(.a(gate109inter0), .b(s_54), .O(gate109inter1));
  and2  gate927(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate928(.a(s_54), .O(gate109inter3));
  inv1  gate929(.a(s_55), .O(gate109inter4));
  nand2 gate930(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate931(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate932(.a(G370), .O(gate109inter7));
  inv1  gate933(.a(G371), .O(gate109inter8));
  nand2 gate934(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate935(.a(s_55), .b(gate109inter3), .O(gate109inter10));
  nor2  gate936(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate937(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate938(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1219(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1220(.a(gate112inter0), .b(s_96), .O(gate112inter1));
  and2  gate1221(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1222(.a(s_96), .O(gate112inter3));
  inv1  gate1223(.a(s_97), .O(gate112inter4));
  nand2 gate1224(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1225(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1226(.a(G376), .O(gate112inter7));
  inv1  gate1227(.a(G377), .O(gate112inter8));
  nand2 gate1228(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1229(.a(s_97), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1230(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1231(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1232(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate2101(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2102(.a(gate113inter0), .b(s_222), .O(gate113inter1));
  and2  gate2103(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2104(.a(s_222), .O(gate113inter3));
  inv1  gate2105(.a(s_223), .O(gate113inter4));
  nand2 gate2106(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2107(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2108(.a(G378), .O(gate113inter7));
  inv1  gate2109(.a(G379), .O(gate113inter8));
  nand2 gate2110(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2111(.a(s_223), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2112(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2113(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2114(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1919(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1920(.a(gate116inter0), .b(s_196), .O(gate116inter1));
  and2  gate1921(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1922(.a(s_196), .O(gate116inter3));
  inv1  gate1923(.a(s_197), .O(gate116inter4));
  nand2 gate1924(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1925(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1926(.a(G384), .O(gate116inter7));
  inv1  gate1927(.a(G385), .O(gate116inter8));
  nand2 gate1928(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1929(.a(s_197), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1930(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1931(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1932(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1765(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1766(.a(gate118inter0), .b(s_174), .O(gate118inter1));
  and2  gate1767(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1768(.a(s_174), .O(gate118inter3));
  inv1  gate1769(.a(s_175), .O(gate118inter4));
  nand2 gate1770(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1771(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1772(.a(G388), .O(gate118inter7));
  inv1  gate1773(.a(G389), .O(gate118inter8));
  nand2 gate1774(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1775(.a(s_175), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1776(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1777(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1778(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate785(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate786(.a(gate120inter0), .b(s_34), .O(gate120inter1));
  and2  gate787(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate788(.a(s_34), .O(gate120inter3));
  inv1  gate789(.a(s_35), .O(gate120inter4));
  nand2 gate790(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate791(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate792(.a(G392), .O(gate120inter7));
  inv1  gate793(.a(G393), .O(gate120inter8));
  nand2 gate794(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate795(.a(s_35), .b(gate120inter3), .O(gate120inter10));
  nor2  gate796(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate797(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate798(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1807(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1808(.a(gate121inter0), .b(s_180), .O(gate121inter1));
  and2  gate1809(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1810(.a(s_180), .O(gate121inter3));
  inv1  gate1811(.a(s_181), .O(gate121inter4));
  nand2 gate1812(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1813(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1814(.a(G394), .O(gate121inter7));
  inv1  gate1815(.a(G395), .O(gate121inter8));
  nand2 gate1816(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1817(.a(s_181), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1818(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1819(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1820(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2675(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2676(.a(gate122inter0), .b(s_304), .O(gate122inter1));
  and2  gate2677(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2678(.a(s_304), .O(gate122inter3));
  inv1  gate2679(.a(s_305), .O(gate122inter4));
  nand2 gate2680(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2681(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2682(.a(G396), .O(gate122inter7));
  inv1  gate2683(.a(G397), .O(gate122inter8));
  nand2 gate2684(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2685(.a(s_305), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2686(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2687(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2688(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2801(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2802(.a(gate125inter0), .b(s_322), .O(gate125inter1));
  and2  gate2803(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2804(.a(s_322), .O(gate125inter3));
  inv1  gate2805(.a(s_323), .O(gate125inter4));
  nand2 gate2806(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2807(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2808(.a(G402), .O(gate125inter7));
  inv1  gate2809(.a(G403), .O(gate125inter8));
  nand2 gate2810(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2811(.a(s_323), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2812(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2813(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2814(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1471(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1472(.a(gate126inter0), .b(s_132), .O(gate126inter1));
  and2  gate1473(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1474(.a(s_132), .O(gate126inter3));
  inv1  gate1475(.a(s_133), .O(gate126inter4));
  nand2 gate1476(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1477(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1478(.a(G404), .O(gate126inter7));
  inv1  gate1479(.a(G405), .O(gate126inter8));
  nand2 gate1480(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1481(.a(s_133), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1482(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1483(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1484(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2381(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2382(.a(gate129inter0), .b(s_262), .O(gate129inter1));
  and2  gate2383(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2384(.a(s_262), .O(gate129inter3));
  inv1  gate2385(.a(s_263), .O(gate129inter4));
  nand2 gate2386(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2387(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2388(.a(G410), .O(gate129inter7));
  inv1  gate2389(.a(G411), .O(gate129inter8));
  nand2 gate2390(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2391(.a(s_263), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2392(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2393(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2394(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2003(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2004(.a(gate130inter0), .b(s_208), .O(gate130inter1));
  and2  gate2005(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2006(.a(s_208), .O(gate130inter3));
  inv1  gate2007(.a(s_209), .O(gate130inter4));
  nand2 gate2008(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2009(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2010(.a(G412), .O(gate130inter7));
  inv1  gate2011(.a(G413), .O(gate130inter8));
  nand2 gate2012(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2013(.a(s_209), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2014(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2015(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2016(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1709(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1710(.a(gate131inter0), .b(s_166), .O(gate131inter1));
  and2  gate1711(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1712(.a(s_166), .O(gate131inter3));
  inv1  gate1713(.a(s_167), .O(gate131inter4));
  nand2 gate1714(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1715(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1716(.a(G414), .O(gate131inter7));
  inv1  gate1717(.a(G415), .O(gate131inter8));
  nand2 gate1718(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1719(.a(s_167), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1720(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1721(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1722(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate911(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate912(.a(gate133inter0), .b(s_52), .O(gate133inter1));
  and2  gate913(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate914(.a(s_52), .O(gate133inter3));
  inv1  gate915(.a(s_53), .O(gate133inter4));
  nand2 gate916(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate917(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate918(.a(G418), .O(gate133inter7));
  inv1  gate919(.a(G419), .O(gate133inter8));
  nand2 gate920(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate921(.a(s_53), .b(gate133inter3), .O(gate133inter10));
  nor2  gate922(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate923(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate924(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate2997(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2998(.a(gate134inter0), .b(s_350), .O(gate134inter1));
  and2  gate2999(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate3000(.a(s_350), .O(gate134inter3));
  inv1  gate3001(.a(s_351), .O(gate134inter4));
  nand2 gate3002(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate3003(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate3004(.a(G420), .O(gate134inter7));
  inv1  gate3005(.a(G421), .O(gate134inter8));
  nand2 gate3006(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate3007(.a(s_351), .b(gate134inter3), .O(gate134inter10));
  nor2  gate3008(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate3009(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate3010(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1261(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1262(.a(gate137inter0), .b(s_102), .O(gate137inter1));
  and2  gate1263(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1264(.a(s_102), .O(gate137inter3));
  inv1  gate1265(.a(s_103), .O(gate137inter4));
  nand2 gate1266(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1267(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1268(.a(G426), .O(gate137inter7));
  inv1  gate1269(.a(G429), .O(gate137inter8));
  nand2 gate1270(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1271(.a(s_103), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1272(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1273(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1274(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate3151(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate3152(.a(gate141inter0), .b(s_372), .O(gate141inter1));
  and2  gate3153(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate3154(.a(s_372), .O(gate141inter3));
  inv1  gate3155(.a(s_373), .O(gate141inter4));
  nand2 gate3156(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate3157(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate3158(.a(G450), .O(gate141inter7));
  inv1  gate3159(.a(G453), .O(gate141inter8));
  nand2 gate3160(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate3161(.a(s_373), .b(gate141inter3), .O(gate141inter10));
  nor2  gate3162(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate3163(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate3164(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate3053(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate3054(.a(gate143inter0), .b(s_358), .O(gate143inter1));
  and2  gate3055(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate3056(.a(s_358), .O(gate143inter3));
  inv1  gate3057(.a(s_359), .O(gate143inter4));
  nand2 gate3058(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate3059(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate3060(.a(G462), .O(gate143inter7));
  inv1  gate3061(.a(G465), .O(gate143inter8));
  nand2 gate3062(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate3063(.a(s_359), .b(gate143inter3), .O(gate143inter10));
  nor2  gate3064(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate3065(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate3066(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate3109(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate3110(.a(gate144inter0), .b(s_366), .O(gate144inter1));
  and2  gate3111(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate3112(.a(s_366), .O(gate144inter3));
  inv1  gate3113(.a(s_367), .O(gate144inter4));
  nand2 gate3114(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate3115(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate3116(.a(G468), .O(gate144inter7));
  inv1  gate3117(.a(G471), .O(gate144inter8));
  nand2 gate3118(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate3119(.a(s_367), .b(gate144inter3), .O(gate144inter10));
  nor2  gate3120(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate3121(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate3122(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2647(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2648(.a(gate147inter0), .b(s_300), .O(gate147inter1));
  and2  gate2649(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2650(.a(s_300), .O(gate147inter3));
  inv1  gate2651(.a(s_301), .O(gate147inter4));
  nand2 gate2652(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2653(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2654(.a(G486), .O(gate147inter7));
  inv1  gate2655(.a(G489), .O(gate147inter8));
  nand2 gate2656(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2657(.a(s_301), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2658(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2659(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2660(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate981(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate982(.a(gate150inter0), .b(s_62), .O(gate150inter1));
  and2  gate983(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate984(.a(s_62), .O(gate150inter3));
  inv1  gate985(.a(s_63), .O(gate150inter4));
  nand2 gate986(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate987(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate988(.a(G504), .O(gate150inter7));
  inv1  gate989(.a(G507), .O(gate150inter8));
  nand2 gate990(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate991(.a(s_63), .b(gate150inter3), .O(gate150inter10));
  nor2  gate992(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate993(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate994(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1233(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1234(.a(gate151inter0), .b(s_98), .O(gate151inter1));
  and2  gate1235(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1236(.a(s_98), .O(gate151inter3));
  inv1  gate1237(.a(s_99), .O(gate151inter4));
  nand2 gate1238(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1239(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1240(.a(G510), .O(gate151inter7));
  inv1  gate1241(.a(G513), .O(gate151inter8));
  nand2 gate1242(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1243(.a(s_99), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1244(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1245(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1246(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1093(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1094(.a(gate156inter0), .b(s_78), .O(gate156inter1));
  and2  gate1095(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1096(.a(s_78), .O(gate156inter3));
  inv1  gate1097(.a(s_79), .O(gate156inter4));
  nand2 gate1098(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1099(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1100(.a(G435), .O(gate156inter7));
  inv1  gate1101(.a(G525), .O(gate156inter8));
  nand2 gate1102(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1103(.a(s_79), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1104(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1105(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1106(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1639(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1640(.a(gate157inter0), .b(s_156), .O(gate157inter1));
  and2  gate1641(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1642(.a(s_156), .O(gate157inter3));
  inv1  gate1643(.a(s_157), .O(gate157inter4));
  nand2 gate1644(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1645(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1646(.a(G438), .O(gate157inter7));
  inv1  gate1647(.a(G528), .O(gate157inter8));
  nand2 gate1648(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1649(.a(s_157), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1650(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1651(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1652(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2493(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2494(.a(gate158inter0), .b(s_278), .O(gate158inter1));
  and2  gate2495(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2496(.a(s_278), .O(gate158inter3));
  inv1  gate2497(.a(s_279), .O(gate158inter4));
  nand2 gate2498(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2499(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2500(.a(G441), .O(gate158inter7));
  inv1  gate2501(.a(G528), .O(gate158inter8));
  nand2 gate2502(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2503(.a(s_279), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2504(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2505(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2506(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1737(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1738(.a(gate159inter0), .b(s_170), .O(gate159inter1));
  and2  gate1739(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1740(.a(s_170), .O(gate159inter3));
  inv1  gate1741(.a(s_171), .O(gate159inter4));
  nand2 gate1742(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1743(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1744(.a(G444), .O(gate159inter7));
  inv1  gate1745(.a(G531), .O(gate159inter8));
  nand2 gate1746(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1747(.a(s_171), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1748(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1749(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1750(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate701(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate702(.a(gate164inter0), .b(s_22), .O(gate164inter1));
  and2  gate703(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate704(.a(s_22), .O(gate164inter3));
  inv1  gate705(.a(s_23), .O(gate164inter4));
  nand2 gate706(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate707(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate708(.a(G459), .O(gate164inter7));
  inv1  gate709(.a(G537), .O(gate164inter8));
  nand2 gate710(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate711(.a(s_23), .b(gate164inter3), .O(gate164inter10));
  nor2  gate712(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate713(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate714(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate1009(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1010(.a(gate165inter0), .b(s_66), .O(gate165inter1));
  and2  gate1011(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1012(.a(s_66), .O(gate165inter3));
  inv1  gate1013(.a(s_67), .O(gate165inter4));
  nand2 gate1014(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1015(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1016(.a(G462), .O(gate165inter7));
  inv1  gate1017(.a(G540), .O(gate165inter8));
  nand2 gate1018(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1019(.a(s_67), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1020(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1021(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1022(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate771(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate772(.a(gate166inter0), .b(s_32), .O(gate166inter1));
  and2  gate773(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate774(.a(s_32), .O(gate166inter3));
  inv1  gate775(.a(s_33), .O(gate166inter4));
  nand2 gate776(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate777(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate778(.a(G465), .O(gate166inter7));
  inv1  gate779(.a(G540), .O(gate166inter8));
  nand2 gate780(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate781(.a(s_33), .b(gate166inter3), .O(gate166inter10));
  nor2  gate782(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate783(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate784(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate3123(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate3124(.a(gate167inter0), .b(s_368), .O(gate167inter1));
  and2  gate3125(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate3126(.a(s_368), .O(gate167inter3));
  inv1  gate3127(.a(s_369), .O(gate167inter4));
  nand2 gate3128(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate3129(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate3130(.a(G468), .O(gate167inter7));
  inv1  gate3131(.a(G543), .O(gate167inter8));
  nand2 gate3132(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate3133(.a(s_369), .b(gate167inter3), .O(gate167inter10));
  nor2  gate3134(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate3135(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate3136(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1793(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1794(.a(gate170inter0), .b(s_178), .O(gate170inter1));
  and2  gate1795(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1796(.a(s_178), .O(gate170inter3));
  inv1  gate1797(.a(s_179), .O(gate170inter4));
  nand2 gate1798(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1799(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1800(.a(G477), .O(gate170inter7));
  inv1  gate1801(.a(G546), .O(gate170inter8));
  nand2 gate1802(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1803(.a(s_179), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1804(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1805(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1806(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1863(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1864(.a(gate171inter0), .b(s_188), .O(gate171inter1));
  and2  gate1865(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1866(.a(s_188), .O(gate171inter3));
  inv1  gate1867(.a(s_189), .O(gate171inter4));
  nand2 gate1868(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1869(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1870(.a(G480), .O(gate171inter7));
  inv1  gate1871(.a(G549), .O(gate171inter8));
  nand2 gate1872(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1873(.a(s_189), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1874(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1875(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1876(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2115(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2116(.a(gate172inter0), .b(s_224), .O(gate172inter1));
  and2  gate2117(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2118(.a(s_224), .O(gate172inter3));
  inv1  gate2119(.a(s_225), .O(gate172inter4));
  nand2 gate2120(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2121(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2122(.a(G483), .O(gate172inter7));
  inv1  gate2123(.a(G549), .O(gate172inter8));
  nand2 gate2124(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2125(.a(s_225), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2126(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2127(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2128(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate953(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate954(.a(gate173inter0), .b(s_58), .O(gate173inter1));
  and2  gate955(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate956(.a(s_58), .O(gate173inter3));
  inv1  gate957(.a(s_59), .O(gate173inter4));
  nand2 gate958(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate959(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate960(.a(G486), .O(gate173inter7));
  inv1  gate961(.a(G552), .O(gate173inter8));
  nand2 gate962(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate963(.a(s_59), .b(gate173inter3), .O(gate173inter10));
  nor2  gate964(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate965(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate966(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2087(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2088(.a(gate176inter0), .b(s_220), .O(gate176inter1));
  and2  gate2089(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2090(.a(s_220), .O(gate176inter3));
  inv1  gate2091(.a(s_221), .O(gate176inter4));
  nand2 gate2092(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2093(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2094(.a(G495), .O(gate176inter7));
  inv1  gate2095(.a(G555), .O(gate176inter8));
  nand2 gate2096(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2097(.a(s_221), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2098(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2099(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2100(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2927(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2928(.a(gate179inter0), .b(s_340), .O(gate179inter1));
  and2  gate2929(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2930(.a(s_340), .O(gate179inter3));
  inv1  gate2931(.a(s_341), .O(gate179inter4));
  nand2 gate2932(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2933(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2934(.a(G504), .O(gate179inter7));
  inv1  gate2935(.a(G561), .O(gate179inter8));
  nand2 gate2936(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2937(.a(s_341), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2938(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2939(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2940(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate2745(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2746(.a(gate180inter0), .b(s_314), .O(gate180inter1));
  and2  gate2747(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2748(.a(s_314), .O(gate180inter3));
  inv1  gate2749(.a(s_315), .O(gate180inter4));
  nand2 gate2750(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2751(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2752(.a(G507), .O(gate180inter7));
  inv1  gate2753(.a(G561), .O(gate180inter8));
  nand2 gate2754(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2755(.a(s_315), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2756(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2757(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2758(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1177(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1178(.a(gate181inter0), .b(s_90), .O(gate181inter1));
  and2  gate1179(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1180(.a(s_90), .O(gate181inter3));
  inv1  gate1181(.a(s_91), .O(gate181inter4));
  nand2 gate1182(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1183(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1184(.a(G510), .O(gate181inter7));
  inv1  gate1185(.a(G564), .O(gate181inter8));
  nand2 gate1186(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1187(.a(s_91), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1188(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1189(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1190(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2395(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2396(.a(gate182inter0), .b(s_264), .O(gate182inter1));
  and2  gate2397(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2398(.a(s_264), .O(gate182inter3));
  inv1  gate2399(.a(s_265), .O(gate182inter4));
  nand2 gate2400(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2401(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2402(.a(G513), .O(gate182inter7));
  inv1  gate2403(.a(G564), .O(gate182inter8));
  nand2 gate2404(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2405(.a(s_265), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2406(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2407(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2408(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate715(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate716(.a(gate183inter0), .b(s_24), .O(gate183inter1));
  and2  gate717(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate718(.a(s_24), .O(gate183inter3));
  inv1  gate719(.a(s_25), .O(gate183inter4));
  nand2 gate720(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate721(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate722(.a(G516), .O(gate183inter7));
  inv1  gate723(.a(G567), .O(gate183inter8));
  nand2 gate724(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate725(.a(s_25), .b(gate183inter3), .O(gate183inter10));
  nor2  gate726(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate727(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate728(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1835(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1836(.a(gate185inter0), .b(s_184), .O(gate185inter1));
  and2  gate1837(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1838(.a(s_184), .O(gate185inter3));
  inv1  gate1839(.a(s_185), .O(gate185inter4));
  nand2 gate1840(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1841(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1842(.a(G570), .O(gate185inter7));
  inv1  gate1843(.a(G571), .O(gate185inter8));
  nand2 gate1844(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1845(.a(s_185), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1846(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1847(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1848(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1121(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1122(.a(gate186inter0), .b(s_82), .O(gate186inter1));
  and2  gate1123(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1124(.a(s_82), .O(gate186inter3));
  inv1  gate1125(.a(s_83), .O(gate186inter4));
  nand2 gate1126(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1127(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1128(.a(G572), .O(gate186inter7));
  inv1  gate1129(.a(G573), .O(gate186inter8));
  nand2 gate1130(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1131(.a(s_83), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1132(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1133(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1134(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1247(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1248(.a(gate187inter0), .b(s_100), .O(gate187inter1));
  and2  gate1249(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1250(.a(s_100), .O(gate187inter3));
  inv1  gate1251(.a(s_101), .O(gate187inter4));
  nand2 gate1252(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1253(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1254(.a(G574), .O(gate187inter7));
  inv1  gate1255(.a(G575), .O(gate187inter8));
  nand2 gate1256(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1257(.a(s_101), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1258(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1259(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1260(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2255(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2256(.a(gate188inter0), .b(s_244), .O(gate188inter1));
  and2  gate2257(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2258(.a(s_244), .O(gate188inter3));
  inv1  gate2259(.a(s_245), .O(gate188inter4));
  nand2 gate2260(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2261(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2262(.a(G576), .O(gate188inter7));
  inv1  gate2263(.a(G577), .O(gate188inter8));
  nand2 gate2264(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2265(.a(s_245), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2266(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2267(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2268(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate3165(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate3166(.a(gate189inter0), .b(s_374), .O(gate189inter1));
  and2  gate3167(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate3168(.a(s_374), .O(gate189inter3));
  inv1  gate3169(.a(s_375), .O(gate189inter4));
  nand2 gate3170(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate3171(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate3172(.a(G578), .O(gate189inter7));
  inv1  gate3173(.a(G579), .O(gate189inter8));
  nand2 gate3174(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate3175(.a(s_375), .b(gate189inter3), .O(gate189inter10));
  nor2  gate3176(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate3177(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate3178(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate967(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate968(.a(gate192inter0), .b(s_60), .O(gate192inter1));
  and2  gate969(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate970(.a(s_60), .O(gate192inter3));
  inv1  gate971(.a(s_61), .O(gate192inter4));
  nand2 gate972(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate973(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate974(.a(G584), .O(gate192inter7));
  inv1  gate975(.a(G585), .O(gate192inter8));
  nand2 gate976(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate977(.a(s_61), .b(gate192inter3), .O(gate192inter10));
  nor2  gate978(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate979(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate980(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2073(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2074(.a(gate193inter0), .b(s_218), .O(gate193inter1));
  and2  gate2075(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2076(.a(s_218), .O(gate193inter3));
  inv1  gate2077(.a(s_219), .O(gate193inter4));
  nand2 gate2078(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2079(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2080(.a(G586), .O(gate193inter7));
  inv1  gate2081(.a(G587), .O(gate193inter8));
  nand2 gate2082(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2083(.a(s_219), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2084(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2085(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2086(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate2703(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2704(.a(gate196inter0), .b(s_308), .O(gate196inter1));
  and2  gate2705(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2706(.a(s_308), .O(gate196inter3));
  inv1  gate2707(.a(s_309), .O(gate196inter4));
  nand2 gate2708(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2709(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2710(.a(G592), .O(gate196inter7));
  inv1  gate2711(.a(G593), .O(gate196inter8));
  nand2 gate2712(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2713(.a(s_309), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2714(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2715(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2716(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1821(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1822(.a(gate197inter0), .b(s_182), .O(gate197inter1));
  and2  gate1823(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1824(.a(s_182), .O(gate197inter3));
  inv1  gate1825(.a(s_183), .O(gate197inter4));
  nand2 gate1826(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1827(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1828(.a(G594), .O(gate197inter7));
  inv1  gate1829(.a(G595), .O(gate197inter8));
  nand2 gate1830(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1831(.a(s_183), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1832(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1833(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1834(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate2045(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2046(.a(gate198inter0), .b(s_214), .O(gate198inter1));
  and2  gate2047(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2048(.a(s_214), .O(gate198inter3));
  inv1  gate2049(.a(s_215), .O(gate198inter4));
  nand2 gate2050(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2051(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2052(.a(G596), .O(gate198inter7));
  inv1  gate2053(.a(G597), .O(gate198inter8));
  nand2 gate2054(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2055(.a(s_215), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2056(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2057(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2058(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1317(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1318(.a(gate201inter0), .b(s_110), .O(gate201inter1));
  and2  gate1319(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1320(.a(s_110), .O(gate201inter3));
  inv1  gate1321(.a(s_111), .O(gate201inter4));
  nand2 gate1322(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1323(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1324(.a(G602), .O(gate201inter7));
  inv1  gate1325(.a(G607), .O(gate201inter8));
  nand2 gate1326(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1327(.a(s_111), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1328(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1329(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1330(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2857(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2858(.a(gate203inter0), .b(s_330), .O(gate203inter1));
  and2  gate2859(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2860(.a(s_330), .O(gate203inter3));
  inv1  gate2861(.a(s_331), .O(gate203inter4));
  nand2 gate2862(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2863(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2864(.a(G602), .O(gate203inter7));
  inv1  gate2865(.a(G612), .O(gate203inter8));
  nand2 gate2866(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2867(.a(s_331), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2868(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2869(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2870(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate2815(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2816(.a(gate204inter0), .b(s_324), .O(gate204inter1));
  and2  gate2817(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2818(.a(s_324), .O(gate204inter3));
  inv1  gate2819(.a(s_325), .O(gate204inter4));
  nand2 gate2820(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2821(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2822(.a(G607), .O(gate204inter7));
  inv1  gate2823(.a(G617), .O(gate204inter8));
  nand2 gate2824(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2825(.a(s_325), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2826(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2827(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2828(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2689(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2690(.a(gate206inter0), .b(s_306), .O(gate206inter1));
  and2  gate2691(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2692(.a(s_306), .O(gate206inter3));
  inv1  gate2693(.a(s_307), .O(gate206inter4));
  nand2 gate2694(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2695(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2696(.a(G632), .O(gate206inter7));
  inv1  gate2697(.a(G637), .O(gate206inter8));
  nand2 gate2698(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2699(.a(s_307), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2700(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2701(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2702(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2983(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2984(.a(gate207inter0), .b(s_348), .O(gate207inter1));
  and2  gate2985(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2986(.a(s_348), .O(gate207inter3));
  inv1  gate2987(.a(s_349), .O(gate207inter4));
  nand2 gate2988(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2989(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2990(.a(G622), .O(gate207inter7));
  inv1  gate2991(.a(G632), .O(gate207inter8));
  nand2 gate2992(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2993(.a(s_349), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2994(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2995(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2996(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate827(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate828(.a(gate208inter0), .b(s_40), .O(gate208inter1));
  and2  gate829(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate830(.a(s_40), .O(gate208inter3));
  inv1  gate831(.a(s_41), .O(gate208inter4));
  nand2 gate832(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate833(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate834(.a(G627), .O(gate208inter7));
  inv1  gate835(.a(G637), .O(gate208inter8));
  nand2 gate836(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate837(.a(s_41), .b(gate208inter3), .O(gate208inter10));
  nor2  gate838(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate839(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate840(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2479(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2480(.a(gate209inter0), .b(s_276), .O(gate209inter1));
  and2  gate2481(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2482(.a(s_276), .O(gate209inter3));
  inv1  gate2483(.a(s_277), .O(gate209inter4));
  nand2 gate2484(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2485(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2486(.a(G602), .O(gate209inter7));
  inv1  gate2487(.a(G666), .O(gate209inter8));
  nand2 gate2488(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2489(.a(s_277), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2490(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2491(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2492(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2409(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2410(.a(gate210inter0), .b(s_266), .O(gate210inter1));
  and2  gate2411(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2412(.a(s_266), .O(gate210inter3));
  inv1  gate2413(.a(s_267), .O(gate210inter4));
  nand2 gate2414(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2415(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2416(.a(G607), .O(gate210inter7));
  inv1  gate2417(.a(G666), .O(gate210inter8));
  nand2 gate2418(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2419(.a(s_267), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2420(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2421(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2422(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1933(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1934(.a(gate211inter0), .b(s_198), .O(gate211inter1));
  and2  gate1935(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1936(.a(s_198), .O(gate211inter3));
  inv1  gate1937(.a(s_199), .O(gate211inter4));
  nand2 gate1938(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1939(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1940(.a(G612), .O(gate211inter7));
  inv1  gate1941(.a(G669), .O(gate211inter8));
  nand2 gate1942(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1943(.a(s_199), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1944(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1945(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1946(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1163(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1164(.a(gate216inter0), .b(s_88), .O(gate216inter1));
  and2  gate1165(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1166(.a(s_88), .O(gate216inter3));
  inv1  gate1167(.a(s_89), .O(gate216inter4));
  nand2 gate1168(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1169(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1170(.a(G617), .O(gate216inter7));
  inv1  gate1171(.a(G675), .O(gate216inter8));
  nand2 gate1172(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1173(.a(s_89), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1174(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1175(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1176(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1891(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1892(.a(gate217inter0), .b(s_192), .O(gate217inter1));
  and2  gate1893(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1894(.a(s_192), .O(gate217inter3));
  inv1  gate1895(.a(s_193), .O(gate217inter4));
  nand2 gate1896(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1897(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1898(.a(G622), .O(gate217inter7));
  inv1  gate1899(.a(G678), .O(gate217inter8));
  nand2 gate1900(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1901(.a(s_193), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1902(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1903(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1904(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate645(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate646(.a(gate222inter0), .b(s_14), .O(gate222inter1));
  and2  gate647(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate648(.a(s_14), .O(gate222inter3));
  inv1  gate649(.a(s_15), .O(gate222inter4));
  nand2 gate650(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate651(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate652(.a(G632), .O(gate222inter7));
  inv1  gate653(.a(G684), .O(gate222inter8));
  nand2 gate654(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate655(.a(s_15), .b(gate222inter3), .O(gate222inter10));
  nor2  gate656(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate657(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate658(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1555(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1556(.a(gate224inter0), .b(s_144), .O(gate224inter1));
  and2  gate1557(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1558(.a(s_144), .O(gate224inter3));
  inv1  gate1559(.a(s_145), .O(gate224inter4));
  nand2 gate1560(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1561(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1562(.a(G637), .O(gate224inter7));
  inv1  gate1563(.a(G687), .O(gate224inter8));
  nand2 gate1564(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1565(.a(s_145), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1566(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1567(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1568(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate2367(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate2368(.a(gate226inter0), .b(s_260), .O(gate226inter1));
  and2  gate2369(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate2370(.a(s_260), .O(gate226inter3));
  inv1  gate2371(.a(s_261), .O(gate226inter4));
  nand2 gate2372(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate2373(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate2374(.a(G692), .O(gate226inter7));
  inv1  gate2375(.a(G693), .O(gate226inter8));
  nand2 gate2376(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate2377(.a(s_261), .b(gate226inter3), .O(gate226inter10));
  nor2  gate2378(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate2379(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate2380(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2717(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2718(.a(gate229inter0), .b(s_310), .O(gate229inter1));
  and2  gate2719(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2720(.a(s_310), .O(gate229inter3));
  inv1  gate2721(.a(s_311), .O(gate229inter4));
  nand2 gate2722(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2723(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2724(.a(G698), .O(gate229inter7));
  inv1  gate2725(.a(G699), .O(gate229inter8));
  nand2 gate2726(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2727(.a(s_311), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2728(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2729(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2730(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2661(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2662(.a(gate231inter0), .b(s_302), .O(gate231inter1));
  and2  gate2663(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2664(.a(s_302), .O(gate231inter3));
  inv1  gate2665(.a(s_303), .O(gate231inter4));
  nand2 gate2666(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2667(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2668(.a(G702), .O(gate231inter7));
  inv1  gate2669(.a(G703), .O(gate231inter8));
  nand2 gate2670(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2671(.a(s_303), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2672(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2673(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2674(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2787(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2788(.a(gate233inter0), .b(s_320), .O(gate233inter1));
  and2  gate2789(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2790(.a(s_320), .O(gate233inter3));
  inv1  gate2791(.a(s_321), .O(gate233inter4));
  nand2 gate2792(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2793(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2794(.a(G242), .O(gate233inter7));
  inv1  gate2795(.a(G718), .O(gate233inter8));
  nand2 gate2796(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2797(.a(s_321), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2798(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2799(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2800(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1541(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1542(.a(gate234inter0), .b(s_142), .O(gate234inter1));
  and2  gate1543(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1544(.a(s_142), .O(gate234inter3));
  inv1  gate1545(.a(s_143), .O(gate234inter4));
  nand2 gate1546(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1547(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1548(.a(G245), .O(gate234inter7));
  inv1  gate1549(.a(G721), .O(gate234inter8));
  nand2 gate1550(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1551(.a(s_143), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1552(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1553(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1554(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2311(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2312(.a(gate236inter0), .b(s_252), .O(gate236inter1));
  and2  gate2313(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2314(.a(s_252), .O(gate236inter3));
  inv1  gate2315(.a(s_253), .O(gate236inter4));
  nand2 gate2316(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2317(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2318(.a(G251), .O(gate236inter7));
  inv1  gate2319(.a(G727), .O(gate236inter8));
  nand2 gate2320(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2321(.a(s_253), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2322(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2323(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2324(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1513(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1514(.a(gate237inter0), .b(s_138), .O(gate237inter1));
  and2  gate1515(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1516(.a(s_138), .O(gate237inter3));
  inv1  gate1517(.a(s_139), .O(gate237inter4));
  nand2 gate1518(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1519(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1520(.a(G254), .O(gate237inter7));
  inv1  gate1521(.a(G706), .O(gate237inter8));
  nand2 gate1522(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1523(.a(s_139), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1524(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1525(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1526(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate2437(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2438(.a(gate238inter0), .b(s_270), .O(gate238inter1));
  and2  gate2439(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2440(.a(s_270), .O(gate238inter3));
  inv1  gate2441(.a(s_271), .O(gate238inter4));
  nand2 gate2442(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2443(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2444(.a(G257), .O(gate238inter7));
  inv1  gate2445(.a(G709), .O(gate238inter8));
  nand2 gate2446(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2447(.a(s_271), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2448(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2449(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2450(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate869(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate870(.a(gate241inter0), .b(s_46), .O(gate241inter1));
  and2  gate871(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate872(.a(s_46), .O(gate241inter3));
  inv1  gate873(.a(s_47), .O(gate241inter4));
  nand2 gate874(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate875(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate876(.a(G242), .O(gate241inter7));
  inv1  gate877(.a(G730), .O(gate241inter8));
  nand2 gate878(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate879(.a(s_47), .b(gate241inter3), .O(gate241inter10));
  nor2  gate880(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate881(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate882(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1415(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1416(.a(gate246inter0), .b(s_124), .O(gate246inter1));
  and2  gate1417(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1418(.a(s_124), .O(gate246inter3));
  inv1  gate1419(.a(s_125), .O(gate246inter4));
  nand2 gate1420(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1421(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1422(.a(G724), .O(gate246inter7));
  inv1  gate1423(.a(G736), .O(gate246inter8));
  nand2 gate1424(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1425(.a(s_125), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1426(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1427(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1428(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2227(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2228(.a(gate248inter0), .b(s_240), .O(gate248inter1));
  and2  gate2229(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2230(.a(s_240), .O(gate248inter3));
  inv1  gate2231(.a(s_241), .O(gate248inter4));
  nand2 gate2232(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2233(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2234(.a(G727), .O(gate248inter7));
  inv1  gate2235(.a(G739), .O(gate248inter8));
  nand2 gate2236(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2237(.a(s_241), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2238(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2239(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2240(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1681(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1682(.a(gate249inter0), .b(s_162), .O(gate249inter1));
  and2  gate1683(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1684(.a(s_162), .O(gate249inter3));
  inv1  gate1685(.a(s_163), .O(gate249inter4));
  nand2 gate1686(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1687(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1688(.a(G254), .O(gate249inter7));
  inv1  gate1689(.a(G742), .O(gate249inter8));
  nand2 gate1690(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1691(.a(s_163), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1692(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1693(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1694(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1625(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1626(.a(gate260inter0), .b(s_154), .O(gate260inter1));
  and2  gate1627(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1628(.a(s_154), .O(gate260inter3));
  inv1  gate1629(.a(s_155), .O(gate260inter4));
  nand2 gate1630(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1631(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1632(.a(G760), .O(gate260inter7));
  inv1  gate1633(.a(G761), .O(gate260inter8));
  nand2 gate1634(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1635(.a(s_155), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1636(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1637(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1638(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate855(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate856(.a(gate263inter0), .b(s_44), .O(gate263inter1));
  and2  gate857(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate858(.a(s_44), .O(gate263inter3));
  inv1  gate859(.a(s_45), .O(gate263inter4));
  nand2 gate860(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate861(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate862(.a(G766), .O(gate263inter7));
  inv1  gate863(.a(G767), .O(gate263inter8));
  nand2 gate864(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate865(.a(s_45), .b(gate263inter3), .O(gate263inter10));
  nor2  gate866(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate867(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate868(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1345(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1346(.a(gate265inter0), .b(s_114), .O(gate265inter1));
  and2  gate1347(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1348(.a(s_114), .O(gate265inter3));
  inv1  gate1349(.a(s_115), .O(gate265inter4));
  nand2 gate1350(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1351(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1352(.a(G642), .O(gate265inter7));
  inv1  gate1353(.a(G770), .O(gate265inter8));
  nand2 gate1354(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1355(.a(s_115), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1356(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1357(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1358(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate3011(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate3012(.a(gate273inter0), .b(s_352), .O(gate273inter1));
  and2  gate3013(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate3014(.a(s_352), .O(gate273inter3));
  inv1  gate3015(.a(s_353), .O(gate273inter4));
  nand2 gate3016(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate3017(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate3018(.a(G642), .O(gate273inter7));
  inv1  gate3019(.a(G794), .O(gate273inter8));
  nand2 gate3020(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate3021(.a(s_353), .b(gate273inter3), .O(gate273inter10));
  nor2  gate3022(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate3023(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate3024(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2955(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2956(.a(gate276inter0), .b(s_344), .O(gate276inter1));
  and2  gate2957(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2958(.a(s_344), .O(gate276inter3));
  inv1  gate2959(.a(s_345), .O(gate276inter4));
  nand2 gate2960(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2961(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2962(.a(G773), .O(gate276inter7));
  inv1  gate2963(.a(G797), .O(gate276inter8));
  nand2 gate2964(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2965(.a(s_345), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2966(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2967(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2968(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1401(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1402(.a(gate277inter0), .b(s_122), .O(gate277inter1));
  and2  gate1403(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1404(.a(s_122), .O(gate277inter3));
  inv1  gate1405(.a(s_123), .O(gate277inter4));
  nand2 gate1406(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1407(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1408(.a(G648), .O(gate277inter7));
  inv1  gate1409(.a(G800), .O(gate277inter8));
  nand2 gate1410(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1411(.a(s_123), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1412(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1413(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1414(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate2143(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2144(.a(gate278inter0), .b(s_228), .O(gate278inter1));
  and2  gate2145(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2146(.a(s_228), .O(gate278inter3));
  inv1  gate2147(.a(s_229), .O(gate278inter4));
  nand2 gate2148(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2149(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2150(.a(G776), .O(gate278inter7));
  inv1  gate2151(.a(G800), .O(gate278inter8));
  nand2 gate2152(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2153(.a(s_229), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2154(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2155(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2156(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate757(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate758(.a(gate282inter0), .b(s_30), .O(gate282inter1));
  and2  gate759(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate760(.a(s_30), .O(gate282inter3));
  inv1  gate761(.a(s_31), .O(gate282inter4));
  nand2 gate762(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate763(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate764(.a(G782), .O(gate282inter7));
  inv1  gate765(.a(G806), .O(gate282inter8));
  nand2 gate766(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate767(.a(s_31), .b(gate282inter3), .O(gate282inter10));
  nor2  gate768(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate769(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate770(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1191(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1192(.a(gate284inter0), .b(s_92), .O(gate284inter1));
  and2  gate1193(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1194(.a(s_92), .O(gate284inter3));
  inv1  gate1195(.a(s_93), .O(gate284inter4));
  nand2 gate1196(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1197(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1198(.a(G785), .O(gate284inter7));
  inv1  gate1199(.a(G809), .O(gate284inter8));
  nand2 gate1200(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1201(.a(s_93), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1202(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1203(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1204(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2521(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2522(.a(gate285inter0), .b(s_282), .O(gate285inter1));
  and2  gate2523(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2524(.a(s_282), .O(gate285inter3));
  inv1  gate2525(.a(s_283), .O(gate285inter4));
  nand2 gate2526(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2527(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2528(.a(G660), .O(gate285inter7));
  inv1  gate2529(.a(G812), .O(gate285inter8));
  nand2 gate2530(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2531(.a(s_283), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2532(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2533(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2534(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2843(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2844(.a(gate286inter0), .b(s_328), .O(gate286inter1));
  and2  gate2845(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2846(.a(s_328), .O(gate286inter3));
  inv1  gate2847(.a(s_329), .O(gate286inter4));
  nand2 gate2848(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2849(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2850(.a(G788), .O(gate286inter7));
  inv1  gate2851(.a(G812), .O(gate286inter8));
  nand2 gate2852(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2853(.a(s_329), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2854(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2855(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2856(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate589(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate590(.a(gate287inter0), .b(s_6), .O(gate287inter1));
  and2  gate591(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate592(.a(s_6), .O(gate287inter3));
  inv1  gate593(.a(s_7), .O(gate287inter4));
  nand2 gate594(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate595(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate596(.a(G663), .O(gate287inter7));
  inv1  gate597(.a(G815), .O(gate287inter8));
  nand2 gate598(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate599(.a(s_7), .b(gate287inter3), .O(gate287inter10));
  nor2  gate600(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate601(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate602(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate2633(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2634(.a(gate288inter0), .b(s_298), .O(gate288inter1));
  and2  gate2635(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2636(.a(s_298), .O(gate288inter3));
  inv1  gate2637(.a(s_299), .O(gate288inter4));
  nand2 gate2638(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2639(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2640(.a(G791), .O(gate288inter7));
  inv1  gate2641(.a(G815), .O(gate288inter8));
  nand2 gate2642(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2643(.a(s_299), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2644(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2645(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2646(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1289(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1290(.a(gate290inter0), .b(s_106), .O(gate290inter1));
  and2  gate1291(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1292(.a(s_106), .O(gate290inter3));
  inv1  gate1293(.a(s_107), .O(gate290inter4));
  nand2 gate1294(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1295(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1296(.a(G820), .O(gate290inter7));
  inv1  gate1297(.a(G821), .O(gate290inter8));
  nand2 gate1298(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1299(.a(s_107), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1300(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1301(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1302(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2283(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2284(.a(gate294inter0), .b(s_248), .O(gate294inter1));
  and2  gate2285(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2286(.a(s_248), .O(gate294inter3));
  inv1  gate2287(.a(s_249), .O(gate294inter4));
  nand2 gate2288(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2289(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2290(.a(G832), .O(gate294inter7));
  inv1  gate2291(.a(G833), .O(gate294inter8));
  nand2 gate2292(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2293(.a(s_249), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2294(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2295(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2296(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1275(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1276(.a(gate296inter0), .b(s_104), .O(gate296inter1));
  and2  gate1277(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1278(.a(s_104), .O(gate296inter3));
  inv1  gate1279(.a(s_105), .O(gate296inter4));
  nand2 gate1280(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1281(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1282(.a(G826), .O(gate296inter7));
  inv1  gate1283(.a(G827), .O(gate296inter8));
  nand2 gate1284(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1285(.a(s_105), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1286(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1287(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1288(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate673(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate674(.a(gate387inter0), .b(s_18), .O(gate387inter1));
  and2  gate675(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate676(.a(s_18), .O(gate387inter3));
  inv1  gate677(.a(s_19), .O(gate387inter4));
  nand2 gate678(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate679(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate680(.a(G1), .O(gate387inter7));
  inv1  gate681(.a(G1036), .O(gate387inter8));
  nand2 gate682(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate683(.a(s_19), .b(gate387inter3), .O(gate387inter10));
  nor2  gate684(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate685(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate686(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2297(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2298(.a(gate389inter0), .b(s_250), .O(gate389inter1));
  and2  gate2299(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2300(.a(s_250), .O(gate389inter3));
  inv1  gate2301(.a(s_251), .O(gate389inter4));
  nand2 gate2302(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2303(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2304(.a(G3), .O(gate389inter7));
  inv1  gate2305(.a(G1042), .O(gate389inter8));
  nand2 gate2306(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2307(.a(s_251), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2308(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2309(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2310(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2157(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2158(.a(gate391inter0), .b(s_230), .O(gate391inter1));
  and2  gate2159(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2160(.a(s_230), .O(gate391inter3));
  inv1  gate2161(.a(s_231), .O(gate391inter4));
  nand2 gate2162(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2163(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2164(.a(G5), .O(gate391inter7));
  inv1  gate2165(.a(G1048), .O(gate391inter8));
  nand2 gate2166(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2167(.a(s_231), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2168(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2169(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2170(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate3095(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate3096(.a(gate396inter0), .b(s_364), .O(gate396inter1));
  and2  gate3097(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate3098(.a(s_364), .O(gate396inter3));
  inv1  gate3099(.a(s_365), .O(gate396inter4));
  nand2 gate3100(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate3101(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate3102(.a(G10), .O(gate396inter7));
  inv1  gate3103(.a(G1063), .O(gate396inter8));
  nand2 gate3104(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate3105(.a(s_365), .b(gate396inter3), .O(gate396inter10));
  nor2  gate3106(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate3107(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate3108(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2451(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2452(.a(gate398inter0), .b(s_272), .O(gate398inter1));
  and2  gate2453(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2454(.a(s_272), .O(gate398inter3));
  inv1  gate2455(.a(s_273), .O(gate398inter4));
  nand2 gate2456(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2457(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2458(.a(G12), .O(gate398inter7));
  inv1  gate2459(.a(G1069), .O(gate398inter8));
  nand2 gate2460(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2461(.a(s_273), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2462(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2463(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2464(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1485(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1486(.a(gate399inter0), .b(s_134), .O(gate399inter1));
  and2  gate1487(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1488(.a(s_134), .O(gate399inter3));
  inv1  gate1489(.a(s_135), .O(gate399inter4));
  nand2 gate1490(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1491(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1492(.a(G13), .O(gate399inter7));
  inv1  gate1493(.a(G1072), .O(gate399inter8));
  nand2 gate1494(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1495(.a(s_135), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1496(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1497(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1498(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1499(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1500(.a(gate401inter0), .b(s_136), .O(gate401inter1));
  and2  gate1501(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1502(.a(s_136), .O(gate401inter3));
  inv1  gate1503(.a(s_137), .O(gate401inter4));
  nand2 gate1504(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1505(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1506(.a(G15), .O(gate401inter7));
  inv1  gate1507(.a(G1078), .O(gate401inter8));
  nand2 gate1508(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1509(.a(s_137), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1510(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1511(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1512(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1905(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1906(.a(gate405inter0), .b(s_194), .O(gate405inter1));
  and2  gate1907(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1908(.a(s_194), .O(gate405inter3));
  inv1  gate1909(.a(s_195), .O(gate405inter4));
  nand2 gate1910(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1911(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1912(.a(G19), .O(gate405inter7));
  inv1  gate1913(.a(G1090), .O(gate405inter8));
  nand2 gate1914(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1915(.a(s_195), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1916(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1917(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1918(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1023(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1024(.a(gate406inter0), .b(s_68), .O(gate406inter1));
  and2  gate1025(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1026(.a(s_68), .O(gate406inter3));
  inv1  gate1027(.a(s_69), .O(gate406inter4));
  nand2 gate1028(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1029(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1030(.a(G20), .O(gate406inter7));
  inv1  gate1031(.a(G1093), .O(gate406inter8));
  nand2 gate1032(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1033(.a(s_69), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1034(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1035(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1036(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1331(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1332(.a(gate409inter0), .b(s_112), .O(gate409inter1));
  and2  gate1333(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1334(.a(s_112), .O(gate409inter3));
  inv1  gate1335(.a(s_113), .O(gate409inter4));
  nand2 gate1336(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1337(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1338(.a(G23), .O(gate409inter7));
  inv1  gate1339(.a(G1102), .O(gate409inter8));
  nand2 gate1340(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1341(.a(s_113), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1342(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1343(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1344(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1597(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1598(.a(gate413inter0), .b(s_150), .O(gate413inter1));
  and2  gate1599(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1600(.a(s_150), .O(gate413inter3));
  inv1  gate1601(.a(s_151), .O(gate413inter4));
  nand2 gate1602(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1603(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1604(.a(G27), .O(gate413inter7));
  inv1  gate1605(.a(G1114), .O(gate413inter8));
  nand2 gate1606(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1607(.a(s_151), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1608(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1609(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1610(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2129(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2130(.a(gate415inter0), .b(s_226), .O(gate415inter1));
  and2  gate2131(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2132(.a(s_226), .O(gate415inter3));
  inv1  gate2133(.a(s_227), .O(gate415inter4));
  nand2 gate2134(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2135(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2136(.a(G29), .O(gate415inter7));
  inv1  gate2137(.a(G1120), .O(gate415inter8));
  nand2 gate2138(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2139(.a(s_227), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2140(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2141(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2142(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1877(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1878(.a(gate416inter0), .b(s_190), .O(gate416inter1));
  and2  gate1879(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1880(.a(s_190), .O(gate416inter3));
  inv1  gate1881(.a(s_191), .O(gate416inter4));
  nand2 gate1882(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1883(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1884(.a(G30), .O(gate416inter7));
  inv1  gate1885(.a(G1123), .O(gate416inter8));
  nand2 gate1886(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1887(.a(s_191), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1888(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1889(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1890(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate3025(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate3026(.a(gate418inter0), .b(s_354), .O(gate418inter1));
  and2  gate3027(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate3028(.a(s_354), .O(gate418inter3));
  inv1  gate3029(.a(s_355), .O(gate418inter4));
  nand2 gate3030(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate3031(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate3032(.a(G32), .O(gate418inter7));
  inv1  gate3033(.a(G1129), .O(gate418inter8));
  nand2 gate3034(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate3035(.a(s_355), .b(gate418inter3), .O(gate418inter10));
  nor2  gate3036(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate3037(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate3038(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2423(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2424(.a(gate419inter0), .b(s_268), .O(gate419inter1));
  and2  gate2425(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2426(.a(s_268), .O(gate419inter3));
  inv1  gate2427(.a(s_269), .O(gate419inter4));
  nand2 gate2428(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2429(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2430(.a(G1), .O(gate419inter7));
  inv1  gate2431(.a(G1132), .O(gate419inter8));
  nand2 gate2432(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2433(.a(s_269), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2434(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2435(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2436(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1583(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1584(.a(gate420inter0), .b(s_148), .O(gate420inter1));
  and2  gate1585(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1586(.a(s_148), .O(gate420inter3));
  inv1  gate1587(.a(s_149), .O(gate420inter4));
  nand2 gate1588(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1589(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1590(.a(G1036), .O(gate420inter7));
  inv1  gate1591(.a(G1132), .O(gate420inter8));
  nand2 gate1592(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1593(.a(s_149), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1594(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1595(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1596(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1947(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1948(.a(gate423inter0), .b(s_200), .O(gate423inter1));
  and2  gate1949(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1950(.a(s_200), .O(gate423inter3));
  inv1  gate1951(.a(s_201), .O(gate423inter4));
  nand2 gate1952(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1953(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1954(.a(G3), .O(gate423inter7));
  inv1  gate1955(.a(G1138), .O(gate423inter8));
  nand2 gate1956(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1957(.a(s_201), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1958(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1959(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1960(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1653(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1654(.a(gate426inter0), .b(s_158), .O(gate426inter1));
  and2  gate1655(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1656(.a(s_158), .O(gate426inter3));
  inv1  gate1657(.a(s_159), .O(gate426inter4));
  nand2 gate1658(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1659(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1660(.a(G1045), .O(gate426inter7));
  inv1  gate1661(.a(G1141), .O(gate426inter8));
  nand2 gate1662(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1663(.a(s_159), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1664(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1665(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1666(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2941(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2942(.a(gate427inter0), .b(s_342), .O(gate427inter1));
  and2  gate2943(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2944(.a(s_342), .O(gate427inter3));
  inv1  gate2945(.a(s_343), .O(gate427inter4));
  nand2 gate2946(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2947(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2948(.a(G5), .O(gate427inter7));
  inv1  gate2949(.a(G1144), .O(gate427inter8));
  nand2 gate2950(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2951(.a(s_343), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2952(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2953(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2954(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1037(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1038(.a(gate428inter0), .b(s_70), .O(gate428inter1));
  and2  gate1039(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1040(.a(s_70), .O(gate428inter3));
  inv1  gate1041(.a(s_71), .O(gate428inter4));
  nand2 gate1042(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1043(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1044(.a(G1048), .O(gate428inter7));
  inv1  gate1045(.a(G1144), .O(gate428inter8));
  nand2 gate1046(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1047(.a(s_71), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1048(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1049(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1050(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate939(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate940(.a(gate429inter0), .b(s_56), .O(gate429inter1));
  and2  gate941(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate942(.a(s_56), .O(gate429inter3));
  inv1  gate943(.a(s_57), .O(gate429inter4));
  nand2 gate944(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate945(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate946(.a(G6), .O(gate429inter7));
  inv1  gate947(.a(G1147), .O(gate429inter8));
  nand2 gate948(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate949(.a(s_57), .b(gate429inter3), .O(gate429inter10));
  nor2  gate950(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate951(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate952(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate2017(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2018(.a(gate430inter0), .b(s_210), .O(gate430inter1));
  and2  gate2019(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2020(.a(s_210), .O(gate430inter3));
  inv1  gate2021(.a(s_211), .O(gate430inter4));
  nand2 gate2022(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2023(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2024(.a(G1051), .O(gate430inter7));
  inv1  gate2025(.a(G1147), .O(gate430inter8));
  nand2 gate2026(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2027(.a(s_211), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2028(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2029(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2030(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1373(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1374(.a(gate431inter0), .b(s_118), .O(gate431inter1));
  and2  gate1375(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1376(.a(s_118), .O(gate431inter3));
  inv1  gate1377(.a(s_119), .O(gate431inter4));
  nand2 gate1378(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1379(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1380(.a(G7), .O(gate431inter7));
  inv1  gate1381(.a(G1150), .O(gate431inter8));
  nand2 gate1382(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1383(.a(s_119), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1384(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1385(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1386(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate799(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate800(.a(gate433inter0), .b(s_36), .O(gate433inter1));
  and2  gate801(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate802(.a(s_36), .O(gate433inter3));
  inv1  gate803(.a(s_37), .O(gate433inter4));
  nand2 gate804(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate805(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate806(.a(G8), .O(gate433inter7));
  inv1  gate807(.a(G1153), .O(gate433inter8));
  nand2 gate808(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate809(.a(s_37), .b(gate433inter3), .O(gate433inter10));
  nor2  gate810(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate811(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate812(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate2535(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2536(.a(gate434inter0), .b(s_284), .O(gate434inter1));
  and2  gate2537(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2538(.a(s_284), .O(gate434inter3));
  inv1  gate2539(.a(s_285), .O(gate434inter4));
  nand2 gate2540(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2541(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2542(.a(G1057), .O(gate434inter7));
  inv1  gate2543(.a(G1153), .O(gate434inter8));
  nand2 gate2544(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2545(.a(s_285), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2546(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2547(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2548(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2899(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2900(.a(gate435inter0), .b(s_336), .O(gate435inter1));
  and2  gate2901(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2902(.a(s_336), .O(gate435inter3));
  inv1  gate2903(.a(s_337), .O(gate435inter4));
  nand2 gate2904(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2905(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2906(.a(G9), .O(gate435inter7));
  inv1  gate2907(.a(G1156), .O(gate435inter8));
  nand2 gate2908(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2909(.a(s_337), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2910(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2911(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2912(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1527(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1528(.a(gate440inter0), .b(s_140), .O(gate440inter1));
  and2  gate1529(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1530(.a(s_140), .O(gate440inter3));
  inv1  gate1531(.a(s_141), .O(gate440inter4));
  nand2 gate1532(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1533(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1534(.a(G1066), .O(gate440inter7));
  inv1  gate1535(.a(G1162), .O(gate440inter8));
  nand2 gate1536(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1537(.a(s_141), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1538(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1539(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1540(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate2171(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2172(.a(gate441inter0), .b(s_232), .O(gate441inter1));
  and2  gate2173(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2174(.a(s_232), .O(gate441inter3));
  inv1  gate2175(.a(s_233), .O(gate441inter4));
  nand2 gate2176(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2177(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2178(.a(G12), .O(gate441inter7));
  inv1  gate2179(.a(G1165), .O(gate441inter8));
  nand2 gate2180(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2181(.a(s_233), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2182(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2183(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2184(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate897(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate898(.a(gate442inter0), .b(s_50), .O(gate442inter1));
  and2  gate899(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate900(.a(s_50), .O(gate442inter3));
  inv1  gate901(.a(s_51), .O(gate442inter4));
  nand2 gate902(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate903(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate904(.a(G1069), .O(gate442inter7));
  inv1  gate905(.a(G1165), .O(gate442inter8));
  nand2 gate906(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate907(.a(s_51), .b(gate442inter3), .O(gate442inter10));
  nor2  gate908(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate909(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate910(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1135(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1136(.a(gate443inter0), .b(s_84), .O(gate443inter1));
  and2  gate1137(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1138(.a(s_84), .O(gate443inter3));
  inv1  gate1139(.a(s_85), .O(gate443inter4));
  nand2 gate1140(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1141(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1142(.a(G13), .O(gate443inter7));
  inv1  gate1143(.a(G1168), .O(gate443inter8));
  nand2 gate1144(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1145(.a(s_85), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1146(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1147(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1148(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate3067(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate3068(.a(gate444inter0), .b(s_360), .O(gate444inter1));
  and2  gate3069(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate3070(.a(s_360), .O(gate444inter3));
  inv1  gate3071(.a(s_361), .O(gate444inter4));
  nand2 gate3072(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate3073(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate3074(.a(G1072), .O(gate444inter7));
  inv1  gate3075(.a(G1168), .O(gate444inter8));
  nand2 gate3076(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate3077(.a(s_361), .b(gate444inter3), .O(gate444inter10));
  nor2  gate3078(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate3079(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate3080(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1961(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1962(.a(gate451inter0), .b(s_202), .O(gate451inter1));
  and2  gate1963(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1964(.a(s_202), .O(gate451inter3));
  inv1  gate1965(.a(s_203), .O(gate451inter4));
  nand2 gate1966(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1967(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1968(.a(G17), .O(gate451inter7));
  inv1  gate1969(.a(G1180), .O(gate451inter8));
  nand2 gate1970(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1971(.a(s_203), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1972(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1973(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1974(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate883(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate884(.a(gate452inter0), .b(s_48), .O(gate452inter1));
  and2  gate885(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate886(.a(s_48), .O(gate452inter3));
  inv1  gate887(.a(s_49), .O(gate452inter4));
  nand2 gate888(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate889(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate890(.a(G1084), .O(gate452inter7));
  inv1  gate891(.a(G1180), .O(gate452inter8));
  nand2 gate892(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate893(.a(s_49), .b(gate452inter3), .O(gate452inter10));
  nor2  gate894(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate895(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate896(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate3193(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate3194(.a(gate453inter0), .b(s_378), .O(gate453inter1));
  and2  gate3195(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate3196(.a(s_378), .O(gate453inter3));
  inv1  gate3197(.a(s_379), .O(gate453inter4));
  nand2 gate3198(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate3199(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate3200(.a(G18), .O(gate453inter7));
  inv1  gate3201(.a(G1183), .O(gate453inter8));
  nand2 gate3202(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate3203(.a(s_379), .b(gate453inter3), .O(gate453inter10));
  nor2  gate3204(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate3205(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate3206(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate2549(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2550(.a(gate454inter0), .b(s_286), .O(gate454inter1));
  and2  gate2551(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2552(.a(s_286), .O(gate454inter3));
  inv1  gate2553(.a(s_287), .O(gate454inter4));
  nand2 gate2554(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2555(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2556(.a(G1087), .O(gate454inter7));
  inv1  gate2557(.a(G1183), .O(gate454inter8));
  nand2 gate2558(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2559(.a(s_287), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2560(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2561(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2562(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate631(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate632(.a(gate458inter0), .b(s_12), .O(gate458inter1));
  and2  gate633(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate634(.a(s_12), .O(gate458inter3));
  inv1  gate635(.a(s_13), .O(gate458inter4));
  nand2 gate636(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate637(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate638(.a(G1093), .O(gate458inter7));
  inv1  gate639(.a(G1189), .O(gate458inter8));
  nand2 gate640(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate641(.a(s_13), .b(gate458inter3), .O(gate458inter10));
  nor2  gate642(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate643(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate644(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2353(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2354(.a(gate460inter0), .b(s_258), .O(gate460inter1));
  and2  gate2355(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2356(.a(s_258), .O(gate460inter3));
  inv1  gate2357(.a(s_259), .O(gate460inter4));
  nand2 gate2358(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2359(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2360(.a(G1096), .O(gate460inter7));
  inv1  gate2361(.a(G1192), .O(gate460inter8));
  nand2 gate2362(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2363(.a(s_259), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2364(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2365(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2366(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate3039(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate3040(.a(gate463inter0), .b(s_356), .O(gate463inter1));
  and2  gate3041(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate3042(.a(s_356), .O(gate463inter3));
  inv1  gate3043(.a(s_357), .O(gate463inter4));
  nand2 gate3044(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate3045(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate3046(.a(G23), .O(gate463inter7));
  inv1  gate3047(.a(G1198), .O(gate463inter8));
  nand2 gate3048(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate3049(.a(s_357), .b(gate463inter3), .O(gate463inter10));
  nor2  gate3050(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate3051(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate3052(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2619(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2620(.a(gate465inter0), .b(s_296), .O(gate465inter1));
  and2  gate2621(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2622(.a(s_296), .O(gate465inter3));
  inv1  gate2623(.a(s_297), .O(gate465inter4));
  nand2 gate2624(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2625(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2626(.a(G24), .O(gate465inter7));
  inv1  gate2627(.a(G1201), .O(gate465inter8));
  nand2 gate2628(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2629(.a(s_297), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2630(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2631(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2632(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1303(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1304(.a(gate469inter0), .b(s_108), .O(gate469inter1));
  and2  gate1305(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1306(.a(s_108), .O(gate469inter3));
  inv1  gate1307(.a(s_109), .O(gate469inter4));
  nand2 gate1308(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1309(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1310(.a(G26), .O(gate469inter7));
  inv1  gate1311(.a(G1207), .O(gate469inter8));
  nand2 gate1312(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1313(.a(s_109), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1314(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1315(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1316(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2185(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2186(.a(gate470inter0), .b(s_234), .O(gate470inter1));
  and2  gate2187(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2188(.a(s_234), .O(gate470inter3));
  inv1  gate2189(.a(s_235), .O(gate470inter4));
  nand2 gate2190(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2191(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2192(.a(G1111), .O(gate470inter7));
  inv1  gate2193(.a(G1207), .O(gate470inter8));
  nand2 gate2194(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2195(.a(s_235), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2196(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2197(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2198(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1443(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1444(.a(gate473inter0), .b(s_128), .O(gate473inter1));
  and2  gate1445(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1446(.a(s_128), .O(gate473inter3));
  inv1  gate1447(.a(s_129), .O(gate473inter4));
  nand2 gate1448(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1449(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1450(.a(G28), .O(gate473inter7));
  inv1  gate1451(.a(G1213), .O(gate473inter8));
  nand2 gate1452(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1453(.a(s_129), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1454(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1455(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1456(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2339(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2340(.a(gate482inter0), .b(s_256), .O(gate482inter1));
  and2  gate2341(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2342(.a(s_256), .O(gate482inter3));
  inv1  gate2343(.a(s_257), .O(gate482inter4));
  nand2 gate2344(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2345(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2346(.a(G1129), .O(gate482inter7));
  inv1  gate2347(.a(G1225), .O(gate482inter8));
  nand2 gate2348(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2349(.a(s_257), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2350(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2351(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2352(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1359(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1360(.a(gate486inter0), .b(s_116), .O(gate486inter1));
  and2  gate1361(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1362(.a(s_116), .O(gate486inter3));
  inv1  gate1363(.a(s_117), .O(gate486inter4));
  nand2 gate1364(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1365(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1366(.a(G1234), .O(gate486inter7));
  inv1  gate1367(.a(G1235), .O(gate486inter8));
  nand2 gate1368(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1369(.a(s_117), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1370(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1371(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1372(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1695(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1696(.a(gate487inter0), .b(s_164), .O(gate487inter1));
  and2  gate1697(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1698(.a(s_164), .O(gate487inter3));
  inv1  gate1699(.a(s_165), .O(gate487inter4));
  nand2 gate1700(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1701(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1702(.a(G1236), .O(gate487inter7));
  inv1  gate1703(.a(G1237), .O(gate487inter8));
  nand2 gate1704(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1705(.a(s_165), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1706(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1707(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1708(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2871(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2872(.a(gate488inter0), .b(s_332), .O(gate488inter1));
  and2  gate2873(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2874(.a(s_332), .O(gate488inter3));
  inv1  gate2875(.a(s_333), .O(gate488inter4));
  nand2 gate2876(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2877(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2878(.a(G1238), .O(gate488inter7));
  inv1  gate2879(.a(G1239), .O(gate488inter8));
  nand2 gate2880(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2881(.a(s_333), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2882(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2883(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2884(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate2591(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2592(.a(gate489inter0), .b(s_292), .O(gate489inter1));
  and2  gate2593(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2594(.a(s_292), .O(gate489inter3));
  inv1  gate2595(.a(s_293), .O(gate489inter4));
  nand2 gate2596(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2597(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2598(.a(G1240), .O(gate489inter7));
  inv1  gate2599(.a(G1241), .O(gate489inter8));
  nand2 gate2600(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2601(.a(s_293), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2602(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2603(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2604(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate2829(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2830(.a(gate490inter0), .b(s_326), .O(gate490inter1));
  and2  gate2831(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2832(.a(s_326), .O(gate490inter3));
  inv1  gate2833(.a(s_327), .O(gate490inter4));
  nand2 gate2834(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2835(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2836(.a(G1242), .O(gate490inter7));
  inv1  gate2837(.a(G1243), .O(gate490inter8));
  nand2 gate2838(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2839(.a(s_327), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2840(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2841(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2842(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1205(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1206(.a(gate491inter0), .b(s_94), .O(gate491inter1));
  and2  gate1207(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1208(.a(s_94), .O(gate491inter3));
  inv1  gate1209(.a(s_95), .O(gate491inter4));
  nand2 gate1210(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1211(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1212(.a(G1244), .O(gate491inter7));
  inv1  gate1213(.a(G1245), .O(gate491inter8));
  nand2 gate1214(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1215(.a(s_95), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1216(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1217(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1218(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1429(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1430(.a(gate492inter0), .b(s_126), .O(gate492inter1));
  and2  gate1431(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1432(.a(s_126), .O(gate492inter3));
  inv1  gate1433(.a(s_127), .O(gate492inter4));
  nand2 gate1434(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1435(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1436(.a(G1246), .O(gate492inter7));
  inv1  gate1437(.a(G1247), .O(gate492inter8));
  nand2 gate1438(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1439(.a(s_127), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1440(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1441(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1442(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1667(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1668(.a(gate493inter0), .b(s_160), .O(gate493inter1));
  and2  gate1669(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1670(.a(s_160), .O(gate493inter3));
  inv1  gate1671(.a(s_161), .O(gate493inter4));
  nand2 gate1672(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1673(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1674(.a(G1248), .O(gate493inter7));
  inv1  gate1675(.a(G1249), .O(gate493inter8));
  nand2 gate1676(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1677(.a(s_161), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1678(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1679(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1680(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2759(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2760(.a(gate494inter0), .b(s_316), .O(gate494inter1));
  and2  gate2761(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2762(.a(s_316), .O(gate494inter3));
  inv1  gate2763(.a(s_317), .O(gate494inter4));
  nand2 gate2764(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2765(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2766(.a(G1250), .O(gate494inter7));
  inv1  gate2767(.a(G1251), .O(gate494inter8));
  nand2 gate2768(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2769(.a(s_317), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2770(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2771(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2772(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2731(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2732(.a(gate497inter0), .b(s_312), .O(gate497inter1));
  and2  gate2733(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2734(.a(s_312), .O(gate497inter3));
  inv1  gate2735(.a(s_313), .O(gate497inter4));
  nand2 gate2736(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2737(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2738(.a(G1256), .O(gate497inter7));
  inv1  gate2739(.a(G1257), .O(gate497inter8));
  nand2 gate2740(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2741(.a(s_313), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2742(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2743(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2744(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2605(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2606(.a(gate499inter0), .b(s_294), .O(gate499inter1));
  and2  gate2607(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2608(.a(s_294), .O(gate499inter3));
  inv1  gate2609(.a(s_295), .O(gate499inter4));
  nand2 gate2610(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2611(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2612(.a(G1260), .O(gate499inter7));
  inv1  gate2613(.a(G1261), .O(gate499inter8));
  nand2 gate2614(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2615(.a(s_295), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2616(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2617(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2618(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate687(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate688(.a(gate500inter0), .b(s_20), .O(gate500inter1));
  and2  gate689(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate690(.a(s_20), .O(gate500inter3));
  inv1  gate691(.a(s_21), .O(gate500inter4));
  nand2 gate692(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate693(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate694(.a(G1262), .O(gate500inter7));
  inv1  gate695(.a(G1263), .O(gate500inter8));
  nand2 gate696(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate697(.a(s_21), .b(gate500inter3), .O(gate500inter10));
  nor2  gate698(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate699(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate700(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2325(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2326(.a(gate503inter0), .b(s_254), .O(gate503inter1));
  and2  gate2327(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2328(.a(s_254), .O(gate503inter3));
  inv1  gate2329(.a(s_255), .O(gate503inter4));
  nand2 gate2330(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2331(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2332(.a(G1268), .O(gate503inter7));
  inv1  gate2333(.a(G1269), .O(gate503inter8));
  nand2 gate2334(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2335(.a(s_255), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2336(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2337(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2338(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate603(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate604(.a(gate505inter0), .b(s_8), .O(gate505inter1));
  and2  gate605(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate606(.a(s_8), .O(gate505inter3));
  inv1  gate607(.a(s_9), .O(gate505inter4));
  nand2 gate608(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate609(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate610(.a(G1272), .O(gate505inter7));
  inv1  gate611(.a(G1273), .O(gate505inter8));
  nand2 gate612(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate613(.a(s_9), .b(gate505inter3), .O(gate505inter10));
  nor2  gate614(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate615(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate616(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2031(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2032(.a(gate511inter0), .b(s_212), .O(gate511inter1));
  and2  gate2033(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2034(.a(s_212), .O(gate511inter3));
  inv1  gate2035(.a(s_213), .O(gate511inter4));
  nand2 gate2036(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2037(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2038(.a(G1284), .O(gate511inter7));
  inv1  gate2039(.a(G1285), .O(gate511inter8));
  nand2 gate2040(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2041(.a(s_213), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2042(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2043(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2044(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1569(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1570(.a(gate512inter0), .b(s_146), .O(gate512inter1));
  and2  gate1571(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1572(.a(s_146), .O(gate512inter3));
  inv1  gate1573(.a(s_147), .O(gate512inter4));
  nand2 gate1574(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1575(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1576(.a(G1286), .O(gate512inter7));
  inv1  gate1577(.a(G1287), .O(gate512inter8));
  nand2 gate1578(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1579(.a(s_147), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1580(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1581(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1582(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate743(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate744(.a(gate513inter0), .b(s_28), .O(gate513inter1));
  and2  gate745(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate746(.a(s_28), .O(gate513inter3));
  inv1  gate747(.a(s_29), .O(gate513inter4));
  nand2 gate748(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate749(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate750(.a(G1288), .O(gate513inter7));
  inv1  gate751(.a(G1289), .O(gate513inter8));
  nand2 gate752(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate753(.a(s_29), .b(gate513inter3), .O(gate513inter10));
  nor2  gate754(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate755(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate756(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate2969(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2970(.a(gate514inter0), .b(s_346), .O(gate514inter1));
  and2  gate2971(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2972(.a(s_346), .O(gate514inter3));
  inv1  gate2973(.a(s_347), .O(gate514inter4));
  nand2 gate2974(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2975(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2976(.a(G1290), .O(gate514inter7));
  inv1  gate2977(.a(G1291), .O(gate514inter8));
  nand2 gate2978(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2979(.a(s_347), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2980(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2981(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2982(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule