module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1163(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1164(.a(gate9inter0), .b(s_88), .O(gate9inter1));
  and2  gate1165(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1166(.a(s_88), .O(gate9inter3));
  inv1  gate1167(.a(s_89), .O(gate9inter4));
  nand2 gate1168(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1169(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1170(.a(G1), .O(gate9inter7));
  inv1  gate1171(.a(G2), .O(gate9inter8));
  nand2 gate1172(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1173(.a(s_89), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1174(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1175(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1176(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate589(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate590(.a(gate12inter0), .b(s_6), .O(gate12inter1));
  and2  gate591(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate592(.a(s_6), .O(gate12inter3));
  inv1  gate593(.a(s_7), .O(gate12inter4));
  nand2 gate594(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate595(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate596(.a(G7), .O(gate12inter7));
  inv1  gate597(.a(G8), .O(gate12inter8));
  nand2 gate598(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate599(.a(s_7), .b(gate12inter3), .O(gate12inter10));
  nor2  gate600(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate601(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate602(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1303(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1304(.a(gate21inter0), .b(s_108), .O(gate21inter1));
  and2  gate1305(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1306(.a(s_108), .O(gate21inter3));
  inv1  gate1307(.a(s_109), .O(gate21inter4));
  nand2 gate1308(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1309(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1310(.a(G25), .O(gate21inter7));
  inv1  gate1311(.a(G26), .O(gate21inter8));
  nand2 gate1312(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1313(.a(s_109), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1314(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1315(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1316(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate757(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate758(.a(gate28inter0), .b(s_30), .O(gate28inter1));
  and2  gate759(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate760(.a(s_30), .O(gate28inter3));
  inv1  gate761(.a(s_31), .O(gate28inter4));
  nand2 gate762(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate763(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate764(.a(G10), .O(gate28inter7));
  inv1  gate765(.a(G14), .O(gate28inter8));
  nand2 gate766(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate767(.a(s_31), .b(gate28inter3), .O(gate28inter10));
  nor2  gate768(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate769(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate770(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1611(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1612(.a(gate30inter0), .b(s_152), .O(gate30inter1));
  and2  gate1613(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1614(.a(s_152), .O(gate30inter3));
  inv1  gate1615(.a(s_153), .O(gate30inter4));
  nand2 gate1616(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1617(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1618(.a(G11), .O(gate30inter7));
  inv1  gate1619(.a(G15), .O(gate30inter8));
  nand2 gate1620(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1621(.a(s_153), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1622(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1623(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1624(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1541(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1542(.a(gate34inter0), .b(s_142), .O(gate34inter1));
  and2  gate1543(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1544(.a(s_142), .O(gate34inter3));
  inv1  gate1545(.a(s_143), .O(gate34inter4));
  nand2 gate1546(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1547(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1548(.a(G25), .O(gate34inter7));
  inv1  gate1549(.a(G29), .O(gate34inter8));
  nand2 gate1550(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1551(.a(s_143), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1552(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1553(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1554(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate813(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate814(.a(gate43inter0), .b(s_38), .O(gate43inter1));
  and2  gate815(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate816(.a(s_38), .O(gate43inter3));
  inv1  gate817(.a(s_39), .O(gate43inter4));
  nand2 gate818(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate819(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate820(.a(G3), .O(gate43inter7));
  inv1  gate821(.a(G269), .O(gate43inter8));
  nand2 gate822(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate823(.a(s_39), .b(gate43inter3), .O(gate43inter10));
  nor2  gate824(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate825(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate826(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1233(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1234(.a(gate50inter0), .b(s_98), .O(gate50inter1));
  and2  gate1235(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1236(.a(s_98), .O(gate50inter3));
  inv1  gate1237(.a(s_99), .O(gate50inter4));
  nand2 gate1238(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1239(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1240(.a(G10), .O(gate50inter7));
  inv1  gate1241(.a(G278), .O(gate50inter8));
  nand2 gate1242(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1243(.a(s_99), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1244(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1245(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1246(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2157(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2158(.a(gate53inter0), .b(s_230), .O(gate53inter1));
  and2  gate2159(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2160(.a(s_230), .O(gate53inter3));
  inv1  gate2161(.a(s_231), .O(gate53inter4));
  nand2 gate2162(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2163(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2164(.a(G13), .O(gate53inter7));
  inv1  gate2165(.a(G284), .O(gate53inter8));
  nand2 gate2166(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2167(.a(s_231), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2168(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2169(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2170(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1275(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1276(.a(gate54inter0), .b(s_104), .O(gate54inter1));
  and2  gate1277(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1278(.a(s_104), .O(gate54inter3));
  inv1  gate1279(.a(s_105), .O(gate54inter4));
  nand2 gate1280(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1281(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1282(.a(G14), .O(gate54inter7));
  inv1  gate1283(.a(G284), .O(gate54inter8));
  nand2 gate1284(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1285(.a(s_105), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1286(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1287(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1288(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1877(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1878(.a(gate56inter0), .b(s_190), .O(gate56inter1));
  and2  gate1879(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1880(.a(s_190), .O(gate56inter3));
  inv1  gate1881(.a(s_191), .O(gate56inter4));
  nand2 gate1882(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1883(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1884(.a(G16), .O(gate56inter7));
  inv1  gate1885(.a(G287), .O(gate56inter8));
  nand2 gate1886(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1887(.a(s_191), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1888(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1889(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1890(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate967(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate968(.a(gate59inter0), .b(s_60), .O(gate59inter1));
  and2  gate969(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate970(.a(s_60), .O(gate59inter3));
  inv1  gate971(.a(s_61), .O(gate59inter4));
  nand2 gate972(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate973(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate974(.a(G19), .O(gate59inter7));
  inv1  gate975(.a(G293), .O(gate59inter8));
  nand2 gate976(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate977(.a(s_61), .b(gate59inter3), .O(gate59inter10));
  nor2  gate978(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate979(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate980(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1849(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1850(.a(gate60inter0), .b(s_186), .O(gate60inter1));
  and2  gate1851(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1852(.a(s_186), .O(gate60inter3));
  inv1  gate1853(.a(s_187), .O(gate60inter4));
  nand2 gate1854(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1855(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1856(.a(G20), .O(gate60inter7));
  inv1  gate1857(.a(G293), .O(gate60inter8));
  nand2 gate1858(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1859(.a(s_187), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1860(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1861(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1862(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1793(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1794(.a(gate72inter0), .b(s_178), .O(gate72inter1));
  and2  gate1795(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1796(.a(s_178), .O(gate72inter3));
  inv1  gate1797(.a(s_179), .O(gate72inter4));
  nand2 gate1798(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1799(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1800(.a(G32), .O(gate72inter7));
  inv1  gate1801(.a(G311), .O(gate72inter8));
  nand2 gate1802(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1803(.a(s_179), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1804(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1805(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1806(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate2115(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2116(.a(gate73inter0), .b(s_224), .O(gate73inter1));
  and2  gate2117(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2118(.a(s_224), .O(gate73inter3));
  inv1  gate2119(.a(s_225), .O(gate73inter4));
  nand2 gate2120(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2121(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2122(.a(G1), .O(gate73inter7));
  inv1  gate2123(.a(G314), .O(gate73inter8));
  nand2 gate2124(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2125(.a(s_225), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2126(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2127(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2128(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate659(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate660(.a(gate74inter0), .b(s_16), .O(gate74inter1));
  and2  gate661(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate662(.a(s_16), .O(gate74inter3));
  inv1  gate663(.a(s_17), .O(gate74inter4));
  nand2 gate664(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate665(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate666(.a(G5), .O(gate74inter7));
  inv1  gate667(.a(G314), .O(gate74inter8));
  nand2 gate668(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate669(.a(s_17), .b(gate74inter3), .O(gate74inter10));
  nor2  gate670(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate671(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate672(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1947(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1948(.a(gate75inter0), .b(s_200), .O(gate75inter1));
  and2  gate1949(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1950(.a(s_200), .O(gate75inter3));
  inv1  gate1951(.a(s_201), .O(gate75inter4));
  nand2 gate1952(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1953(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1954(.a(G9), .O(gate75inter7));
  inv1  gate1955(.a(G317), .O(gate75inter8));
  nand2 gate1956(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1957(.a(s_201), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1958(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1959(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1960(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1387(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1388(.a(gate76inter0), .b(s_120), .O(gate76inter1));
  and2  gate1389(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1390(.a(s_120), .O(gate76inter3));
  inv1  gate1391(.a(s_121), .O(gate76inter4));
  nand2 gate1392(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1393(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1394(.a(G13), .O(gate76inter7));
  inv1  gate1395(.a(G317), .O(gate76inter8));
  nand2 gate1396(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1397(.a(s_121), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1398(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1399(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1400(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate827(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate828(.a(gate79inter0), .b(s_40), .O(gate79inter1));
  and2  gate829(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate830(.a(s_40), .O(gate79inter3));
  inv1  gate831(.a(s_41), .O(gate79inter4));
  nand2 gate832(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate833(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate834(.a(G10), .O(gate79inter7));
  inv1  gate835(.a(G323), .O(gate79inter8));
  nand2 gate836(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate837(.a(s_41), .b(gate79inter3), .O(gate79inter10));
  nor2  gate838(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate839(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate840(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1863(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1864(.a(gate83inter0), .b(s_188), .O(gate83inter1));
  and2  gate1865(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1866(.a(s_188), .O(gate83inter3));
  inv1  gate1867(.a(s_189), .O(gate83inter4));
  nand2 gate1868(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1869(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1870(.a(G11), .O(gate83inter7));
  inv1  gate1871(.a(G329), .O(gate83inter8));
  nand2 gate1872(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1873(.a(s_189), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1874(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1875(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1876(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate939(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate940(.a(gate85inter0), .b(s_56), .O(gate85inter1));
  and2  gate941(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate942(.a(s_56), .O(gate85inter3));
  inv1  gate943(.a(s_57), .O(gate85inter4));
  nand2 gate944(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate945(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate946(.a(G4), .O(gate85inter7));
  inv1  gate947(.a(G332), .O(gate85inter8));
  nand2 gate948(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate949(.a(s_57), .b(gate85inter3), .O(gate85inter10));
  nor2  gate950(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate951(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate952(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate715(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate716(.a(gate87inter0), .b(s_24), .O(gate87inter1));
  and2  gate717(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate718(.a(s_24), .O(gate87inter3));
  inv1  gate719(.a(s_25), .O(gate87inter4));
  nand2 gate720(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate721(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate722(.a(G12), .O(gate87inter7));
  inv1  gate723(.a(G335), .O(gate87inter8));
  nand2 gate724(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate725(.a(s_25), .b(gate87inter3), .O(gate87inter10));
  nor2  gate726(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate727(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate728(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1289(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1290(.a(gate91inter0), .b(s_106), .O(gate91inter1));
  and2  gate1291(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1292(.a(s_106), .O(gate91inter3));
  inv1  gate1293(.a(s_107), .O(gate91inter4));
  nand2 gate1294(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1295(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1296(.a(G25), .O(gate91inter7));
  inv1  gate1297(.a(G341), .O(gate91inter8));
  nand2 gate1298(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1299(.a(s_107), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1300(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1301(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1302(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate855(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate856(.a(gate97inter0), .b(s_44), .O(gate97inter1));
  and2  gate857(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate858(.a(s_44), .O(gate97inter3));
  inv1  gate859(.a(s_45), .O(gate97inter4));
  nand2 gate860(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate861(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate862(.a(G19), .O(gate97inter7));
  inv1  gate863(.a(G350), .O(gate97inter8));
  nand2 gate864(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate865(.a(s_45), .b(gate97inter3), .O(gate97inter10));
  nor2  gate866(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate867(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate868(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate547(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate548(.a(gate101inter0), .b(s_0), .O(gate101inter1));
  and2  gate549(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate550(.a(s_0), .O(gate101inter3));
  inv1  gate551(.a(s_1), .O(gate101inter4));
  nand2 gate552(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate553(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate554(.a(G20), .O(gate101inter7));
  inv1  gate555(.a(G356), .O(gate101inter8));
  nand2 gate556(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate557(.a(s_1), .b(gate101inter3), .O(gate101inter10));
  nor2  gate558(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate559(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate560(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1037(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1038(.a(gate105inter0), .b(s_70), .O(gate105inter1));
  and2  gate1039(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1040(.a(s_70), .O(gate105inter3));
  inv1  gate1041(.a(s_71), .O(gate105inter4));
  nand2 gate1042(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1043(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1044(.a(G362), .O(gate105inter7));
  inv1  gate1045(.a(G363), .O(gate105inter8));
  nand2 gate1046(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1047(.a(s_71), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1048(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1049(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1050(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1373(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1374(.a(gate107inter0), .b(s_118), .O(gate107inter1));
  and2  gate1375(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1376(.a(s_118), .O(gate107inter3));
  inv1  gate1377(.a(s_119), .O(gate107inter4));
  nand2 gate1378(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1379(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1380(.a(G366), .O(gate107inter7));
  inv1  gate1381(.a(G367), .O(gate107inter8));
  nand2 gate1382(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1383(.a(s_119), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1384(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1385(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1386(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1415(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1416(.a(gate110inter0), .b(s_124), .O(gate110inter1));
  and2  gate1417(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1418(.a(s_124), .O(gate110inter3));
  inv1  gate1419(.a(s_125), .O(gate110inter4));
  nand2 gate1420(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1421(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1422(.a(G372), .O(gate110inter7));
  inv1  gate1423(.a(G373), .O(gate110inter8));
  nand2 gate1424(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1425(.a(s_125), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1426(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1427(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1428(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate743(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate744(.a(gate111inter0), .b(s_28), .O(gate111inter1));
  and2  gate745(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate746(.a(s_28), .O(gate111inter3));
  inv1  gate747(.a(s_29), .O(gate111inter4));
  nand2 gate748(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate749(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate750(.a(G374), .O(gate111inter7));
  inv1  gate751(.a(G375), .O(gate111inter8));
  nand2 gate752(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate753(.a(s_29), .b(gate111inter3), .O(gate111inter10));
  nor2  gate754(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate755(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate756(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1009(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1010(.a(gate112inter0), .b(s_66), .O(gate112inter1));
  and2  gate1011(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1012(.a(s_66), .O(gate112inter3));
  inv1  gate1013(.a(s_67), .O(gate112inter4));
  nand2 gate1014(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1015(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1016(.a(G376), .O(gate112inter7));
  inv1  gate1017(.a(G377), .O(gate112inter8));
  nand2 gate1018(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1019(.a(s_67), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1020(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1021(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1022(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1107(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1108(.a(gate118inter0), .b(s_80), .O(gate118inter1));
  and2  gate1109(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1110(.a(s_80), .O(gate118inter3));
  inv1  gate1111(.a(s_81), .O(gate118inter4));
  nand2 gate1112(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1113(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1114(.a(G388), .O(gate118inter7));
  inv1  gate1115(.a(G389), .O(gate118inter8));
  nand2 gate1116(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1117(.a(s_81), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1118(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1119(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1120(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1975(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1976(.a(gate121inter0), .b(s_204), .O(gate121inter1));
  and2  gate1977(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1978(.a(s_204), .O(gate121inter3));
  inv1  gate1979(.a(s_205), .O(gate121inter4));
  nand2 gate1980(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1981(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1982(.a(G394), .O(gate121inter7));
  inv1  gate1983(.a(G395), .O(gate121inter8));
  nand2 gate1984(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1985(.a(s_205), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1986(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1987(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1988(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1835(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1836(.a(gate123inter0), .b(s_184), .O(gate123inter1));
  and2  gate1837(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1838(.a(s_184), .O(gate123inter3));
  inv1  gate1839(.a(s_185), .O(gate123inter4));
  nand2 gate1840(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1841(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1842(.a(G398), .O(gate123inter7));
  inv1  gate1843(.a(G399), .O(gate123inter8));
  nand2 gate1844(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1845(.a(s_185), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1846(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1847(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1848(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate603(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate604(.a(gate131inter0), .b(s_8), .O(gate131inter1));
  and2  gate605(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate606(.a(s_8), .O(gate131inter3));
  inv1  gate607(.a(s_9), .O(gate131inter4));
  nand2 gate608(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate609(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate610(.a(G414), .O(gate131inter7));
  inv1  gate611(.a(G415), .O(gate131inter8));
  nand2 gate612(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate613(.a(s_9), .b(gate131inter3), .O(gate131inter10));
  nor2  gate614(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate615(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate616(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1121(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1122(.a(gate132inter0), .b(s_82), .O(gate132inter1));
  and2  gate1123(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1124(.a(s_82), .O(gate132inter3));
  inv1  gate1125(.a(s_83), .O(gate132inter4));
  nand2 gate1126(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1127(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1128(.a(G416), .O(gate132inter7));
  inv1  gate1129(.a(G417), .O(gate132inter8));
  nand2 gate1130(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1131(.a(s_83), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1132(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1133(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1134(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate911(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate912(.a(gate135inter0), .b(s_52), .O(gate135inter1));
  and2  gate913(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate914(.a(s_52), .O(gate135inter3));
  inv1  gate915(.a(s_53), .O(gate135inter4));
  nand2 gate916(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate917(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate918(.a(G422), .O(gate135inter7));
  inv1  gate919(.a(G423), .O(gate135inter8));
  nand2 gate920(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate921(.a(s_53), .b(gate135inter3), .O(gate135inter10));
  nor2  gate922(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate923(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate924(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate673(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate674(.a(gate138inter0), .b(s_18), .O(gate138inter1));
  and2  gate675(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate676(.a(s_18), .O(gate138inter3));
  inv1  gate677(.a(s_19), .O(gate138inter4));
  nand2 gate678(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate679(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate680(.a(G432), .O(gate138inter7));
  inv1  gate681(.a(G435), .O(gate138inter8));
  nand2 gate682(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate683(.a(s_19), .b(gate138inter3), .O(gate138inter10));
  nor2  gate684(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate685(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate686(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1191(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1192(.a(gate141inter0), .b(s_92), .O(gate141inter1));
  and2  gate1193(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1194(.a(s_92), .O(gate141inter3));
  inv1  gate1195(.a(s_93), .O(gate141inter4));
  nand2 gate1196(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1197(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1198(.a(G450), .O(gate141inter7));
  inv1  gate1199(.a(G453), .O(gate141inter8));
  nand2 gate1200(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1201(.a(s_93), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1202(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1203(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1204(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate897(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate898(.a(gate144inter0), .b(s_50), .O(gate144inter1));
  and2  gate899(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate900(.a(s_50), .O(gate144inter3));
  inv1  gate901(.a(s_51), .O(gate144inter4));
  nand2 gate902(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate903(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate904(.a(G468), .O(gate144inter7));
  inv1  gate905(.a(G471), .O(gate144inter8));
  nand2 gate906(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate907(.a(s_51), .b(gate144inter3), .O(gate144inter10));
  nor2  gate908(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate909(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate910(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate841(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate842(.a(gate153inter0), .b(s_42), .O(gate153inter1));
  and2  gate843(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate844(.a(s_42), .O(gate153inter3));
  inv1  gate845(.a(s_43), .O(gate153inter4));
  nand2 gate846(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate847(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate848(.a(G426), .O(gate153inter7));
  inv1  gate849(.a(G522), .O(gate153inter8));
  nand2 gate850(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate851(.a(s_43), .b(gate153inter3), .O(gate153inter10));
  nor2  gate852(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate853(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate854(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1401(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1402(.a(gate155inter0), .b(s_122), .O(gate155inter1));
  and2  gate1403(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1404(.a(s_122), .O(gate155inter3));
  inv1  gate1405(.a(s_123), .O(gate155inter4));
  nand2 gate1406(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1407(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1408(.a(G432), .O(gate155inter7));
  inv1  gate1409(.a(G525), .O(gate155inter8));
  nand2 gate1410(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1411(.a(s_123), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1412(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1413(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1414(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1639(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1640(.a(gate157inter0), .b(s_156), .O(gate157inter1));
  and2  gate1641(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1642(.a(s_156), .O(gate157inter3));
  inv1  gate1643(.a(s_157), .O(gate157inter4));
  nand2 gate1644(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1645(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1646(.a(G438), .O(gate157inter7));
  inv1  gate1647(.a(G528), .O(gate157inter8));
  nand2 gate1648(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1649(.a(s_157), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1650(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1651(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1652(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1079(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1080(.a(gate165inter0), .b(s_76), .O(gate165inter1));
  and2  gate1081(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1082(.a(s_76), .O(gate165inter3));
  inv1  gate1083(.a(s_77), .O(gate165inter4));
  nand2 gate1084(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1085(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1086(.a(G462), .O(gate165inter7));
  inv1  gate1087(.a(G540), .O(gate165inter8));
  nand2 gate1088(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1089(.a(s_77), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1090(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1091(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1092(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1247(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1248(.a(gate169inter0), .b(s_100), .O(gate169inter1));
  and2  gate1249(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1250(.a(s_100), .O(gate169inter3));
  inv1  gate1251(.a(s_101), .O(gate169inter4));
  nand2 gate1252(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1253(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1254(.a(G474), .O(gate169inter7));
  inv1  gate1255(.a(G546), .O(gate169inter8));
  nand2 gate1256(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1257(.a(s_101), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1258(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1259(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1260(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1065(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1066(.a(gate170inter0), .b(s_74), .O(gate170inter1));
  and2  gate1067(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1068(.a(s_74), .O(gate170inter3));
  inv1  gate1069(.a(s_75), .O(gate170inter4));
  nand2 gate1070(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1071(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1072(.a(G477), .O(gate170inter7));
  inv1  gate1073(.a(G546), .O(gate170inter8));
  nand2 gate1074(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1075(.a(s_75), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1076(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1077(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1078(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1667(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1668(.a(gate171inter0), .b(s_160), .O(gate171inter1));
  and2  gate1669(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1670(.a(s_160), .O(gate171inter3));
  inv1  gate1671(.a(s_161), .O(gate171inter4));
  nand2 gate1672(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1673(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1674(.a(G480), .O(gate171inter7));
  inv1  gate1675(.a(G549), .O(gate171inter8));
  nand2 gate1676(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1677(.a(s_161), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1678(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1679(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1680(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1765(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1766(.a(gate172inter0), .b(s_174), .O(gate172inter1));
  and2  gate1767(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1768(.a(s_174), .O(gate172inter3));
  inv1  gate1769(.a(s_175), .O(gate172inter4));
  nand2 gate1770(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1771(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1772(.a(G483), .O(gate172inter7));
  inv1  gate1773(.a(G549), .O(gate172inter8));
  nand2 gate1774(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1775(.a(s_175), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1776(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1777(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1778(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1149(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1150(.a(gate174inter0), .b(s_86), .O(gate174inter1));
  and2  gate1151(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1152(.a(s_86), .O(gate174inter3));
  inv1  gate1153(.a(s_87), .O(gate174inter4));
  nand2 gate1154(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1155(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1156(.a(G489), .O(gate174inter7));
  inv1  gate1157(.a(G552), .O(gate174inter8));
  nand2 gate1158(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1159(.a(s_87), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1160(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1161(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1162(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate981(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate982(.a(gate175inter0), .b(s_62), .O(gate175inter1));
  and2  gate983(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate984(.a(s_62), .O(gate175inter3));
  inv1  gate985(.a(s_63), .O(gate175inter4));
  nand2 gate986(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate987(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate988(.a(G492), .O(gate175inter7));
  inv1  gate989(.a(G555), .O(gate175inter8));
  nand2 gate990(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate991(.a(s_63), .b(gate175inter3), .O(gate175inter10));
  nor2  gate992(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate993(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate994(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate729(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate730(.a(gate177inter0), .b(s_26), .O(gate177inter1));
  and2  gate731(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate732(.a(s_26), .O(gate177inter3));
  inv1  gate733(.a(s_27), .O(gate177inter4));
  nand2 gate734(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate735(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate736(.a(G498), .O(gate177inter7));
  inv1  gate737(.a(G558), .O(gate177inter8));
  nand2 gate738(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate739(.a(s_27), .b(gate177inter3), .O(gate177inter10));
  nor2  gate740(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate741(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate742(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1345(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1346(.a(gate182inter0), .b(s_114), .O(gate182inter1));
  and2  gate1347(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1348(.a(s_114), .O(gate182inter3));
  inv1  gate1349(.a(s_115), .O(gate182inter4));
  nand2 gate1350(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1351(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1352(.a(G513), .O(gate182inter7));
  inv1  gate1353(.a(G564), .O(gate182inter8));
  nand2 gate1354(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1355(.a(s_115), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1356(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1357(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1358(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1625(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1626(.a(gate184inter0), .b(s_154), .O(gate184inter1));
  and2  gate1627(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1628(.a(s_154), .O(gate184inter3));
  inv1  gate1629(.a(s_155), .O(gate184inter4));
  nand2 gate1630(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1631(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1632(.a(G519), .O(gate184inter7));
  inv1  gate1633(.a(G567), .O(gate184inter8));
  nand2 gate1634(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1635(.a(s_155), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1636(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1637(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1638(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1471(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1472(.a(gate187inter0), .b(s_132), .O(gate187inter1));
  and2  gate1473(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1474(.a(s_132), .O(gate187inter3));
  inv1  gate1475(.a(s_133), .O(gate187inter4));
  nand2 gate1476(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1477(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1478(.a(G574), .O(gate187inter7));
  inv1  gate1479(.a(G575), .O(gate187inter8));
  nand2 gate1480(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1481(.a(s_133), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1482(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1483(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1484(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate617(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate618(.a(gate195inter0), .b(s_10), .O(gate195inter1));
  and2  gate619(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate620(.a(s_10), .O(gate195inter3));
  inv1  gate621(.a(s_11), .O(gate195inter4));
  nand2 gate622(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate623(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate624(.a(G590), .O(gate195inter7));
  inv1  gate625(.a(G591), .O(gate195inter8));
  nand2 gate626(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate627(.a(s_11), .b(gate195inter3), .O(gate195inter10));
  nor2  gate628(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate629(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate630(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1443(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1444(.a(gate202inter0), .b(s_128), .O(gate202inter1));
  and2  gate1445(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1446(.a(s_128), .O(gate202inter3));
  inv1  gate1447(.a(s_129), .O(gate202inter4));
  nand2 gate1448(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1449(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1450(.a(G612), .O(gate202inter7));
  inv1  gate1451(.a(G617), .O(gate202inter8));
  nand2 gate1452(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1453(.a(s_129), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1454(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1455(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1456(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate883(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate884(.a(gate203inter0), .b(s_48), .O(gate203inter1));
  and2  gate885(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate886(.a(s_48), .O(gate203inter3));
  inv1  gate887(.a(s_49), .O(gate203inter4));
  nand2 gate888(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate889(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate890(.a(G602), .O(gate203inter7));
  inv1  gate891(.a(G612), .O(gate203inter8));
  nand2 gate892(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate893(.a(s_49), .b(gate203inter3), .O(gate203inter10));
  nor2  gate894(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate895(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate896(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1961(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1962(.a(gate204inter0), .b(s_202), .O(gate204inter1));
  and2  gate1963(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1964(.a(s_202), .O(gate204inter3));
  inv1  gate1965(.a(s_203), .O(gate204inter4));
  nand2 gate1966(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1967(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1968(.a(G607), .O(gate204inter7));
  inv1  gate1969(.a(G617), .O(gate204inter8));
  nand2 gate1970(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1971(.a(s_203), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1972(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1973(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1974(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2073(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2074(.a(gate208inter0), .b(s_218), .O(gate208inter1));
  and2  gate2075(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2076(.a(s_218), .O(gate208inter3));
  inv1  gate2077(.a(s_219), .O(gate208inter4));
  nand2 gate2078(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2079(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2080(.a(G627), .O(gate208inter7));
  inv1  gate2081(.a(G637), .O(gate208inter8));
  nand2 gate2082(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2083(.a(s_219), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2084(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2085(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2086(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate631(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate632(.a(gate212inter0), .b(s_12), .O(gate212inter1));
  and2  gate633(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate634(.a(s_12), .O(gate212inter3));
  inv1  gate635(.a(s_13), .O(gate212inter4));
  nand2 gate636(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate637(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate638(.a(G617), .O(gate212inter7));
  inv1  gate639(.a(G669), .O(gate212inter8));
  nand2 gate640(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate641(.a(s_13), .b(gate212inter3), .O(gate212inter10));
  nor2  gate642(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate643(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate644(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate645(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate646(.a(gate213inter0), .b(s_14), .O(gate213inter1));
  and2  gate647(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate648(.a(s_14), .O(gate213inter3));
  inv1  gate649(.a(s_15), .O(gate213inter4));
  nand2 gate650(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate651(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate652(.a(G602), .O(gate213inter7));
  inv1  gate653(.a(G672), .O(gate213inter8));
  nand2 gate654(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate655(.a(s_15), .b(gate213inter3), .O(gate213inter10));
  nor2  gate656(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate657(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate658(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate799(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate800(.a(gate228inter0), .b(s_36), .O(gate228inter1));
  and2  gate801(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate802(.a(s_36), .O(gate228inter3));
  inv1  gate803(.a(s_37), .O(gate228inter4));
  nand2 gate804(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate805(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate806(.a(G696), .O(gate228inter7));
  inv1  gate807(.a(G697), .O(gate228inter8));
  nand2 gate808(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate809(.a(s_37), .b(gate228inter3), .O(gate228inter10));
  nor2  gate810(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate811(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate812(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1989(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1990(.a(gate229inter0), .b(s_206), .O(gate229inter1));
  and2  gate1991(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1992(.a(s_206), .O(gate229inter3));
  inv1  gate1993(.a(s_207), .O(gate229inter4));
  nand2 gate1994(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1995(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1996(.a(G698), .O(gate229inter7));
  inv1  gate1997(.a(G699), .O(gate229inter8));
  nand2 gate1998(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1999(.a(s_207), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2000(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2001(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2002(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate687(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate688(.a(gate233inter0), .b(s_20), .O(gate233inter1));
  and2  gate689(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate690(.a(s_20), .O(gate233inter3));
  inv1  gate691(.a(s_21), .O(gate233inter4));
  nand2 gate692(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate693(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate694(.a(G242), .O(gate233inter7));
  inv1  gate695(.a(G718), .O(gate233inter8));
  nand2 gate696(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate697(.a(s_21), .b(gate233inter3), .O(gate233inter10));
  nor2  gate698(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate699(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate700(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2017(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2018(.a(gate238inter0), .b(s_210), .O(gate238inter1));
  and2  gate2019(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2020(.a(s_210), .O(gate238inter3));
  inv1  gate2021(.a(s_211), .O(gate238inter4));
  nand2 gate2022(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2023(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2024(.a(G257), .O(gate238inter7));
  inv1  gate2025(.a(G709), .O(gate238inter8));
  nand2 gate2026(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2027(.a(s_211), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2028(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2029(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2030(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1317(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1318(.a(gate240inter0), .b(s_110), .O(gate240inter1));
  and2  gate1319(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1320(.a(s_110), .O(gate240inter3));
  inv1  gate1321(.a(s_111), .O(gate240inter4));
  nand2 gate1322(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1323(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1324(.a(G263), .O(gate240inter7));
  inv1  gate1325(.a(G715), .O(gate240inter8));
  nand2 gate1326(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1327(.a(s_111), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1328(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1329(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1330(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate869(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate870(.a(gate245inter0), .b(s_46), .O(gate245inter1));
  and2  gate871(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate872(.a(s_46), .O(gate245inter3));
  inv1  gate873(.a(s_47), .O(gate245inter4));
  nand2 gate874(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate875(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate876(.a(G248), .O(gate245inter7));
  inv1  gate877(.a(G736), .O(gate245inter8));
  nand2 gate878(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate879(.a(s_47), .b(gate245inter3), .O(gate245inter10));
  nor2  gate880(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate881(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate882(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1779(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1780(.a(gate253inter0), .b(s_176), .O(gate253inter1));
  and2  gate1781(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1782(.a(s_176), .O(gate253inter3));
  inv1  gate1783(.a(s_177), .O(gate253inter4));
  nand2 gate1784(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1785(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1786(.a(G260), .O(gate253inter7));
  inv1  gate1787(.a(G748), .O(gate253inter8));
  nand2 gate1788(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1789(.a(s_177), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1790(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1791(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1792(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1597(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1598(.a(gate254inter0), .b(s_150), .O(gate254inter1));
  and2  gate1599(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1600(.a(s_150), .O(gate254inter3));
  inv1  gate1601(.a(s_151), .O(gate254inter4));
  nand2 gate1602(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1603(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1604(.a(G712), .O(gate254inter7));
  inv1  gate1605(.a(G748), .O(gate254inter8));
  nand2 gate1606(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1607(.a(s_151), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1608(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1609(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1610(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1485(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1486(.a(gate257inter0), .b(s_134), .O(gate257inter1));
  and2  gate1487(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1488(.a(s_134), .O(gate257inter3));
  inv1  gate1489(.a(s_135), .O(gate257inter4));
  nand2 gate1490(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1491(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1492(.a(G754), .O(gate257inter7));
  inv1  gate1493(.a(G755), .O(gate257inter8));
  nand2 gate1494(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1495(.a(s_135), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1496(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1497(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1498(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate953(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate954(.a(gate258inter0), .b(s_58), .O(gate258inter1));
  and2  gate955(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate956(.a(s_58), .O(gate258inter3));
  inv1  gate957(.a(s_59), .O(gate258inter4));
  nand2 gate958(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate959(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate960(.a(G756), .O(gate258inter7));
  inv1  gate961(.a(G757), .O(gate258inter8));
  nand2 gate962(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate963(.a(s_59), .b(gate258inter3), .O(gate258inter10));
  nor2  gate964(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate965(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate966(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2129(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2130(.a(gate263inter0), .b(s_226), .O(gate263inter1));
  and2  gate2131(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2132(.a(s_226), .O(gate263inter3));
  inv1  gate2133(.a(s_227), .O(gate263inter4));
  nand2 gate2134(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2135(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2136(.a(G766), .O(gate263inter7));
  inv1  gate2137(.a(G767), .O(gate263inter8));
  nand2 gate2138(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2139(.a(s_227), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2140(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2141(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2142(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1331(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1332(.a(gate266inter0), .b(s_112), .O(gate266inter1));
  and2  gate1333(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1334(.a(s_112), .O(gate266inter3));
  inv1  gate1335(.a(s_113), .O(gate266inter4));
  nand2 gate1336(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1337(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1338(.a(G645), .O(gate266inter7));
  inv1  gate1339(.a(G773), .O(gate266inter8));
  nand2 gate1340(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1341(.a(s_113), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1342(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1343(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1344(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1205(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1206(.a(gate268inter0), .b(s_94), .O(gate268inter1));
  and2  gate1207(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1208(.a(s_94), .O(gate268inter3));
  inv1  gate1209(.a(s_95), .O(gate268inter4));
  nand2 gate1210(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1211(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1212(.a(G651), .O(gate268inter7));
  inv1  gate1213(.a(G779), .O(gate268inter8));
  nand2 gate1214(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1215(.a(s_95), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1216(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1217(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1218(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1555(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1556(.a(gate272inter0), .b(s_144), .O(gate272inter1));
  and2  gate1557(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1558(.a(s_144), .O(gate272inter3));
  inv1  gate1559(.a(s_145), .O(gate272inter4));
  nand2 gate1560(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1561(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1562(.a(G663), .O(gate272inter7));
  inv1  gate1563(.a(G791), .O(gate272inter8));
  nand2 gate1564(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1565(.a(s_145), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1566(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1567(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1568(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2101(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2102(.a(gate281inter0), .b(s_222), .O(gate281inter1));
  and2  gate2103(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2104(.a(s_222), .O(gate281inter3));
  inv1  gate2105(.a(s_223), .O(gate281inter4));
  nand2 gate2106(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2107(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2108(.a(G654), .O(gate281inter7));
  inv1  gate2109(.a(G806), .O(gate281inter8));
  nand2 gate2110(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2111(.a(s_223), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2112(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2113(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2114(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate561(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate562(.a(gate289inter0), .b(s_2), .O(gate289inter1));
  and2  gate563(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate564(.a(s_2), .O(gate289inter3));
  inv1  gate565(.a(s_3), .O(gate289inter4));
  nand2 gate566(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate567(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate568(.a(G818), .O(gate289inter7));
  inv1  gate569(.a(G819), .O(gate289inter8));
  nand2 gate570(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate571(.a(s_3), .b(gate289inter3), .O(gate289inter10));
  nor2  gate572(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate573(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate574(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate925(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate926(.a(gate295inter0), .b(s_54), .O(gate295inter1));
  and2  gate927(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate928(.a(s_54), .O(gate295inter3));
  inv1  gate929(.a(s_55), .O(gate295inter4));
  nand2 gate930(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate931(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate932(.a(G830), .O(gate295inter7));
  inv1  gate933(.a(G831), .O(gate295inter8));
  nand2 gate934(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate935(.a(s_55), .b(gate295inter3), .O(gate295inter10));
  nor2  gate936(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate937(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate938(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1177(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1178(.a(gate396inter0), .b(s_90), .O(gate396inter1));
  and2  gate1179(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1180(.a(s_90), .O(gate396inter3));
  inv1  gate1181(.a(s_91), .O(gate396inter4));
  nand2 gate1182(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1183(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1184(.a(G10), .O(gate396inter7));
  inv1  gate1185(.a(G1063), .O(gate396inter8));
  nand2 gate1186(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1187(.a(s_91), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1188(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1189(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1190(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1569(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1570(.a(gate402inter0), .b(s_146), .O(gate402inter1));
  and2  gate1571(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1572(.a(s_146), .O(gate402inter3));
  inv1  gate1573(.a(s_147), .O(gate402inter4));
  nand2 gate1574(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1575(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1576(.a(G16), .O(gate402inter7));
  inv1  gate1577(.a(G1081), .O(gate402inter8));
  nand2 gate1578(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1579(.a(s_147), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1580(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1581(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1582(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate995(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate996(.a(gate403inter0), .b(s_64), .O(gate403inter1));
  and2  gate997(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate998(.a(s_64), .O(gate403inter3));
  inv1  gate999(.a(s_65), .O(gate403inter4));
  nand2 gate1000(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1001(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1002(.a(G17), .O(gate403inter7));
  inv1  gate1003(.a(G1084), .O(gate403inter8));
  nand2 gate1004(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1005(.a(s_65), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1006(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1007(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1008(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2003(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2004(.a(gate407inter0), .b(s_208), .O(gate407inter1));
  and2  gate2005(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2006(.a(s_208), .O(gate407inter3));
  inv1  gate2007(.a(s_209), .O(gate407inter4));
  nand2 gate2008(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2009(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2010(.a(G21), .O(gate407inter7));
  inv1  gate2011(.a(G1096), .O(gate407inter8));
  nand2 gate2012(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2013(.a(s_209), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2014(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2015(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2016(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1821(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1822(.a(gate409inter0), .b(s_182), .O(gate409inter1));
  and2  gate1823(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1824(.a(s_182), .O(gate409inter3));
  inv1  gate1825(.a(s_183), .O(gate409inter4));
  nand2 gate1826(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1827(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1828(.a(G23), .O(gate409inter7));
  inv1  gate1829(.a(G1102), .O(gate409inter8));
  nand2 gate1830(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1831(.a(s_183), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1832(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1833(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1834(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1219(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1220(.a(gate413inter0), .b(s_96), .O(gate413inter1));
  and2  gate1221(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1222(.a(s_96), .O(gate413inter3));
  inv1  gate1223(.a(s_97), .O(gate413inter4));
  nand2 gate1224(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1225(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1226(.a(G27), .O(gate413inter7));
  inv1  gate1227(.a(G1114), .O(gate413inter8));
  nand2 gate1228(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1229(.a(s_97), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1230(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1231(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1232(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate785(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate786(.a(gate417inter0), .b(s_34), .O(gate417inter1));
  and2  gate787(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate788(.a(s_34), .O(gate417inter3));
  inv1  gate789(.a(s_35), .O(gate417inter4));
  nand2 gate790(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate791(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate792(.a(G31), .O(gate417inter7));
  inv1  gate793(.a(G1126), .O(gate417inter8));
  nand2 gate794(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate795(.a(s_35), .b(gate417inter3), .O(gate417inter10));
  nor2  gate796(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate797(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate798(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1807(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1808(.a(gate420inter0), .b(s_180), .O(gate420inter1));
  and2  gate1809(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1810(.a(s_180), .O(gate420inter3));
  inv1  gate1811(.a(s_181), .O(gate420inter4));
  nand2 gate1812(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1813(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1814(.a(G1036), .O(gate420inter7));
  inv1  gate1815(.a(G1132), .O(gate420inter8));
  nand2 gate1816(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1817(.a(s_181), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1818(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1819(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1820(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1653(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1654(.a(gate421inter0), .b(s_158), .O(gate421inter1));
  and2  gate1655(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1656(.a(s_158), .O(gate421inter3));
  inv1  gate1657(.a(s_159), .O(gate421inter4));
  nand2 gate1658(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1659(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1660(.a(G2), .O(gate421inter7));
  inv1  gate1661(.a(G1135), .O(gate421inter8));
  nand2 gate1662(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1663(.a(s_159), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1664(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1665(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1666(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1709(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1710(.a(gate422inter0), .b(s_166), .O(gate422inter1));
  and2  gate1711(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1712(.a(s_166), .O(gate422inter3));
  inv1  gate1713(.a(s_167), .O(gate422inter4));
  nand2 gate1714(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1715(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1716(.a(G1039), .O(gate422inter7));
  inv1  gate1717(.a(G1135), .O(gate422inter8));
  nand2 gate1718(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1719(.a(s_167), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1720(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1721(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1722(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1751(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1752(.a(gate426inter0), .b(s_172), .O(gate426inter1));
  and2  gate1753(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1754(.a(s_172), .O(gate426inter3));
  inv1  gate1755(.a(s_173), .O(gate426inter4));
  nand2 gate1756(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1757(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1758(.a(G1045), .O(gate426inter7));
  inv1  gate1759(.a(G1141), .O(gate426inter8));
  nand2 gate1760(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1761(.a(s_173), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1762(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1763(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1764(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2087(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2088(.a(gate432inter0), .b(s_220), .O(gate432inter1));
  and2  gate2089(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2090(.a(s_220), .O(gate432inter3));
  inv1  gate2091(.a(s_221), .O(gate432inter4));
  nand2 gate2092(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2093(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2094(.a(G1054), .O(gate432inter7));
  inv1  gate2095(.a(G1150), .O(gate432inter8));
  nand2 gate2096(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2097(.a(s_221), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2098(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2099(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2100(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1737(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1738(.a(gate435inter0), .b(s_170), .O(gate435inter1));
  and2  gate1739(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1740(.a(s_170), .O(gate435inter3));
  inv1  gate1741(.a(s_171), .O(gate435inter4));
  nand2 gate1742(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1743(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1744(.a(G9), .O(gate435inter7));
  inv1  gate1745(.a(G1156), .O(gate435inter8));
  nand2 gate1746(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1747(.a(s_171), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1748(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1749(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1750(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1919(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1920(.a(gate442inter0), .b(s_196), .O(gate442inter1));
  and2  gate1921(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1922(.a(s_196), .O(gate442inter3));
  inv1  gate1923(.a(s_197), .O(gate442inter4));
  nand2 gate1924(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1925(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1926(.a(G1069), .O(gate442inter7));
  inv1  gate1927(.a(G1165), .O(gate442inter8));
  nand2 gate1928(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1929(.a(s_197), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1930(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1931(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1932(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2143(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2144(.a(gate444inter0), .b(s_228), .O(gate444inter1));
  and2  gate2145(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2146(.a(s_228), .O(gate444inter3));
  inv1  gate2147(.a(s_229), .O(gate444inter4));
  nand2 gate2148(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2149(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2150(.a(G1072), .O(gate444inter7));
  inv1  gate2151(.a(G1168), .O(gate444inter8));
  nand2 gate2152(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2153(.a(s_229), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2154(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2155(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2156(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1583(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1584(.a(gate446inter0), .b(s_148), .O(gate446inter1));
  and2  gate1585(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1586(.a(s_148), .O(gate446inter3));
  inv1  gate1587(.a(s_149), .O(gate446inter4));
  nand2 gate1588(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1589(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1590(.a(G1075), .O(gate446inter7));
  inv1  gate1591(.a(G1171), .O(gate446inter8));
  nand2 gate1592(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1593(.a(s_149), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1594(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1595(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1596(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1023(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1024(.a(gate447inter0), .b(s_68), .O(gate447inter1));
  and2  gate1025(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1026(.a(s_68), .O(gate447inter3));
  inv1  gate1027(.a(s_69), .O(gate447inter4));
  nand2 gate1028(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1029(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1030(.a(G15), .O(gate447inter7));
  inv1  gate1031(.a(G1174), .O(gate447inter8));
  nand2 gate1032(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1033(.a(s_69), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1034(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1035(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1036(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1527(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1528(.a(gate448inter0), .b(s_140), .O(gate448inter1));
  and2  gate1529(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1530(.a(s_140), .O(gate448inter3));
  inv1  gate1531(.a(s_141), .O(gate448inter4));
  nand2 gate1532(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1533(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1534(.a(G1078), .O(gate448inter7));
  inv1  gate1535(.a(G1174), .O(gate448inter8));
  nand2 gate1536(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1537(.a(s_141), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1538(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1539(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1540(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1457(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1458(.a(gate454inter0), .b(s_130), .O(gate454inter1));
  and2  gate1459(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1460(.a(s_130), .O(gate454inter3));
  inv1  gate1461(.a(s_131), .O(gate454inter4));
  nand2 gate1462(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1463(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1464(.a(G1087), .O(gate454inter7));
  inv1  gate1465(.a(G1183), .O(gate454inter8));
  nand2 gate1466(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1467(.a(s_131), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1468(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1469(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1470(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1359(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1360(.a(gate456inter0), .b(s_116), .O(gate456inter1));
  and2  gate1361(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1362(.a(s_116), .O(gate456inter3));
  inv1  gate1363(.a(s_117), .O(gate456inter4));
  nand2 gate1364(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1365(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1366(.a(G1090), .O(gate456inter7));
  inv1  gate1367(.a(G1186), .O(gate456inter8));
  nand2 gate1368(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1369(.a(s_117), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1370(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1371(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1372(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1051(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1052(.a(gate462inter0), .b(s_72), .O(gate462inter1));
  and2  gate1053(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1054(.a(s_72), .O(gate462inter3));
  inv1  gate1055(.a(s_73), .O(gate462inter4));
  nand2 gate1056(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1057(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1058(.a(G1099), .O(gate462inter7));
  inv1  gate1059(.a(G1195), .O(gate462inter8));
  nand2 gate1060(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1061(.a(s_73), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1062(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1063(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1064(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1513(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1514(.a(gate469inter0), .b(s_138), .O(gate469inter1));
  and2  gate1515(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1516(.a(s_138), .O(gate469inter3));
  inv1  gate1517(.a(s_139), .O(gate469inter4));
  nand2 gate1518(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1519(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1520(.a(G26), .O(gate469inter7));
  inv1  gate1521(.a(G1207), .O(gate469inter8));
  nand2 gate1522(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1523(.a(s_139), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1524(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1525(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1526(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1499(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1500(.a(gate477inter0), .b(s_136), .O(gate477inter1));
  and2  gate1501(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1502(.a(s_136), .O(gate477inter3));
  inv1  gate1503(.a(s_137), .O(gate477inter4));
  nand2 gate1504(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1505(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1506(.a(G30), .O(gate477inter7));
  inv1  gate1507(.a(G1219), .O(gate477inter8));
  nand2 gate1508(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1509(.a(s_137), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1510(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1511(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1512(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate701(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate702(.a(gate479inter0), .b(s_22), .O(gate479inter1));
  and2  gate703(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate704(.a(s_22), .O(gate479inter3));
  inv1  gate705(.a(s_23), .O(gate479inter4));
  nand2 gate706(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate707(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate708(.a(G31), .O(gate479inter7));
  inv1  gate709(.a(G1222), .O(gate479inter8));
  nand2 gate710(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate711(.a(s_23), .b(gate479inter3), .O(gate479inter10));
  nor2  gate712(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate713(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate714(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1933(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1934(.a(gate480inter0), .b(s_198), .O(gate480inter1));
  and2  gate1935(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1936(.a(s_198), .O(gate480inter3));
  inv1  gate1937(.a(s_199), .O(gate480inter4));
  nand2 gate1938(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1939(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1940(.a(G1126), .O(gate480inter7));
  inv1  gate1941(.a(G1222), .O(gate480inter8));
  nand2 gate1942(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1943(.a(s_199), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1944(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1945(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1946(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate771(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate772(.a(gate481inter0), .b(s_32), .O(gate481inter1));
  and2  gate773(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate774(.a(s_32), .O(gate481inter3));
  inv1  gate775(.a(s_33), .O(gate481inter4));
  nand2 gate776(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate777(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate778(.a(G32), .O(gate481inter7));
  inv1  gate779(.a(G1225), .O(gate481inter8));
  nand2 gate780(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate781(.a(s_33), .b(gate481inter3), .O(gate481inter10));
  nor2  gate782(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate783(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate784(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1093(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1094(.a(gate482inter0), .b(s_78), .O(gate482inter1));
  and2  gate1095(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1096(.a(s_78), .O(gate482inter3));
  inv1  gate1097(.a(s_79), .O(gate482inter4));
  nand2 gate1098(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1099(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1100(.a(G1129), .O(gate482inter7));
  inv1  gate1101(.a(G1225), .O(gate482inter8));
  nand2 gate1102(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1103(.a(s_79), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1104(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1105(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1106(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1681(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1682(.a(gate484inter0), .b(s_162), .O(gate484inter1));
  and2  gate1683(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1684(.a(s_162), .O(gate484inter3));
  inv1  gate1685(.a(s_163), .O(gate484inter4));
  nand2 gate1686(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1687(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1688(.a(G1230), .O(gate484inter7));
  inv1  gate1689(.a(G1231), .O(gate484inter8));
  nand2 gate1690(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1691(.a(s_163), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1692(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1693(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1694(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate2059(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2060(.a(gate487inter0), .b(s_216), .O(gate487inter1));
  and2  gate2061(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2062(.a(s_216), .O(gate487inter3));
  inv1  gate2063(.a(s_217), .O(gate487inter4));
  nand2 gate2064(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2065(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2066(.a(G1236), .O(gate487inter7));
  inv1  gate2067(.a(G1237), .O(gate487inter8));
  nand2 gate2068(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2069(.a(s_217), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2070(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2071(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2072(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2045(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2046(.a(gate493inter0), .b(s_214), .O(gate493inter1));
  and2  gate2047(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2048(.a(s_214), .O(gate493inter3));
  inv1  gate2049(.a(s_215), .O(gate493inter4));
  nand2 gate2050(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2051(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2052(.a(G1248), .O(gate493inter7));
  inv1  gate2053(.a(G1249), .O(gate493inter8));
  nand2 gate2054(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2055(.a(s_215), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2056(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2057(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2058(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate575(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate576(.a(gate494inter0), .b(s_4), .O(gate494inter1));
  and2  gate577(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate578(.a(s_4), .O(gate494inter3));
  inv1  gate579(.a(s_5), .O(gate494inter4));
  nand2 gate580(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate581(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate582(.a(G1250), .O(gate494inter7));
  inv1  gate583(.a(G1251), .O(gate494inter8));
  nand2 gate584(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate585(.a(s_5), .b(gate494inter3), .O(gate494inter10));
  nor2  gate586(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate587(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate588(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1135(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1136(.a(gate496inter0), .b(s_84), .O(gate496inter1));
  and2  gate1137(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1138(.a(s_84), .O(gate496inter3));
  inv1  gate1139(.a(s_85), .O(gate496inter4));
  nand2 gate1140(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1141(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1142(.a(G1254), .O(gate496inter7));
  inv1  gate1143(.a(G1255), .O(gate496inter8));
  nand2 gate1144(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1145(.a(s_85), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1146(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1147(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1148(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate2031(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2032(.a(gate497inter0), .b(s_212), .O(gate497inter1));
  and2  gate2033(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2034(.a(s_212), .O(gate497inter3));
  inv1  gate2035(.a(s_213), .O(gate497inter4));
  nand2 gate2036(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2037(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2038(.a(G1256), .O(gate497inter7));
  inv1  gate2039(.a(G1257), .O(gate497inter8));
  nand2 gate2040(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2041(.a(s_213), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2042(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2043(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2044(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1429(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1430(.a(gate499inter0), .b(s_126), .O(gate499inter1));
  and2  gate1431(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1432(.a(s_126), .O(gate499inter3));
  inv1  gate1433(.a(s_127), .O(gate499inter4));
  nand2 gate1434(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1435(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1436(.a(G1260), .O(gate499inter7));
  inv1  gate1437(.a(G1261), .O(gate499inter8));
  nand2 gate1438(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1439(.a(s_127), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1440(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1441(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1442(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1905(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1906(.a(gate501inter0), .b(s_194), .O(gate501inter1));
  and2  gate1907(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1908(.a(s_194), .O(gate501inter3));
  inv1  gate1909(.a(s_195), .O(gate501inter4));
  nand2 gate1910(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1911(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1912(.a(G1264), .O(gate501inter7));
  inv1  gate1913(.a(G1265), .O(gate501inter8));
  nand2 gate1914(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1915(.a(s_195), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1916(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1917(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1918(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1891(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1892(.a(gate502inter0), .b(s_192), .O(gate502inter1));
  and2  gate1893(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1894(.a(s_192), .O(gate502inter3));
  inv1  gate1895(.a(s_193), .O(gate502inter4));
  nand2 gate1896(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1897(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1898(.a(G1266), .O(gate502inter7));
  inv1  gate1899(.a(G1267), .O(gate502inter8));
  nand2 gate1900(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1901(.a(s_193), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1902(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1903(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1904(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1695(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1696(.a(gate509inter0), .b(s_164), .O(gate509inter1));
  and2  gate1697(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1698(.a(s_164), .O(gate509inter3));
  inv1  gate1699(.a(s_165), .O(gate509inter4));
  nand2 gate1700(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1701(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1702(.a(G1280), .O(gate509inter7));
  inv1  gate1703(.a(G1281), .O(gate509inter8));
  nand2 gate1704(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1705(.a(s_165), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1706(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1707(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1708(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1261(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1262(.a(gate512inter0), .b(s_102), .O(gate512inter1));
  and2  gate1263(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1264(.a(s_102), .O(gate512inter3));
  inv1  gate1265(.a(s_103), .O(gate512inter4));
  nand2 gate1266(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1267(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1268(.a(G1286), .O(gate512inter7));
  inv1  gate1269(.a(G1287), .O(gate512inter8));
  nand2 gate1270(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1271(.a(s_103), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1272(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1273(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1274(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1723(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1724(.a(gate513inter0), .b(s_168), .O(gate513inter1));
  and2  gate1725(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1726(.a(s_168), .O(gate513inter3));
  inv1  gate1727(.a(s_169), .O(gate513inter4));
  nand2 gate1728(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1729(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1730(.a(G1288), .O(gate513inter7));
  inv1  gate1731(.a(G1289), .O(gate513inter8));
  nand2 gate1732(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1733(.a(s_169), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1734(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1735(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1736(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule