module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2213(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2214(.a(gate14inter0), .b(s_238), .O(gate14inter1));
  and2  gate2215(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2216(.a(s_238), .O(gate14inter3));
  inv1  gate2217(.a(s_239), .O(gate14inter4));
  nand2 gate2218(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2219(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2220(.a(G11), .O(gate14inter7));
  inv1  gate2221(.a(G12), .O(gate14inter8));
  nand2 gate2222(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2223(.a(s_239), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2224(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2225(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2226(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate799(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate800(.a(gate15inter0), .b(s_36), .O(gate15inter1));
  and2  gate801(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate802(.a(s_36), .O(gate15inter3));
  inv1  gate803(.a(s_37), .O(gate15inter4));
  nand2 gate804(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate805(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate806(.a(G13), .O(gate15inter7));
  inv1  gate807(.a(G14), .O(gate15inter8));
  nand2 gate808(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate809(.a(s_37), .b(gate15inter3), .O(gate15inter10));
  nor2  gate810(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate811(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate812(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2073(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2074(.a(gate18inter0), .b(s_218), .O(gate18inter1));
  and2  gate2075(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2076(.a(s_218), .O(gate18inter3));
  inv1  gate2077(.a(s_219), .O(gate18inter4));
  nand2 gate2078(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2079(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2080(.a(G19), .O(gate18inter7));
  inv1  gate2081(.a(G20), .O(gate18inter8));
  nand2 gate2082(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2083(.a(s_219), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2084(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2085(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2086(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate547(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate548(.a(gate19inter0), .b(s_0), .O(gate19inter1));
  and2  gate549(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate550(.a(s_0), .O(gate19inter3));
  inv1  gate551(.a(s_1), .O(gate19inter4));
  nand2 gate552(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate553(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate554(.a(G21), .O(gate19inter7));
  inv1  gate555(.a(G22), .O(gate19inter8));
  nand2 gate556(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate557(.a(s_1), .b(gate19inter3), .O(gate19inter10));
  nor2  gate558(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate559(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate560(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1709(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1710(.a(gate22inter0), .b(s_166), .O(gate22inter1));
  and2  gate1711(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1712(.a(s_166), .O(gate22inter3));
  inv1  gate1713(.a(s_167), .O(gate22inter4));
  nand2 gate1714(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1715(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1716(.a(G27), .O(gate22inter7));
  inv1  gate1717(.a(G28), .O(gate22inter8));
  nand2 gate1718(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1719(.a(s_167), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1720(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1721(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1722(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2143(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2144(.a(gate23inter0), .b(s_228), .O(gate23inter1));
  and2  gate2145(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2146(.a(s_228), .O(gate23inter3));
  inv1  gate2147(.a(s_229), .O(gate23inter4));
  nand2 gate2148(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2149(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2150(.a(G29), .O(gate23inter7));
  inv1  gate2151(.a(G30), .O(gate23inter8));
  nand2 gate2152(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2153(.a(s_229), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2154(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2155(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2156(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1597(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1598(.a(gate29inter0), .b(s_150), .O(gate29inter1));
  and2  gate1599(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1600(.a(s_150), .O(gate29inter3));
  inv1  gate1601(.a(s_151), .O(gate29inter4));
  nand2 gate1602(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1603(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1604(.a(G3), .O(gate29inter7));
  inv1  gate1605(.a(G7), .O(gate29inter8));
  nand2 gate1606(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1607(.a(s_151), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1608(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1609(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1610(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate659(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate660(.a(gate31inter0), .b(s_16), .O(gate31inter1));
  and2  gate661(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate662(.a(s_16), .O(gate31inter3));
  inv1  gate663(.a(s_17), .O(gate31inter4));
  nand2 gate664(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate665(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate666(.a(G4), .O(gate31inter7));
  inv1  gate667(.a(G8), .O(gate31inter8));
  nand2 gate668(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate669(.a(s_17), .b(gate31inter3), .O(gate31inter10));
  nor2  gate670(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate671(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate672(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1975(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1976(.a(gate32inter0), .b(s_204), .O(gate32inter1));
  and2  gate1977(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1978(.a(s_204), .O(gate32inter3));
  inv1  gate1979(.a(s_205), .O(gate32inter4));
  nand2 gate1980(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1981(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1982(.a(G12), .O(gate32inter7));
  inv1  gate1983(.a(G16), .O(gate32inter8));
  nand2 gate1984(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1985(.a(s_205), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1986(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1987(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1988(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1163(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1164(.a(gate36inter0), .b(s_88), .O(gate36inter1));
  and2  gate1165(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1166(.a(s_88), .O(gate36inter3));
  inv1  gate1167(.a(s_89), .O(gate36inter4));
  nand2 gate1168(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1169(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1170(.a(G26), .O(gate36inter7));
  inv1  gate1171(.a(G30), .O(gate36inter8));
  nand2 gate1172(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1173(.a(s_89), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1174(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1175(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1176(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate771(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate772(.a(gate38inter0), .b(s_32), .O(gate38inter1));
  and2  gate773(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate774(.a(s_32), .O(gate38inter3));
  inv1  gate775(.a(s_33), .O(gate38inter4));
  nand2 gate776(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate777(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate778(.a(G27), .O(gate38inter7));
  inv1  gate779(.a(G31), .O(gate38inter8));
  nand2 gate780(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate781(.a(s_33), .b(gate38inter3), .O(gate38inter10));
  nor2  gate782(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate783(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate784(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1079(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1080(.a(gate40inter0), .b(s_76), .O(gate40inter1));
  and2  gate1081(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1082(.a(s_76), .O(gate40inter3));
  inv1  gate1083(.a(s_77), .O(gate40inter4));
  nand2 gate1084(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1085(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1086(.a(G28), .O(gate40inter7));
  inv1  gate1087(.a(G32), .O(gate40inter8));
  nand2 gate1088(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1089(.a(s_77), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1090(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1091(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1092(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1821(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1822(.a(gate41inter0), .b(s_182), .O(gate41inter1));
  and2  gate1823(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1824(.a(s_182), .O(gate41inter3));
  inv1  gate1825(.a(s_183), .O(gate41inter4));
  nand2 gate1826(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1827(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1828(.a(G1), .O(gate41inter7));
  inv1  gate1829(.a(G266), .O(gate41inter8));
  nand2 gate1830(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1831(.a(s_183), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1832(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1833(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1834(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2647(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2648(.a(gate42inter0), .b(s_300), .O(gate42inter1));
  and2  gate2649(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2650(.a(s_300), .O(gate42inter3));
  inv1  gate2651(.a(s_301), .O(gate42inter4));
  nand2 gate2652(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2653(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2654(.a(G2), .O(gate42inter7));
  inv1  gate2655(.a(G266), .O(gate42inter8));
  nand2 gate2656(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2657(.a(s_301), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2658(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2659(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2660(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2115(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2116(.a(gate51inter0), .b(s_224), .O(gate51inter1));
  and2  gate2117(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2118(.a(s_224), .O(gate51inter3));
  inv1  gate2119(.a(s_225), .O(gate51inter4));
  nand2 gate2120(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2121(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2122(.a(G11), .O(gate51inter7));
  inv1  gate2123(.a(G281), .O(gate51inter8));
  nand2 gate2124(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2125(.a(s_225), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2126(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2127(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2128(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1135(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1136(.a(gate55inter0), .b(s_84), .O(gate55inter1));
  and2  gate1137(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1138(.a(s_84), .O(gate55inter3));
  inv1  gate1139(.a(s_85), .O(gate55inter4));
  nand2 gate1140(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1141(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1142(.a(G15), .O(gate55inter7));
  inv1  gate1143(.a(G287), .O(gate55inter8));
  nand2 gate1144(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1145(.a(s_85), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1146(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1147(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1148(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1499(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1500(.a(gate57inter0), .b(s_136), .O(gate57inter1));
  and2  gate1501(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1502(.a(s_136), .O(gate57inter3));
  inv1  gate1503(.a(s_137), .O(gate57inter4));
  nand2 gate1504(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1505(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1506(.a(G17), .O(gate57inter7));
  inv1  gate1507(.a(G290), .O(gate57inter8));
  nand2 gate1508(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1509(.a(s_137), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1510(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1511(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1512(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2269(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2270(.a(gate59inter0), .b(s_246), .O(gate59inter1));
  and2  gate2271(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2272(.a(s_246), .O(gate59inter3));
  inv1  gate2273(.a(s_247), .O(gate59inter4));
  nand2 gate2274(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2275(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2276(.a(G19), .O(gate59inter7));
  inv1  gate2277(.a(G293), .O(gate59inter8));
  nand2 gate2278(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2279(.a(s_247), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2280(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2281(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2282(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1121(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1122(.a(gate65inter0), .b(s_82), .O(gate65inter1));
  and2  gate1123(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1124(.a(s_82), .O(gate65inter3));
  inv1  gate1125(.a(s_83), .O(gate65inter4));
  nand2 gate1126(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1127(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1128(.a(G25), .O(gate65inter7));
  inv1  gate1129(.a(G302), .O(gate65inter8));
  nand2 gate1130(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1131(.a(s_83), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1132(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1133(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1134(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2563(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2564(.a(gate67inter0), .b(s_288), .O(gate67inter1));
  and2  gate2565(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2566(.a(s_288), .O(gate67inter3));
  inv1  gate2567(.a(s_289), .O(gate67inter4));
  nand2 gate2568(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2569(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2570(.a(G27), .O(gate67inter7));
  inv1  gate2571(.a(G305), .O(gate67inter8));
  nand2 gate2572(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2573(.a(s_289), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2574(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2575(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2576(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate897(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate898(.a(gate71inter0), .b(s_50), .O(gate71inter1));
  and2  gate899(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate900(.a(s_50), .O(gate71inter3));
  inv1  gate901(.a(s_51), .O(gate71inter4));
  nand2 gate902(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate903(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate904(.a(G31), .O(gate71inter7));
  inv1  gate905(.a(G311), .O(gate71inter8));
  nand2 gate906(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate907(.a(s_51), .b(gate71inter3), .O(gate71inter10));
  nor2  gate908(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate909(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate910(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1779(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1780(.a(gate73inter0), .b(s_176), .O(gate73inter1));
  and2  gate1781(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1782(.a(s_176), .O(gate73inter3));
  inv1  gate1783(.a(s_177), .O(gate73inter4));
  nand2 gate1784(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1785(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1786(.a(G1), .O(gate73inter7));
  inv1  gate1787(.a(G314), .O(gate73inter8));
  nand2 gate1788(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1789(.a(s_177), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1790(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1791(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1792(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1247(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1248(.a(gate74inter0), .b(s_100), .O(gate74inter1));
  and2  gate1249(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1250(.a(s_100), .O(gate74inter3));
  inv1  gate1251(.a(s_101), .O(gate74inter4));
  nand2 gate1252(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1253(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1254(.a(G5), .O(gate74inter7));
  inv1  gate1255(.a(G314), .O(gate74inter8));
  nand2 gate1256(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1257(.a(s_101), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1258(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1259(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1260(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1751(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1752(.a(gate75inter0), .b(s_172), .O(gate75inter1));
  and2  gate1753(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1754(.a(s_172), .O(gate75inter3));
  inv1  gate1755(.a(s_173), .O(gate75inter4));
  nand2 gate1756(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1757(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1758(.a(G9), .O(gate75inter7));
  inv1  gate1759(.a(G317), .O(gate75inter8));
  nand2 gate1760(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1761(.a(s_173), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1762(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1763(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1764(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1023(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1024(.a(gate84inter0), .b(s_68), .O(gate84inter1));
  and2  gate1025(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1026(.a(s_68), .O(gate84inter3));
  inv1  gate1027(.a(s_69), .O(gate84inter4));
  nand2 gate1028(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1029(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1030(.a(G15), .O(gate84inter7));
  inv1  gate1031(.a(G329), .O(gate84inter8));
  nand2 gate1032(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1033(.a(s_69), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1034(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1035(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1036(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1065(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1066(.a(gate86inter0), .b(s_74), .O(gate86inter1));
  and2  gate1067(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1068(.a(s_74), .O(gate86inter3));
  inv1  gate1069(.a(s_75), .O(gate86inter4));
  nand2 gate1070(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1071(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1072(.a(G8), .O(gate86inter7));
  inv1  gate1073(.a(G332), .O(gate86inter8));
  nand2 gate1074(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1075(.a(s_75), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1076(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1077(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1078(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate575(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate576(.a(gate87inter0), .b(s_4), .O(gate87inter1));
  and2  gate577(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate578(.a(s_4), .O(gate87inter3));
  inv1  gate579(.a(s_5), .O(gate87inter4));
  nand2 gate580(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate581(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate582(.a(G12), .O(gate87inter7));
  inv1  gate583(.a(G335), .O(gate87inter8));
  nand2 gate584(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate585(.a(s_5), .b(gate87inter3), .O(gate87inter10));
  nor2  gate586(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate587(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate588(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1863(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1864(.a(gate88inter0), .b(s_188), .O(gate88inter1));
  and2  gate1865(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1866(.a(s_188), .O(gate88inter3));
  inv1  gate1867(.a(s_189), .O(gate88inter4));
  nand2 gate1868(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1869(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1870(.a(G16), .O(gate88inter7));
  inv1  gate1871(.a(G335), .O(gate88inter8));
  nand2 gate1872(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1873(.a(s_189), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1874(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1875(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1876(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate939(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate940(.a(gate90inter0), .b(s_56), .O(gate90inter1));
  and2  gate941(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate942(.a(s_56), .O(gate90inter3));
  inv1  gate943(.a(s_57), .O(gate90inter4));
  nand2 gate944(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate945(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate946(.a(G21), .O(gate90inter7));
  inv1  gate947(.a(G338), .O(gate90inter8));
  nand2 gate948(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate949(.a(s_57), .b(gate90inter3), .O(gate90inter10));
  nor2  gate950(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate951(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate952(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1289(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1290(.a(gate95inter0), .b(s_106), .O(gate95inter1));
  and2  gate1291(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1292(.a(s_106), .O(gate95inter3));
  inv1  gate1293(.a(s_107), .O(gate95inter4));
  nand2 gate1294(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1295(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1296(.a(G26), .O(gate95inter7));
  inv1  gate1297(.a(G347), .O(gate95inter8));
  nand2 gate1298(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1299(.a(s_107), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1300(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1301(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1302(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate2633(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate2634(.a(gate98inter0), .b(s_298), .O(gate98inter1));
  and2  gate2635(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate2636(.a(s_298), .O(gate98inter3));
  inv1  gate2637(.a(s_299), .O(gate98inter4));
  nand2 gate2638(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2639(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2640(.a(G23), .O(gate98inter7));
  inv1  gate2641(.a(G350), .O(gate98inter8));
  nand2 gate2642(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2643(.a(s_299), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2644(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2645(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2646(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2157(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2158(.a(gate99inter0), .b(s_230), .O(gate99inter1));
  and2  gate2159(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2160(.a(s_230), .O(gate99inter3));
  inv1  gate2161(.a(s_231), .O(gate99inter4));
  nand2 gate2162(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2163(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2164(.a(G27), .O(gate99inter7));
  inv1  gate2165(.a(G353), .O(gate99inter8));
  nand2 gate2166(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2167(.a(s_231), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2168(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2169(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2170(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2437(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2438(.a(gate101inter0), .b(s_270), .O(gate101inter1));
  and2  gate2439(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2440(.a(s_270), .O(gate101inter3));
  inv1  gate2441(.a(s_271), .O(gate101inter4));
  nand2 gate2442(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2443(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2444(.a(G20), .O(gate101inter7));
  inv1  gate2445(.a(G356), .O(gate101inter8));
  nand2 gate2446(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2447(.a(s_271), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2448(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2449(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2450(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1793(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1794(.a(gate102inter0), .b(s_178), .O(gate102inter1));
  and2  gate1795(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1796(.a(s_178), .O(gate102inter3));
  inv1  gate1797(.a(s_179), .O(gate102inter4));
  nand2 gate1798(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1799(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1800(.a(G24), .O(gate102inter7));
  inv1  gate1801(.a(G356), .O(gate102inter8));
  nand2 gate1802(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1803(.a(s_179), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1804(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1805(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1806(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate2451(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2452(.a(gate103inter0), .b(s_272), .O(gate103inter1));
  and2  gate2453(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2454(.a(s_272), .O(gate103inter3));
  inv1  gate2455(.a(s_273), .O(gate103inter4));
  nand2 gate2456(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2457(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2458(.a(G28), .O(gate103inter7));
  inv1  gate2459(.a(G359), .O(gate103inter8));
  nand2 gate2460(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2461(.a(s_273), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2462(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2463(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2464(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1919(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1920(.a(gate106inter0), .b(s_196), .O(gate106inter1));
  and2  gate1921(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1922(.a(s_196), .O(gate106inter3));
  inv1  gate1923(.a(s_197), .O(gate106inter4));
  nand2 gate1924(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1925(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1926(.a(G364), .O(gate106inter7));
  inv1  gate1927(.a(G365), .O(gate106inter8));
  nand2 gate1928(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1929(.a(s_197), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1930(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1931(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1932(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1653(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1654(.a(gate109inter0), .b(s_158), .O(gate109inter1));
  and2  gate1655(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1656(.a(s_158), .O(gate109inter3));
  inv1  gate1657(.a(s_159), .O(gate109inter4));
  nand2 gate1658(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1659(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1660(.a(G370), .O(gate109inter7));
  inv1  gate1661(.a(G371), .O(gate109inter8));
  nand2 gate1662(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1663(.a(s_159), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1664(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1665(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1666(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1625(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1626(.a(gate112inter0), .b(s_154), .O(gate112inter1));
  and2  gate1627(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1628(.a(s_154), .O(gate112inter3));
  inv1  gate1629(.a(s_155), .O(gate112inter4));
  nand2 gate1630(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1631(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1632(.a(G376), .O(gate112inter7));
  inv1  gate1633(.a(G377), .O(gate112inter8));
  nand2 gate1634(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1635(.a(s_155), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1636(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1637(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1638(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate813(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate814(.a(gate115inter0), .b(s_38), .O(gate115inter1));
  and2  gate815(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate816(.a(s_38), .O(gate115inter3));
  inv1  gate817(.a(s_39), .O(gate115inter4));
  nand2 gate818(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate819(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate820(.a(G382), .O(gate115inter7));
  inv1  gate821(.a(G383), .O(gate115inter8));
  nand2 gate822(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate823(.a(s_39), .b(gate115inter3), .O(gate115inter10));
  nor2  gate824(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate825(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate826(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1933(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1934(.a(gate117inter0), .b(s_198), .O(gate117inter1));
  and2  gate1935(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1936(.a(s_198), .O(gate117inter3));
  inv1  gate1937(.a(s_199), .O(gate117inter4));
  nand2 gate1938(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1939(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1940(.a(G386), .O(gate117inter7));
  inv1  gate1941(.a(G387), .O(gate117inter8));
  nand2 gate1942(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1943(.a(s_199), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1944(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1945(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1946(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1373(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1374(.a(gate119inter0), .b(s_118), .O(gate119inter1));
  and2  gate1375(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1376(.a(s_118), .O(gate119inter3));
  inv1  gate1377(.a(s_119), .O(gate119inter4));
  nand2 gate1378(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1379(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1380(.a(G390), .O(gate119inter7));
  inv1  gate1381(.a(G391), .O(gate119inter8));
  nand2 gate1382(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1383(.a(s_119), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1384(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1385(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1386(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1051(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1052(.a(gate120inter0), .b(s_72), .O(gate120inter1));
  and2  gate1053(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1054(.a(s_72), .O(gate120inter3));
  inv1  gate1055(.a(s_73), .O(gate120inter4));
  nand2 gate1056(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1057(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1058(.a(G392), .O(gate120inter7));
  inv1  gate1059(.a(G393), .O(gate120inter8));
  nand2 gate1060(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1061(.a(s_73), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1062(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1063(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1064(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate2367(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2368(.a(gate121inter0), .b(s_260), .O(gate121inter1));
  and2  gate2369(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2370(.a(s_260), .O(gate121inter3));
  inv1  gate2371(.a(s_261), .O(gate121inter4));
  nand2 gate2372(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2373(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2374(.a(G394), .O(gate121inter7));
  inv1  gate2375(.a(G395), .O(gate121inter8));
  nand2 gate2376(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2377(.a(s_261), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2378(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2379(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2380(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1849(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1850(.a(gate125inter0), .b(s_186), .O(gate125inter1));
  and2  gate1851(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1852(.a(s_186), .O(gate125inter3));
  inv1  gate1853(.a(s_187), .O(gate125inter4));
  nand2 gate1854(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1855(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1856(.a(G402), .O(gate125inter7));
  inv1  gate1857(.a(G403), .O(gate125inter8));
  nand2 gate1858(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1859(.a(s_187), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1860(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1861(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1862(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2059(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2060(.a(gate127inter0), .b(s_216), .O(gate127inter1));
  and2  gate2061(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2062(.a(s_216), .O(gate127inter3));
  inv1  gate2063(.a(s_217), .O(gate127inter4));
  nand2 gate2064(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2065(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2066(.a(G406), .O(gate127inter7));
  inv1  gate2067(.a(G407), .O(gate127inter8));
  nand2 gate2068(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2069(.a(s_217), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2070(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2071(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2072(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate2591(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2592(.a(gate128inter0), .b(s_292), .O(gate128inter1));
  and2  gate2593(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2594(.a(s_292), .O(gate128inter3));
  inv1  gate2595(.a(s_293), .O(gate128inter4));
  nand2 gate2596(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2597(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2598(.a(G408), .O(gate128inter7));
  inv1  gate2599(.a(G409), .O(gate128inter8));
  nand2 gate2600(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2601(.a(s_293), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2602(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2603(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2604(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate561(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate562(.a(gate130inter0), .b(s_2), .O(gate130inter1));
  and2  gate563(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate564(.a(s_2), .O(gate130inter3));
  inv1  gate565(.a(s_3), .O(gate130inter4));
  nand2 gate566(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate567(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate568(.a(G412), .O(gate130inter7));
  inv1  gate569(.a(G413), .O(gate130inter8));
  nand2 gate570(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate571(.a(s_3), .b(gate130inter3), .O(gate130inter10));
  nor2  gate572(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate573(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate574(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1639(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1640(.a(gate133inter0), .b(s_156), .O(gate133inter1));
  and2  gate1641(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1642(.a(s_156), .O(gate133inter3));
  inv1  gate1643(.a(s_157), .O(gate133inter4));
  nand2 gate1644(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1645(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1646(.a(G418), .O(gate133inter7));
  inv1  gate1647(.a(G419), .O(gate133inter8));
  nand2 gate1648(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1649(.a(s_157), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1650(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1651(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1652(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate2283(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2284(.a(gate134inter0), .b(s_248), .O(gate134inter1));
  and2  gate2285(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2286(.a(s_248), .O(gate134inter3));
  inv1  gate2287(.a(s_249), .O(gate134inter4));
  nand2 gate2288(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2289(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2290(.a(G420), .O(gate134inter7));
  inv1  gate2291(.a(G421), .O(gate134inter8));
  nand2 gate2292(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2293(.a(s_249), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2294(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2295(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2296(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2479(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2480(.a(gate143inter0), .b(s_276), .O(gate143inter1));
  and2  gate2481(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2482(.a(s_276), .O(gate143inter3));
  inv1  gate2483(.a(s_277), .O(gate143inter4));
  nand2 gate2484(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2485(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2486(.a(G462), .O(gate143inter7));
  inv1  gate2487(.a(G465), .O(gate143inter8));
  nand2 gate2488(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2489(.a(s_277), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2490(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2491(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2492(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate995(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate996(.a(gate144inter0), .b(s_64), .O(gate144inter1));
  and2  gate997(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate998(.a(s_64), .O(gate144inter3));
  inv1  gate999(.a(s_65), .O(gate144inter4));
  nand2 gate1000(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1001(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1002(.a(G468), .O(gate144inter7));
  inv1  gate1003(.a(G471), .O(gate144inter8));
  nand2 gate1004(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1005(.a(s_65), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1006(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1007(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1008(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2353(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2354(.a(gate145inter0), .b(s_258), .O(gate145inter1));
  and2  gate2355(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2356(.a(s_258), .O(gate145inter3));
  inv1  gate2357(.a(s_259), .O(gate145inter4));
  nand2 gate2358(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2359(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2360(.a(G474), .O(gate145inter7));
  inv1  gate2361(.a(G477), .O(gate145inter8));
  nand2 gate2362(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2363(.a(s_259), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2364(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2365(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2366(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1303(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1304(.a(gate146inter0), .b(s_108), .O(gate146inter1));
  and2  gate1305(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1306(.a(s_108), .O(gate146inter3));
  inv1  gate1307(.a(s_109), .O(gate146inter4));
  nand2 gate1308(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1309(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1310(.a(G480), .O(gate146inter7));
  inv1  gate1311(.a(G483), .O(gate146inter8));
  nand2 gate1312(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1313(.a(s_109), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1314(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1315(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1316(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2311(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2312(.a(gate149inter0), .b(s_252), .O(gate149inter1));
  and2  gate2313(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2314(.a(s_252), .O(gate149inter3));
  inv1  gate2315(.a(s_253), .O(gate149inter4));
  nand2 gate2316(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2317(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2318(.a(G498), .O(gate149inter7));
  inv1  gate2319(.a(G501), .O(gate149inter8));
  nand2 gate2320(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2321(.a(s_253), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2322(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2323(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2324(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1107(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1108(.a(gate154inter0), .b(s_80), .O(gate154inter1));
  and2  gate1109(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1110(.a(s_80), .O(gate154inter3));
  inv1  gate1111(.a(s_81), .O(gate154inter4));
  nand2 gate1112(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1113(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1114(.a(G429), .O(gate154inter7));
  inv1  gate1115(.a(G522), .O(gate154inter8));
  nand2 gate1116(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1117(.a(s_81), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1118(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1119(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1120(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate883(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate884(.a(gate155inter0), .b(s_48), .O(gate155inter1));
  and2  gate885(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate886(.a(s_48), .O(gate155inter3));
  inv1  gate887(.a(s_49), .O(gate155inter4));
  nand2 gate888(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate889(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate890(.a(G432), .O(gate155inter7));
  inv1  gate891(.a(G525), .O(gate155inter8));
  nand2 gate892(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate893(.a(s_49), .b(gate155inter3), .O(gate155inter10));
  nor2  gate894(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate895(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate896(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate589(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate590(.a(gate157inter0), .b(s_6), .O(gate157inter1));
  and2  gate591(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate592(.a(s_6), .O(gate157inter3));
  inv1  gate593(.a(s_7), .O(gate157inter4));
  nand2 gate594(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate595(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate596(.a(G438), .O(gate157inter7));
  inv1  gate597(.a(G528), .O(gate157inter8));
  nand2 gate598(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate599(.a(s_7), .b(gate157inter3), .O(gate157inter10));
  nor2  gate600(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate601(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate602(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1471(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1472(.a(gate159inter0), .b(s_132), .O(gate159inter1));
  and2  gate1473(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1474(.a(s_132), .O(gate159inter3));
  inv1  gate1475(.a(s_133), .O(gate159inter4));
  nand2 gate1476(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1477(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1478(.a(G444), .O(gate159inter7));
  inv1  gate1479(.a(G531), .O(gate159inter8));
  nand2 gate1480(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1481(.a(s_133), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1482(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1483(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1484(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2521(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2522(.a(gate165inter0), .b(s_282), .O(gate165inter1));
  and2  gate2523(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2524(.a(s_282), .O(gate165inter3));
  inv1  gate2525(.a(s_283), .O(gate165inter4));
  nand2 gate2526(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2527(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2528(.a(G462), .O(gate165inter7));
  inv1  gate2529(.a(G540), .O(gate165inter8));
  nand2 gate2530(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2531(.a(s_283), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2532(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2533(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2534(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2493(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2494(.a(gate169inter0), .b(s_278), .O(gate169inter1));
  and2  gate2495(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2496(.a(s_278), .O(gate169inter3));
  inv1  gate2497(.a(s_279), .O(gate169inter4));
  nand2 gate2498(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2499(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2500(.a(G474), .O(gate169inter7));
  inv1  gate2501(.a(G546), .O(gate169inter8));
  nand2 gate2502(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2503(.a(s_279), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2504(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2505(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2506(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2031(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2032(.a(gate171inter0), .b(s_212), .O(gate171inter1));
  and2  gate2033(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2034(.a(s_212), .O(gate171inter3));
  inv1  gate2035(.a(s_213), .O(gate171inter4));
  nand2 gate2036(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2037(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2038(.a(G480), .O(gate171inter7));
  inv1  gate2039(.a(G549), .O(gate171inter8));
  nand2 gate2040(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2041(.a(s_213), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2042(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2043(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2044(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1723(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1724(.a(gate173inter0), .b(s_168), .O(gate173inter1));
  and2  gate1725(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1726(.a(s_168), .O(gate173inter3));
  inv1  gate1727(.a(s_169), .O(gate173inter4));
  nand2 gate1728(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1729(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1730(.a(G486), .O(gate173inter7));
  inv1  gate1731(.a(G552), .O(gate173inter8));
  nand2 gate1732(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1733(.a(s_169), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1734(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1735(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1736(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1359(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1360(.a(gate181inter0), .b(s_116), .O(gate181inter1));
  and2  gate1361(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1362(.a(s_116), .O(gate181inter3));
  inv1  gate1363(.a(s_117), .O(gate181inter4));
  nand2 gate1364(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1365(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1366(.a(G510), .O(gate181inter7));
  inv1  gate1367(.a(G564), .O(gate181inter8));
  nand2 gate1368(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1369(.a(s_117), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1370(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1371(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1372(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1905(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1906(.a(gate182inter0), .b(s_194), .O(gate182inter1));
  and2  gate1907(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1908(.a(s_194), .O(gate182inter3));
  inv1  gate1909(.a(s_195), .O(gate182inter4));
  nand2 gate1910(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1911(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1912(.a(G513), .O(gate182inter7));
  inv1  gate1913(.a(G564), .O(gate182inter8));
  nand2 gate1914(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1915(.a(s_195), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1916(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1917(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1918(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate631(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate632(.a(gate187inter0), .b(s_12), .O(gate187inter1));
  and2  gate633(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate634(.a(s_12), .O(gate187inter3));
  inv1  gate635(.a(s_13), .O(gate187inter4));
  nand2 gate636(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate637(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate638(.a(G574), .O(gate187inter7));
  inv1  gate639(.a(G575), .O(gate187inter8));
  nand2 gate640(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate641(.a(s_13), .b(gate187inter3), .O(gate187inter10));
  nor2  gate642(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate643(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate644(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2129(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2130(.a(gate190inter0), .b(s_226), .O(gate190inter1));
  and2  gate2131(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2132(.a(s_226), .O(gate190inter3));
  inv1  gate2133(.a(s_227), .O(gate190inter4));
  nand2 gate2134(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2135(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2136(.a(G580), .O(gate190inter7));
  inv1  gate2137(.a(G581), .O(gate190inter8));
  nand2 gate2138(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2139(.a(s_227), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2140(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2141(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2142(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2227(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2228(.a(gate201inter0), .b(s_240), .O(gate201inter1));
  and2  gate2229(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2230(.a(s_240), .O(gate201inter3));
  inv1  gate2231(.a(s_241), .O(gate201inter4));
  nand2 gate2232(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2233(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2234(.a(G602), .O(gate201inter7));
  inv1  gate2235(.a(G607), .O(gate201inter8));
  nand2 gate2236(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2237(.a(s_241), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2238(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2239(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2240(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate715(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate716(.a(gate202inter0), .b(s_24), .O(gate202inter1));
  and2  gate717(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate718(.a(s_24), .O(gate202inter3));
  inv1  gate719(.a(s_25), .O(gate202inter4));
  nand2 gate720(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate721(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate722(.a(G612), .O(gate202inter7));
  inv1  gate723(.a(G617), .O(gate202inter8));
  nand2 gate724(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate725(.a(s_25), .b(gate202inter3), .O(gate202inter10));
  nor2  gate726(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate727(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate728(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1331(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1332(.a(gate204inter0), .b(s_112), .O(gate204inter1));
  and2  gate1333(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1334(.a(s_112), .O(gate204inter3));
  inv1  gate1335(.a(s_113), .O(gate204inter4));
  nand2 gate1336(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1337(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1338(.a(G607), .O(gate204inter7));
  inv1  gate1339(.a(G617), .O(gate204inter8));
  nand2 gate1340(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1341(.a(s_113), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1342(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1343(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1344(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate603(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate604(.a(gate207inter0), .b(s_8), .O(gate207inter1));
  and2  gate605(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate606(.a(s_8), .O(gate207inter3));
  inv1  gate607(.a(s_9), .O(gate207inter4));
  nand2 gate608(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate609(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate610(.a(G622), .O(gate207inter7));
  inv1  gate611(.a(G632), .O(gate207inter8));
  nand2 gate612(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate613(.a(s_9), .b(gate207inter3), .O(gate207inter10));
  nor2  gate614(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate615(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate616(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2423(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2424(.a(gate208inter0), .b(s_268), .O(gate208inter1));
  and2  gate2425(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2426(.a(s_268), .O(gate208inter3));
  inv1  gate2427(.a(s_269), .O(gate208inter4));
  nand2 gate2428(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2429(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2430(.a(G627), .O(gate208inter7));
  inv1  gate2431(.a(G637), .O(gate208inter8));
  nand2 gate2432(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2433(.a(s_269), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2434(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2435(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2436(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2045(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2046(.a(gate209inter0), .b(s_214), .O(gate209inter1));
  and2  gate2047(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2048(.a(s_214), .O(gate209inter3));
  inv1  gate2049(.a(s_215), .O(gate209inter4));
  nand2 gate2050(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2051(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2052(.a(G602), .O(gate209inter7));
  inv1  gate2053(.a(G666), .O(gate209inter8));
  nand2 gate2054(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2055(.a(s_215), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2056(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2057(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2058(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2297(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2298(.a(gate212inter0), .b(s_250), .O(gate212inter1));
  and2  gate2299(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2300(.a(s_250), .O(gate212inter3));
  inv1  gate2301(.a(s_251), .O(gate212inter4));
  nand2 gate2302(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2303(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2304(.a(G617), .O(gate212inter7));
  inv1  gate2305(.a(G669), .O(gate212inter8));
  nand2 gate2306(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2307(.a(s_251), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2308(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2309(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2310(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2255(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2256(.a(gate214inter0), .b(s_244), .O(gate214inter1));
  and2  gate2257(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2258(.a(s_244), .O(gate214inter3));
  inv1  gate2259(.a(s_245), .O(gate214inter4));
  nand2 gate2260(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2261(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2262(.a(G612), .O(gate214inter7));
  inv1  gate2263(.a(G672), .O(gate214inter8));
  nand2 gate2264(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2265(.a(s_245), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2266(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2267(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2268(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1345(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1346(.a(gate216inter0), .b(s_114), .O(gate216inter1));
  and2  gate1347(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1348(.a(s_114), .O(gate216inter3));
  inv1  gate1349(.a(s_115), .O(gate216inter4));
  nand2 gate1350(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1351(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1352(.a(G617), .O(gate216inter7));
  inv1  gate1353(.a(G675), .O(gate216inter8));
  nand2 gate1354(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1355(.a(s_115), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1356(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1357(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1358(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate757(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate758(.a(gate217inter0), .b(s_30), .O(gate217inter1));
  and2  gate759(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate760(.a(s_30), .O(gate217inter3));
  inv1  gate761(.a(s_31), .O(gate217inter4));
  nand2 gate762(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate763(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate764(.a(G622), .O(gate217inter7));
  inv1  gate765(.a(G678), .O(gate217inter8));
  nand2 gate766(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate767(.a(s_31), .b(gate217inter3), .O(gate217inter10));
  nor2  gate768(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate769(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate770(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1457(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1458(.a(gate220inter0), .b(s_130), .O(gate220inter1));
  and2  gate1459(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1460(.a(s_130), .O(gate220inter3));
  inv1  gate1461(.a(s_131), .O(gate220inter4));
  nand2 gate1462(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1463(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1464(.a(G637), .O(gate220inter7));
  inv1  gate1465(.a(G681), .O(gate220inter8));
  nand2 gate1466(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1467(.a(s_131), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1468(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1469(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1470(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1233(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1234(.a(gate221inter0), .b(s_98), .O(gate221inter1));
  and2  gate1235(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1236(.a(s_98), .O(gate221inter3));
  inv1  gate1237(.a(s_99), .O(gate221inter4));
  nand2 gate1238(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1239(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1240(.a(G622), .O(gate221inter7));
  inv1  gate1241(.a(G684), .O(gate221inter8));
  nand2 gate1242(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1243(.a(s_99), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1244(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1245(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1246(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1765(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1766(.a(gate224inter0), .b(s_174), .O(gate224inter1));
  and2  gate1767(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1768(.a(s_174), .O(gate224inter3));
  inv1  gate1769(.a(s_175), .O(gate224inter4));
  nand2 gate1770(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1771(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1772(.a(G637), .O(gate224inter7));
  inv1  gate1773(.a(G687), .O(gate224inter8));
  nand2 gate1774(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1775(.a(s_175), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1776(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1777(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1778(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1541(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1542(.a(gate227inter0), .b(s_142), .O(gate227inter1));
  and2  gate1543(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1544(.a(s_142), .O(gate227inter3));
  inv1  gate1545(.a(s_143), .O(gate227inter4));
  nand2 gate1546(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1547(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1548(.a(G694), .O(gate227inter7));
  inv1  gate1549(.a(G695), .O(gate227inter8));
  nand2 gate1550(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1551(.a(s_143), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1552(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1553(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1554(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate869(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate870(.a(gate230inter0), .b(s_46), .O(gate230inter1));
  and2  gate871(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate872(.a(s_46), .O(gate230inter3));
  inv1  gate873(.a(s_47), .O(gate230inter4));
  nand2 gate874(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate875(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate876(.a(G700), .O(gate230inter7));
  inv1  gate877(.a(G701), .O(gate230inter8));
  nand2 gate878(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate879(.a(s_47), .b(gate230inter3), .O(gate230inter10));
  nor2  gate880(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate881(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate882(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1415(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1416(.a(gate234inter0), .b(s_124), .O(gate234inter1));
  and2  gate1417(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1418(.a(s_124), .O(gate234inter3));
  inv1  gate1419(.a(s_125), .O(gate234inter4));
  nand2 gate1420(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1421(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1422(.a(G245), .O(gate234inter7));
  inv1  gate1423(.a(G721), .O(gate234inter8));
  nand2 gate1424(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1425(.a(s_125), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1426(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1427(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1428(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate981(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate982(.a(gate241inter0), .b(s_62), .O(gate241inter1));
  and2  gate983(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate984(.a(s_62), .O(gate241inter3));
  inv1  gate985(.a(s_63), .O(gate241inter4));
  nand2 gate986(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate987(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate988(.a(G242), .O(gate241inter7));
  inv1  gate989(.a(G730), .O(gate241inter8));
  nand2 gate990(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate991(.a(s_63), .b(gate241inter3), .O(gate241inter10));
  nor2  gate992(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate993(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate994(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1275(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1276(.a(gate243inter0), .b(s_104), .O(gate243inter1));
  and2  gate1277(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1278(.a(s_104), .O(gate243inter3));
  inv1  gate1279(.a(s_105), .O(gate243inter4));
  nand2 gate1280(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1281(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1282(.a(G245), .O(gate243inter7));
  inv1  gate1283(.a(G733), .O(gate243inter8));
  nand2 gate1284(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1285(.a(s_105), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1286(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1287(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1288(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate743(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate744(.a(gate244inter0), .b(s_28), .O(gate244inter1));
  and2  gate745(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate746(.a(s_28), .O(gate244inter3));
  inv1  gate747(.a(s_29), .O(gate244inter4));
  nand2 gate748(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate749(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate750(.a(G721), .O(gate244inter7));
  inv1  gate751(.a(G733), .O(gate244inter8));
  nand2 gate752(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate753(.a(s_29), .b(gate244inter3), .O(gate244inter10));
  nor2  gate754(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate755(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate756(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1835(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1836(.a(gate246inter0), .b(s_184), .O(gate246inter1));
  and2  gate1837(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1838(.a(s_184), .O(gate246inter3));
  inv1  gate1839(.a(s_185), .O(gate246inter4));
  nand2 gate1840(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1841(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1842(.a(G724), .O(gate246inter7));
  inv1  gate1843(.a(G736), .O(gate246inter8));
  nand2 gate1844(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1845(.a(s_185), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1846(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1847(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1848(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate673(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate674(.a(gate247inter0), .b(s_18), .O(gate247inter1));
  and2  gate675(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate676(.a(s_18), .O(gate247inter3));
  inv1  gate677(.a(s_19), .O(gate247inter4));
  nand2 gate678(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate679(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate680(.a(G251), .O(gate247inter7));
  inv1  gate681(.a(G739), .O(gate247inter8));
  nand2 gate682(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate683(.a(s_19), .b(gate247inter3), .O(gate247inter10));
  nor2  gate684(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate685(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate686(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1317(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1318(.a(gate248inter0), .b(s_110), .O(gate248inter1));
  and2  gate1319(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1320(.a(s_110), .O(gate248inter3));
  inv1  gate1321(.a(s_111), .O(gate248inter4));
  nand2 gate1322(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1323(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1324(.a(G727), .O(gate248inter7));
  inv1  gate1325(.a(G739), .O(gate248inter8));
  nand2 gate1326(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1327(.a(s_111), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1328(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1329(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1330(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1387(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1388(.a(gate250inter0), .b(s_120), .O(gate250inter1));
  and2  gate1389(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1390(.a(s_120), .O(gate250inter3));
  inv1  gate1391(.a(s_121), .O(gate250inter4));
  nand2 gate1392(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1393(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1394(.a(G706), .O(gate250inter7));
  inv1  gate1395(.a(G742), .O(gate250inter8));
  nand2 gate1396(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1397(.a(s_121), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1398(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1399(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1400(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1149(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1150(.a(gate252inter0), .b(s_86), .O(gate252inter1));
  and2  gate1151(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1152(.a(s_86), .O(gate252inter3));
  inv1  gate1153(.a(s_87), .O(gate252inter4));
  nand2 gate1154(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1155(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1156(.a(G709), .O(gate252inter7));
  inv1  gate1157(.a(G745), .O(gate252inter8));
  nand2 gate1158(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1159(.a(s_87), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1160(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1161(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1162(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate841(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate842(.a(gate254inter0), .b(s_42), .O(gate254inter1));
  and2  gate843(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate844(.a(s_42), .O(gate254inter3));
  inv1  gate845(.a(s_43), .O(gate254inter4));
  nand2 gate846(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate847(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate848(.a(G712), .O(gate254inter7));
  inv1  gate849(.a(G748), .O(gate254inter8));
  nand2 gate850(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate851(.a(s_43), .b(gate254inter3), .O(gate254inter10));
  nor2  gate852(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate853(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate854(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1961(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1962(.a(gate255inter0), .b(s_202), .O(gate255inter1));
  and2  gate1963(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1964(.a(s_202), .O(gate255inter3));
  inv1  gate1965(.a(s_203), .O(gate255inter4));
  nand2 gate1966(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1967(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1968(.a(G263), .O(gate255inter7));
  inv1  gate1969(.a(G751), .O(gate255inter8));
  nand2 gate1970(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1971(.a(s_203), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1972(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1973(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1974(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2619(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2620(.a(gate258inter0), .b(s_296), .O(gate258inter1));
  and2  gate2621(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2622(.a(s_296), .O(gate258inter3));
  inv1  gate2623(.a(s_297), .O(gate258inter4));
  nand2 gate2624(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2625(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2626(.a(G756), .O(gate258inter7));
  inv1  gate2627(.a(G757), .O(gate258inter8));
  nand2 gate2628(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2629(.a(s_297), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2630(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2631(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2632(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate2185(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2186(.a(gate260inter0), .b(s_234), .O(gate260inter1));
  and2  gate2187(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2188(.a(s_234), .O(gate260inter3));
  inv1  gate2189(.a(s_235), .O(gate260inter4));
  nand2 gate2190(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2191(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2192(.a(G760), .O(gate260inter7));
  inv1  gate2193(.a(G761), .O(gate260inter8));
  nand2 gate2194(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2195(.a(s_235), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2196(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2197(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2198(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2577(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2578(.a(gate261inter0), .b(s_290), .O(gate261inter1));
  and2  gate2579(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2580(.a(s_290), .O(gate261inter3));
  inv1  gate2581(.a(s_291), .O(gate261inter4));
  nand2 gate2582(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2583(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2584(.a(G762), .O(gate261inter7));
  inv1  gate2585(.a(G763), .O(gate261inter8));
  nand2 gate2586(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2587(.a(s_291), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2588(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2589(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2590(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1037(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1038(.a(gate267inter0), .b(s_70), .O(gate267inter1));
  and2  gate1039(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1040(.a(s_70), .O(gate267inter3));
  inv1  gate1041(.a(s_71), .O(gate267inter4));
  nand2 gate1042(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1043(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1044(.a(G648), .O(gate267inter7));
  inv1  gate1045(.a(G776), .O(gate267inter8));
  nand2 gate1046(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1047(.a(s_71), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1048(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1049(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1050(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1261(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1262(.a(gate269inter0), .b(s_102), .O(gate269inter1));
  and2  gate1263(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1264(.a(s_102), .O(gate269inter3));
  inv1  gate1265(.a(s_103), .O(gate269inter4));
  nand2 gate1266(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1267(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1268(.a(G654), .O(gate269inter7));
  inv1  gate1269(.a(G782), .O(gate269inter8));
  nand2 gate1270(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1271(.a(s_103), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1272(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1273(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1274(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate785(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate786(.a(gate271inter0), .b(s_34), .O(gate271inter1));
  and2  gate787(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate788(.a(s_34), .O(gate271inter3));
  inv1  gate789(.a(s_35), .O(gate271inter4));
  nand2 gate790(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate791(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate792(.a(G660), .O(gate271inter7));
  inv1  gate793(.a(G788), .O(gate271inter8));
  nand2 gate794(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate795(.a(s_35), .b(gate271inter3), .O(gate271inter10));
  nor2  gate796(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate797(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate798(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate701(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate702(.a(gate277inter0), .b(s_22), .O(gate277inter1));
  and2  gate703(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate704(.a(s_22), .O(gate277inter3));
  inv1  gate705(.a(s_23), .O(gate277inter4));
  nand2 gate706(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate707(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate708(.a(G648), .O(gate277inter7));
  inv1  gate709(.a(G800), .O(gate277inter8));
  nand2 gate710(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate711(.a(s_23), .b(gate277inter3), .O(gate277inter10));
  nor2  gate712(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate713(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate714(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1667(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1668(.a(gate278inter0), .b(s_160), .O(gate278inter1));
  and2  gate1669(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1670(.a(s_160), .O(gate278inter3));
  inv1  gate1671(.a(s_161), .O(gate278inter4));
  nand2 gate1672(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1673(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1674(.a(G776), .O(gate278inter7));
  inv1  gate1675(.a(G800), .O(gate278inter8));
  nand2 gate1676(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1677(.a(s_161), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1678(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1679(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1680(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate925(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate926(.a(gate279inter0), .b(s_54), .O(gate279inter1));
  and2  gate927(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate928(.a(s_54), .O(gate279inter3));
  inv1  gate929(.a(s_55), .O(gate279inter4));
  nand2 gate930(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate931(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate932(.a(G651), .O(gate279inter7));
  inv1  gate933(.a(G803), .O(gate279inter8));
  nand2 gate934(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate935(.a(s_55), .b(gate279inter3), .O(gate279inter10));
  nor2  gate936(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate937(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate938(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2605(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2606(.a(gate281inter0), .b(s_294), .O(gate281inter1));
  and2  gate2607(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2608(.a(s_294), .O(gate281inter3));
  inv1  gate2609(.a(s_295), .O(gate281inter4));
  nand2 gate2610(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2611(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2612(.a(G654), .O(gate281inter7));
  inv1  gate2613(.a(G806), .O(gate281inter8));
  nand2 gate2614(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2615(.a(s_295), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2616(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2617(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2618(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1429(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1430(.a(gate283inter0), .b(s_126), .O(gate283inter1));
  and2  gate1431(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1432(.a(s_126), .O(gate283inter3));
  inv1  gate1433(.a(s_127), .O(gate283inter4));
  nand2 gate1434(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1435(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1436(.a(G657), .O(gate283inter7));
  inv1  gate1437(.a(G809), .O(gate283inter8));
  nand2 gate1438(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1439(.a(s_127), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1440(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1441(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1442(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2549(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2550(.a(gate289inter0), .b(s_286), .O(gate289inter1));
  and2  gate2551(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2552(.a(s_286), .O(gate289inter3));
  inv1  gate2553(.a(s_287), .O(gate289inter4));
  nand2 gate2554(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2555(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2556(.a(G818), .O(gate289inter7));
  inv1  gate2557(.a(G819), .O(gate289inter8));
  nand2 gate2558(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2559(.a(s_287), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2560(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2561(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2562(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1443(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1444(.a(gate292inter0), .b(s_128), .O(gate292inter1));
  and2  gate1445(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1446(.a(s_128), .O(gate292inter3));
  inv1  gate1447(.a(s_129), .O(gate292inter4));
  nand2 gate1448(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1449(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1450(.a(G824), .O(gate292inter7));
  inv1  gate1451(.a(G825), .O(gate292inter8));
  nand2 gate1452(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1453(.a(s_129), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1454(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1455(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1456(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate953(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate954(.a(gate293inter0), .b(s_58), .O(gate293inter1));
  and2  gate955(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate956(.a(s_58), .O(gate293inter3));
  inv1  gate957(.a(s_59), .O(gate293inter4));
  nand2 gate958(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate959(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate960(.a(G828), .O(gate293inter7));
  inv1  gate961(.a(G829), .O(gate293inter8));
  nand2 gate962(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate963(.a(s_59), .b(gate293inter3), .O(gate293inter10));
  nor2  gate964(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate965(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate966(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1947(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1948(.a(gate295inter0), .b(s_200), .O(gate295inter1));
  and2  gate1949(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1950(.a(s_200), .O(gate295inter3));
  inv1  gate1951(.a(s_201), .O(gate295inter4));
  nand2 gate1952(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1953(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1954(.a(G830), .O(gate295inter7));
  inv1  gate1955(.a(G831), .O(gate295inter8));
  nand2 gate1956(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1957(.a(s_201), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1958(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1959(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1960(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1009(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1010(.a(gate393inter0), .b(s_66), .O(gate393inter1));
  and2  gate1011(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1012(.a(s_66), .O(gate393inter3));
  inv1  gate1013(.a(s_67), .O(gate393inter4));
  nand2 gate1014(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1015(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1016(.a(G7), .O(gate393inter7));
  inv1  gate1017(.a(G1054), .O(gate393inter8));
  nand2 gate1018(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1019(.a(s_67), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1020(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1021(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1022(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1485(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1486(.a(gate397inter0), .b(s_134), .O(gate397inter1));
  and2  gate1487(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1488(.a(s_134), .O(gate397inter3));
  inv1  gate1489(.a(s_135), .O(gate397inter4));
  nand2 gate1490(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1491(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1492(.a(G11), .O(gate397inter7));
  inv1  gate1493(.a(G1066), .O(gate397inter8));
  nand2 gate1494(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1495(.a(s_135), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1496(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1497(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1498(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2101(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2102(.a(gate398inter0), .b(s_222), .O(gate398inter1));
  and2  gate2103(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2104(.a(s_222), .O(gate398inter3));
  inv1  gate2105(.a(s_223), .O(gate398inter4));
  nand2 gate2106(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2107(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2108(.a(G12), .O(gate398inter7));
  inv1  gate2109(.a(G1069), .O(gate398inter8));
  nand2 gate2110(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2111(.a(s_223), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2112(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2113(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2114(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2507(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2508(.a(gate401inter0), .b(s_280), .O(gate401inter1));
  and2  gate2509(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2510(.a(s_280), .O(gate401inter3));
  inv1  gate2511(.a(s_281), .O(gate401inter4));
  nand2 gate2512(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2513(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2514(.a(G15), .O(gate401inter7));
  inv1  gate2515(.a(G1078), .O(gate401inter8));
  nand2 gate2516(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2517(.a(s_281), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2518(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2519(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2520(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate855(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate856(.a(gate404inter0), .b(s_44), .O(gate404inter1));
  and2  gate857(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate858(.a(s_44), .O(gate404inter3));
  inv1  gate859(.a(s_45), .O(gate404inter4));
  nand2 gate860(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate861(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate862(.a(G18), .O(gate404inter7));
  inv1  gate863(.a(G1087), .O(gate404inter8));
  nand2 gate864(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate865(.a(s_45), .b(gate404inter3), .O(gate404inter10));
  nor2  gate866(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate867(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate868(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate827(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate828(.a(gate405inter0), .b(s_40), .O(gate405inter1));
  and2  gate829(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate830(.a(s_40), .O(gate405inter3));
  inv1  gate831(.a(s_41), .O(gate405inter4));
  nand2 gate832(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate833(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate834(.a(G19), .O(gate405inter7));
  inv1  gate835(.a(G1090), .O(gate405inter8));
  nand2 gate836(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate837(.a(s_41), .b(gate405inter3), .O(gate405inter10));
  nor2  gate838(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate839(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate840(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1177(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1178(.a(gate406inter0), .b(s_90), .O(gate406inter1));
  and2  gate1179(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1180(.a(s_90), .O(gate406inter3));
  inv1  gate1181(.a(s_91), .O(gate406inter4));
  nand2 gate1182(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1183(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1184(.a(G20), .O(gate406inter7));
  inv1  gate1185(.a(G1093), .O(gate406inter8));
  nand2 gate1186(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1187(.a(s_91), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1188(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1189(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1190(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate2465(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2466(.a(gate407inter0), .b(s_274), .O(gate407inter1));
  and2  gate2467(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2468(.a(s_274), .O(gate407inter3));
  inv1  gate2469(.a(s_275), .O(gate407inter4));
  nand2 gate2470(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2471(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2472(.a(G21), .O(gate407inter7));
  inv1  gate2473(.a(G1096), .O(gate407inter8));
  nand2 gate2474(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2475(.a(s_275), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2476(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2477(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2478(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate2395(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2396(.a(gate408inter0), .b(s_264), .O(gate408inter1));
  and2  gate2397(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2398(.a(s_264), .O(gate408inter3));
  inv1  gate2399(.a(s_265), .O(gate408inter4));
  nand2 gate2400(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2401(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2402(.a(G22), .O(gate408inter7));
  inv1  gate2403(.a(G1099), .O(gate408inter8));
  nand2 gate2404(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2405(.a(s_265), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2406(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2407(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2408(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1681(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1682(.a(gate416inter0), .b(s_162), .O(gate416inter1));
  and2  gate1683(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1684(.a(s_162), .O(gate416inter3));
  inv1  gate1685(.a(s_163), .O(gate416inter4));
  nand2 gate1686(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1687(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1688(.a(G30), .O(gate416inter7));
  inv1  gate1689(.a(G1123), .O(gate416inter8));
  nand2 gate1690(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1691(.a(s_163), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1692(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1693(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1694(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2409(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2410(.a(gate417inter0), .b(s_266), .O(gate417inter1));
  and2  gate2411(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2412(.a(s_266), .O(gate417inter3));
  inv1  gate2413(.a(s_267), .O(gate417inter4));
  nand2 gate2414(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2415(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2416(.a(G31), .O(gate417inter7));
  inv1  gate2417(.a(G1126), .O(gate417inter8));
  nand2 gate2418(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2419(.a(s_267), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2420(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2421(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2422(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1737(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1738(.a(gate419inter0), .b(s_170), .O(gate419inter1));
  and2  gate1739(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1740(.a(s_170), .O(gate419inter3));
  inv1  gate1741(.a(s_171), .O(gate419inter4));
  nand2 gate1742(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1743(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1744(.a(G1), .O(gate419inter7));
  inv1  gate1745(.a(G1132), .O(gate419inter8));
  nand2 gate1746(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1747(.a(s_171), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1748(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1749(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1750(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2017(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2018(.a(gate420inter0), .b(s_210), .O(gate420inter1));
  and2  gate2019(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2020(.a(s_210), .O(gate420inter3));
  inv1  gate2021(.a(s_211), .O(gate420inter4));
  nand2 gate2022(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2023(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2024(.a(G1036), .O(gate420inter7));
  inv1  gate2025(.a(G1132), .O(gate420inter8));
  nand2 gate2026(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2027(.a(s_211), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2028(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2029(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2030(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1093(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1094(.a(gate424inter0), .b(s_78), .O(gate424inter1));
  and2  gate1095(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1096(.a(s_78), .O(gate424inter3));
  inv1  gate1097(.a(s_79), .O(gate424inter4));
  nand2 gate1098(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1099(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1100(.a(G1042), .O(gate424inter7));
  inv1  gate1101(.a(G1138), .O(gate424inter8));
  nand2 gate1102(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1103(.a(s_79), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1104(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1105(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1106(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1611(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1612(.a(gate425inter0), .b(s_152), .O(gate425inter1));
  and2  gate1613(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1614(.a(s_152), .O(gate425inter3));
  inv1  gate1615(.a(s_153), .O(gate425inter4));
  nand2 gate1616(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1617(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1618(.a(G4), .O(gate425inter7));
  inv1  gate1619(.a(G1141), .O(gate425inter8));
  nand2 gate1620(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1621(.a(s_153), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1622(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1623(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1624(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate617(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate618(.a(gate426inter0), .b(s_10), .O(gate426inter1));
  and2  gate619(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate620(.a(s_10), .O(gate426inter3));
  inv1  gate621(.a(s_11), .O(gate426inter4));
  nand2 gate622(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate623(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate624(.a(G1045), .O(gate426inter7));
  inv1  gate625(.a(G1141), .O(gate426inter8));
  nand2 gate626(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate627(.a(s_11), .b(gate426inter3), .O(gate426inter10));
  nor2  gate628(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate629(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate630(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2535(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2536(.a(gate427inter0), .b(s_284), .O(gate427inter1));
  and2  gate2537(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2538(.a(s_284), .O(gate427inter3));
  inv1  gate2539(.a(s_285), .O(gate427inter4));
  nand2 gate2540(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2541(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2542(.a(G5), .O(gate427inter7));
  inv1  gate2543(.a(G1144), .O(gate427inter8));
  nand2 gate2544(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2545(.a(s_285), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2546(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2547(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2548(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate2381(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2382(.a(gate436inter0), .b(s_262), .O(gate436inter1));
  and2  gate2383(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2384(.a(s_262), .O(gate436inter3));
  inv1  gate2385(.a(s_263), .O(gate436inter4));
  nand2 gate2386(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2387(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2388(.a(G1060), .O(gate436inter7));
  inv1  gate2389(.a(G1156), .O(gate436inter8));
  nand2 gate2390(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2391(.a(s_263), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2392(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2393(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2394(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1205(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1206(.a(gate442inter0), .b(s_94), .O(gate442inter1));
  and2  gate1207(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1208(.a(s_94), .O(gate442inter3));
  inv1  gate1209(.a(s_95), .O(gate442inter4));
  nand2 gate1210(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1211(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1212(.a(G1069), .O(gate442inter7));
  inv1  gate1213(.a(G1165), .O(gate442inter8));
  nand2 gate1214(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1215(.a(s_95), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1216(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1217(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1218(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2171(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2172(.a(gate452inter0), .b(s_232), .O(gate452inter1));
  and2  gate2173(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2174(.a(s_232), .O(gate452inter3));
  inv1  gate2175(.a(s_233), .O(gate452inter4));
  nand2 gate2176(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2177(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2178(.a(G1084), .O(gate452inter7));
  inv1  gate2179(.a(G1180), .O(gate452inter8));
  nand2 gate2180(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2181(.a(s_233), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2182(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2183(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2184(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1401(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1402(.a(gate454inter0), .b(s_122), .O(gate454inter1));
  and2  gate1403(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1404(.a(s_122), .O(gate454inter3));
  inv1  gate1405(.a(s_123), .O(gate454inter4));
  nand2 gate1406(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1407(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1408(.a(G1087), .O(gate454inter7));
  inv1  gate1409(.a(G1183), .O(gate454inter8));
  nand2 gate1410(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1411(.a(s_123), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1412(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1413(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1414(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1989(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1990(.a(gate457inter0), .b(s_206), .O(gate457inter1));
  and2  gate1991(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1992(.a(s_206), .O(gate457inter3));
  inv1  gate1993(.a(s_207), .O(gate457inter4));
  nand2 gate1994(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1995(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1996(.a(G20), .O(gate457inter7));
  inv1  gate1997(.a(G1189), .O(gate457inter8));
  nand2 gate1998(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1999(.a(s_207), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2000(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2001(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2002(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1891(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1892(.a(gate458inter0), .b(s_192), .O(gate458inter1));
  and2  gate1893(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1894(.a(s_192), .O(gate458inter3));
  inv1  gate1895(.a(s_193), .O(gate458inter4));
  nand2 gate1896(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1897(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1898(.a(G1093), .O(gate458inter7));
  inv1  gate1899(.a(G1189), .O(gate458inter8));
  nand2 gate1900(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1901(.a(s_193), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1902(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1903(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1904(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate2199(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2200(.a(gate459inter0), .b(s_236), .O(gate459inter1));
  and2  gate2201(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2202(.a(s_236), .O(gate459inter3));
  inv1  gate2203(.a(s_237), .O(gate459inter4));
  nand2 gate2204(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2205(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2206(.a(G21), .O(gate459inter7));
  inv1  gate2207(.a(G1192), .O(gate459inter8));
  nand2 gate2208(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2209(.a(s_237), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2210(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2211(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2212(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1527(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1528(.a(gate463inter0), .b(s_140), .O(gate463inter1));
  and2  gate1529(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1530(.a(s_140), .O(gate463inter3));
  inv1  gate1531(.a(s_141), .O(gate463inter4));
  nand2 gate1532(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1533(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1534(.a(G23), .O(gate463inter7));
  inv1  gate1535(.a(G1198), .O(gate463inter8));
  nand2 gate1536(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1537(.a(s_141), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1538(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1539(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1540(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate729(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate730(.a(gate464inter0), .b(s_26), .O(gate464inter1));
  and2  gate731(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate732(.a(s_26), .O(gate464inter3));
  inv1  gate733(.a(s_27), .O(gate464inter4));
  nand2 gate734(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate735(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate736(.a(G1102), .O(gate464inter7));
  inv1  gate737(.a(G1198), .O(gate464inter8));
  nand2 gate738(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate739(.a(s_27), .b(gate464inter3), .O(gate464inter10));
  nor2  gate740(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate741(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate742(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate687(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate688(.a(gate470inter0), .b(s_20), .O(gate470inter1));
  and2  gate689(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate690(.a(s_20), .O(gate470inter3));
  inv1  gate691(.a(s_21), .O(gate470inter4));
  nand2 gate692(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate693(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate694(.a(G1111), .O(gate470inter7));
  inv1  gate695(.a(G1207), .O(gate470inter8));
  nand2 gate696(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate697(.a(s_21), .b(gate470inter3), .O(gate470inter10));
  nor2  gate698(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate699(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate700(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1695(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1696(.a(gate473inter0), .b(s_164), .O(gate473inter1));
  and2  gate1697(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1698(.a(s_164), .O(gate473inter3));
  inv1  gate1699(.a(s_165), .O(gate473inter4));
  nand2 gate1700(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1701(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1702(.a(G28), .O(gate473inter7));
  inv1  gate1703(.a(G1213), .O(gate473inter8));
  nand2 gate1704(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1705(.a(s_165), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1706(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1707(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1708(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1569(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1570(.a(gate475inter0), .b(s_146), .O(gate475inter1));
  and2  gate1571(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1572(.a(s_146), .O(gate475inter3));
  inv1  gate1573(.a(s_147), .O(gate475inter4));
  nand2 gate1574(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1575(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1576(.a(G29), .O(gate475inter7));
  inv1  gate1577(.a(G1216), .O(gate475inter8));
  nand2 gate1578(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1579(.a(s_147), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1580(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1581(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1582(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2087(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2088(.a(gate476inter0), .b(s_220), .O(gate476inter1));
  and2  gate2089(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2090(.a(s_220), .O(gate476inter3));
  inv1  gate2091(.a(s_221), .O(gate476inter4));
  nand2 gate2092(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2093(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2094(.a(G1120), .O(gate476inter7));
  inv1  gate2095(.a(G1216), .O(gate476inter8));
  nand2 gate2096(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2097(.a(s_221), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2098(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2099(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2100(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate2339(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2340(.a(gate477inter0), .b(s_256), .O(gate477inter1));
  and2  gate2341(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2342(.a(s_256), .O(gate477inter3));
  inv1  gate2343(.a(s_257), .O(gate477inter4));
  nand2 gate2344(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2345(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2346(.a(G30), .O(gate477inter7));
  inv1  gate2347(.a(G1219), .O(gate477inter8));
  nand2 gate2348(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2349(.a(s_257), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2350(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2351(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2352(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1513(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1514(.a(gate479inter0), .b(s_138), .O(gate479inter1));
  and2  gate1515(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1516(.a(s_138), .O(gate479inter3));
  inv1  gate1517(.a(s_139), .O(gate479inter4));
  nand2 gate1518(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1519(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1520(.a(G31), .O(gate479inter7));
  inv1  gate1521(.a(G1222), .O(gate479inter8));
  nand2 gate1522(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1523(.a(s_139), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1524(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1525(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1526(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1807(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1808(.a(gate480inter0), .b(s_180), .O(gate480inter1));
  and2  gate1809(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1810(.a(s_180), .O(gate480inter3));
  inv1  gate1811(.a(s_181), .O(gate480inter4));
  nand2 gate1812(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1813(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1814(.a(G1126), .O(gate480inter7));
  inv1  gate1815(.a(G1222), .O(gate480inter8));
  nand2 gate1816(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1817(.a(s_181), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1818(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1819(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1820(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1191(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1192(.a(gate481inter0), .b(s_92), .O(gate481inter1));
  and2  gate1193(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1194(.a(s_92), .O(gate481inter3));
  inv1  gate1195(.a(s_93), .O(gate481inter4));
  nand2 gate1196(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1197(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1198(.a(G32), .O(gate481inter7));
  inv1  gate1199(.a(G1225), .O(gate481inter8));
  nand2 gate1200(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1201(.a(s_93), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1202(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1203(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1204(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1219(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1220(.a(gate491inter0), .b(s_96), .O(gate491inter1));
  and2  gate1221(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1222(.a(s_96), .O(gate491inter3));
  inv1  gate1223(.a(s_97), .O(gate491inter4));
  nand2 gate1224(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1225(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1226(.a(G1244), .O(gate491inter7));
  inv1  gate1227(.a(G1245), .O(gate491inter8));
  nand2 gate1228(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1229(.a(s_97), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1230(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1231(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1232(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1555(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1556(.a(gate492inter0), .b(s_144), .O(gate492inter1));
  and2  gate1557(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1558(.a(s_144), .O(gate492inter3));
  inv1  gate1559(.a(s_145), .O(gate492inter4));
  nand2 gate1560(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1561(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1562(.a(G1246), .O(gate492inter7));
  inv1  gate1563(.a(G1247), .O(gate492inter8));
  nand2 gate1564(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1565(.a(s_145), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1566(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1567(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1568(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate2003(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2004(.a(gate494inter0), .b(s_208), .O(gate494inter1));
  and2  gate2005(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2006(.a(s_208), .O(gate494inter3));
  inv1  gate2007(.a(s_209), .O(gate494inter4));
  nand2 gate2008(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2009(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2010(.a(G1250), .O(gate494inter7));
  inv1  gate2011(.a(G1251), .O(gate494inter8));
  nand2 gate2012(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2013(.a(s_209), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2014(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2015(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2016(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2241(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2242(.a(gate495inter0), .b(s_242), .O(gate495inter1));
  and2  gate2243(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2244(.a(s_242), .O(gate495inter3));
  inv1  gate2245(.a(s_243), .O(gate495inter4));
  nand2 gate2246(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2247(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2248(.a(G1252), .O(gate495inter7));
  inv1  gate2249(.a(G1253), .O(gate495inter8));
  nand2 gate2250(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2251(.a(s_243), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2252(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2253(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2254(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate967(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate968(.a(gate497inter0), .b(s_60), .O(gate497inter1));
  and2  gate969(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate970(.a(s_60), .O(gate497inter3));
  inv1  gate971(.a(s_61), .O(gate497inter4));
  nand2 gate972(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate973(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate974(.a(G1256), .O(gate497inter7));
  inv1  gate975(.a(G1257), .O(gate497inter8));
  nand2 gate976(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate977(.a(s_61), .b(gate497inter3), .O(gate497inter10));
  nor2  gate978(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate979(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate980(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1877(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1878(.a(gate498inter0), .b(s_190), .O(gate498inter1));
  and2  gate1879(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1880(.a(s_190), .O(gate498inter3));
  inv1  gate1881(.a(s_191), .O(gate498inter4));
  nand2 gate1882(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1883(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1884(.a(G1258), .O(gate498inter7));
  inv1  gate1885(.a(G1259), .O(gate498inter8));
  nand2 gate1886(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1887(.a(s_191), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1888(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1889(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1890(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2325(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2326(.a(gate501inter0), .b(s_254), .O(gate501inter1));
  and2  gate2327(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2328(.a(s_254), .O(gate501inter3));
  inv1  gate2329(.a(s_255), .O(gate501inter4));
  nand2 gate2330(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2331(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2332(.a(G1264), .O(gate501inter7));
  inv1  gate2333(.a(G1265), .O(gate501inter8));
  nand2 gate2334(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2335(.a(s_255), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2336(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2337(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2338(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1583(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1584(.a(gate506inter0), .b(s_148), .O(gate506inter1));
  and2  gate1585(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1586(.a(s_148), .O(gate506inter3));
  inv1  gate1587(.a(s_149), .O(gate506inter4));
  nand2 gate1588(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1589(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1590(.a(G1274), .O(gate506inter7));
  inv1  gate1591(.a(G1275), .O(gate506inter8));
  nand2 gate1592(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1593(.a(s_149), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1594(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1595(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1596(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate645(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate646(.a(gate509inter0), .b(s_14), .O(gate509inter1));
  and2  gate647(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate648(.a(s_14), .O(gate509inter3));
  inv1  gate649(.a(s_15), .O(gate509inter4));
  nand2 gate650(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate651(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate652(.a(G1280), .O(gate509inter7));
  inv1  gate653(.a(G1281), .O(gate509inter8));
  nand2 gate654(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate655(.a(s_15), .b(gate509inter3), .O(gate509inter10));
  nor2  gate656(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate657(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate658(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate911(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate912(.a(gate511inter0), .b(s_52), .O(gate511inter1));
  and2  gate913(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate914(.a(s_52), .O(gate511inter3));
  inv1  gate915(.a(s_53), .O(gate511inter4));
  nand2 gate916(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate917(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate918(.a(G1284), .O(gate511inter7));
  inv1  gate919(.a(G1285), .O(gate511inter8));
  nand2 gate920(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate921(.a(s_53), .b(gate511inter3), .O(gate511inter10));
  nor2  gate922(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate923(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate924(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule