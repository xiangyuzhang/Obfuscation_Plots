module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2017(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2018(.a(gate9inter0), .b(s_210), .O(gate9inter1));
  and2  gate2019(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2020(.a(s_210), .O(gate9inter3));
  inv1  gate2021(.a(s_211), .O(gate9inter4));
  nand2 gate2022(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2023(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2024(.a(G1), .O(gate9inter7));
  inv1  gate2025(.a(G2), .O(gate9inter8));
  nand2 gate2026(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2027(.a(s_211), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2028(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2029(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2030(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2367(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2368(.a(gate10inter0), .b(s_260), .O(gate10inter1));
  and2  gate2369(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2370(.a(s_260), .O(gate10inter3));
  inv1  gate2371(.a(s_261), .O(gate10inter4));
  nand2 gate2372(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2373(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2374(.a(G3), .O(gate10inter7));
  inv1  gate2375(.a(G4), .O(gate10inter8));
  nand2 gate2376(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2377(.a(s_261), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2378(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2379(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2380(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate561(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate562(.a(gate13inter0), .b(s_2), .O(gate13inter1));
  and2  gate563(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate564(.a(s_2), .O(gate13inter3));
  inv1  gate565(.a(s_3), .O(gate13inter4));
  nand2 gate566(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate567(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate568(.a(G9), .O(gate13inter7));
  inv1  gate569(.a(G10), .O(gate13inter8));
  nand2 gate570(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate571(.a(s_3), .b(gate13inter3), .O(gate13inter10));
  nor2  gate572(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate573(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate574(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1975(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1976(.a(gate14inter0), .b(s_204), .O(gate14inter1));
  and2  gate1977(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1978(.a(s_204), .O(gate14inter3));
  inv1  gate1979(.a(s_205), .O(gate14inter4));
  nand2 gate1980(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1981(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1982(.a(G11), .O(gate14inter7));
  inv1  gate1983(.a(G12), .O(gate14inter8));
  nand2 gate1984(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1985(.a(s_205), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1986(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1987(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1988(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1023(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1024(.a(gate16inter0), .b(s_68), .O(gate16inter1));
  and2  gate1025(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1026(.a(s_68), .O(gate16inter3));
  inv1  gate1027(.a(s_69), .O(gate16inter4));
  nand2 gate1028(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1029(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1030(.a(G15), .O(gate16inter7));
  inv1  gate1031(.a(G16), .O(gate16inter8));
  nand2 gate1032(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1033(.a(s_69), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1034(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1035(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1036(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate631(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate632(.a(gate17inter0), .b(s_12), .O(gate17inter1));
  and2  gate633(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate634(.a(s_12), .O(gate17inter3));
  inv1  gate635(.a(s_13), .O(gate17inter4));
  nand2 gate636(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate637(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate638(.a(G17), .O(gate17inter7));
  inv1  gate639(.a(G18), .O(gate17inter8));
  nand2 gate640(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate641(.a(s_13), .b(gate17inter3), .O(gate17inter10));
  nor2  gate642(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate643(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate644(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate2997(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2998(.a(gate18inter0), .b(s_350), .O(gate18inter1));
  and2  gate2999(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate3000(.a(s_350), .O(gate18inter3));
  inv1  gate3001(.a(s_351), .O(gate18inter4));
  nand2 gate3002(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate3003(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate3004(.a(G19), .O(gate18inter7));
  inv1  gate3005(.a(G20), .O(gate18inter8));
  nand2 gate3006(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate3007(.a(s_351), .b(gate18inter3), .O(gate18inter10));
  nor2  gate3008(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate3009(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate3010(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2983(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2984(.a(gate19inter0), .b(s_348), .O(gate19inter1));
  and2  gate2985(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2986(.a(s_348), .O(gate19inter3));
  inv1  gate2987(.a(s_349), .O(gate19inter4));
  nand2 gate2988(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2989(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2990(.a(G21), .O(gate19inter7));
  inv1  gate2991(.a(G22), .O(gate19inter8));
  nand2 gate2992(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2993(.a(s_349), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2994(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2995(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2996(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1625(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1626(.a(gate20inter0), .b(s_154), .O(gate20inter1));
  and2  gate1627(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1628(.a(s_154), .O(gate20inter3));
  inv1  gate1629(.a(s_155), .O(gate20inter4));
  nand2 gate1630(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1631(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1632(.a(G23), .O(gate20inter7));
  inv1  gate1633(.a(G24), .O(gate20inter8));
  nand2 gate1634(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1635(.a(s_155), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1636(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1637(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1638(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate869(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate870(.a(gate21inter0), .b(s_46), .O(gate21inter1));
  and2  gate871(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate872(.a(s_46), .O(gate21inter3));
  inv1  gate873(.a(s_47), .O(gate21inter4));
  nand2 gate874(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate875(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate876(.a(G25), .O(gate21inter7));
  inv1  gate877(.a(G26), .O(gate21inter8));
  nand2 gate878(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate879(.a(s_47), .b(gate21inter3), .O(gate21inter10));
  nor2  gate880(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate881(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate882(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1681(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1682(.a(gate22inter0), .b(s_162), .O(gate22inter1));
  and2  gate1683(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1684(.a(s_162), .O(gate22inter3));
  inv1  gate1685(.a(s_163), .O(gate22inter4));
  nand2 gate1686(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1687(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1688(.a(G27), .O(gate22inter7));
  inv1  gate1689(.a(G28), .O(gate22inter8));
  nand2 gate1690(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1691(.a(s_163), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1692(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1693(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1694(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1149(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1150(.a(gate23inter0), .b(s_86), .O(gate23inter1));
  and2  gate1151(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1152(.a(s_86), .O(gate23inter3));
  inv1  gate1153(.a(s_87), .O(gate23inter4));
  nand2 gate1154(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1155(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1156(.a(G29), .O(gate23inter7));
  inv1  gate1157(.a(G30), .O(gate23inter8));
  nand2 gate1158(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1159(.a(s_87), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1160(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1161(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1162(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1863(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1864(.a(gate27inter0), .b(s_188), .O(gate27inter1));
  and2  gate1865(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1866(.a(s_188), .O(gate27inter3));
  inv1  gate1867(.a(s_189), .O(gate27inter4));
  nand2 gate1868(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1869(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1870(.a(G2), .O(gate27inter7));
  inv1  gate1871(.a(G6), .O(gate27inter8));
  nand2 gate1872(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1873(.a(s_189), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1874(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1875(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1876(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2381(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2382(.a(gate29inter0), .b(s_262), .O(gate29inter1));
  and2  gate2383(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2384(.a(s_262), .O(gate29inter3));
  inv1  gate2385(.a(s_263), .O(gate29inter4));
  nand2 gate2386(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2387(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2388(.a(G3), .O(gate29inter7));
  inv1  gate2389(.a(G7), .O(gate29inter8));
  nand2 gate2390(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2391(.a(s_263), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2392(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2393(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2394(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2241(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2242(.a(gate31inter0), .b(s_242), .O(gate31inter1));
  and2  gate2243(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2244(.a(s_242), .O(gate31inter3));
  inv1  gate2245(.a(s_243), .O(gate31inter4));
  nand2 gate2246(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2247(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2248(.a(G4), .O(gate31inter7));
  inv1  gate2249(.a(G8), .O(gate31inter8));
  nand2 gate2250(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2251(.a(s_243), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2252(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2253(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2254(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1919(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1920(.a(gate32inter0), .b(s_196), .O(gate32inter1));
  and2  gate1921(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1922(.a(s_196), .O(gate32inter3));
  inv1  gate1923(.a(s_197), .O(gate32inter4));
  nand2 gate1924(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1925(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1926(.a(G12), .O(gate32inter7));
  inv1  gate1927(.a(G16), .O(gate32inter8));
  nand2 gate1928(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1929(.a(s_197), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1930(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1931(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1932(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate547(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate548(.a(gate33inter0), .b(s_0), .O(gate33inter1));
  and2  gate549(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate550(.a(s_0), .O(gate33inter3));
  inv1  gate551(.a(s_1), .O(gate33inter4));
  nand2 gate552(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate553(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate554(.a(G17), .O(gate33inter7));
  inv1  gate555(.a(G21), .O(gate33inter8));
  nand2 gate556(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate557(.a(s_1), .b(gate33inter3), .O(gate33inter10));
  nor2  gate558(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate559(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate560(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1261(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1262(.a(gate35inter0), .b(s_102), .O(gate35inter1));
  and2  gate1263(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1264(.a(s_102), .O(gate35inter3));
  inv1  gate1265(.a(s_103), .O(gate35inter4));
  nand2 gate1266(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1267(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1268(.a(G18), .O(gate35inter7));
  inv1  gate1269(.a(G22), .O(gate35inter8));
  nand2 gate1270(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1271(.a(s_103), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1272(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1273(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1274(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2143(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2144(.a(gate36inter0), .b(s_228), .O(gate36inter1));
  and2  gate2145(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2146(.a(s_228), .O(gate36inter3));
  inv1  gate2147(.a(s_229), .O(gate36inter4));
  nand2 gate2148(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2149(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2150(.a(G26), .O(gate36inter7));
  inv1  gate2151(.a(G30), .O(gate36inter8));
  nand2 gate2152(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2153(.a(s_229), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2154(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2155(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2156(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2969(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2970(.a(gate38inter0), .b(s_346), .O(gate38inter1));
  and2  gate2971(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2972(.a(s_346), .O(gate38inter3));
  inv1  gate2973(.a(s_347), .O(gate38inter4));
  nand2 gate2974(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2975(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2976(.a(G27), .O(gate38inter7));
  inv1  gate2977(.a(G31), .O(gate38inter8));
  nand2 gate2978(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2979(.a(s_347), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2980(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2981(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2982(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1135(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1136(.a(gate42inter0), .b(s_84), .O(gate42inter1));
  and2  gate1137(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1138(.a(s_84), .O(gate42inter3));
  inv1  gate1139(.a(s_85), .O(gate42inter4));
  nand2 gate1140(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1141(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1142(.a(G2), .O(gate42inter7));
  inv1  gate1143(.a(G266), .O(gate42inter8));
  nand2 gate1144(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1145(.a(s_85), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1146(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1147(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1148(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2661(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2662(.a(gate48inter0), .b(s_302), .O(gate48inter1));
  and2  gate2663(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2664(.a(s_302), .O(gate48inter3));
  inv1  gate2665(.a(s_303), .O(gate48inter4));
  nand2 gate2666(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2667(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2668(.a(G8), .O(gate48inter7));
  inv1  gate2669(.a(G275), .O(gate48inter8));
  nand2 gate2670(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2671(.a(s_303), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2672(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2673(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2674(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2073(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2074(.a(gate52inter0), .b(s_218), .O(gate52inter1));
  and2  gate2075(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2076(.a(s_218), .O(gate52inter3));
  inv1  gate2077(.a(s_219), .O(gate52inter4));
  nand2 gate2078(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2079(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2080(.a(G12), .O(gate52inter7));
  inv1  gate2081(.a(G281), .O(gate52inter8));
  nand2 gate2082(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2083(.a(s_219), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2084(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2085(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2086(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate2829(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2830(.a(gate53inter0), .b(s_326), .O(gate53inter1));
  and2  gate2831(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2832(.a(s_326), .O(gate53inter3));
  inv1  gate2833(.a(s_327), .O(gate53inter4));
  nand2 gate2834(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2835(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2836(.a(G13), .O(gate53inter7));
  inv1  gate2837(.a(G284), .O(gate53inter8));
  nand2 gate2838(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2839(.a(s_327), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2840(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2841(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2842(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1611(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1612(.a(gate54inter0), .b(s_152), .O(gate54inter1));
  and2  gate1613(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1614(.a(s_152), .O(gate54inter3));
  inv1  gate1615(.a(s_153), .O(gate54inter4));
  nand2 gate1616(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1617(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1618(.a(G14), .O(gate54inter7));
  inv1  gate1619(.a(G284), .O(gate54inter8));
  nand2 gate1620(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1621(.a(s_153), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1622(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1623(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1624(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate2465(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2466(.a(gate55inter0), .b(s_274), .O(gate55inter1));
  and2  gate2467(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2468(.a(s_274), .O(gate55inter3));
  inv1  gate2469(.a(s_275), .O(gate55inter4));
  nand2 gate2470(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2471(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2472(.a(G15), .O(gate55inter7));
  inv1  gate2473(.a(G287), .O(gate55inter8));
  nand2 gate2474(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2475(.a(s_275), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2476(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2477(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2478(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1779(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1780(.a(gate57inter0), .b(s_176), .O(gate57inter1));
  and2  gate1781(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1782(.a(s_176), .O(gate57inter3));
  inv1  gate1783(.a(s_177), .O(gate57inter4));
  nand2 gate1784(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1785(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1786(.a(G17), .O(gate57inter7));
  inv1  gate1787(.a(G290), .O(gate57inter8));
  nand2 gate1788(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1789(.a(s_177), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1790(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1791(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1792(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate3011(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate3012(.a(gate61inter0), .b(s_352), .O(gate61inter1));
  and2  gate3013(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate3014(.a(s_352), .O(gate61inter3));
  inv1  gate3015(.a(s_353), .O(gate61inter4));
  nand2 gate3016(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate3017(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate3018(.a(G21), .O(gate61inter7));
  inv1  gate3019(.a(G296), .O(gate61inter8));
  nand2 gate3020(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate3021(.a(s_353), .b(gate61inter3), .O(gate61inter10));
  nor2  gate3022(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate3023(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate3024(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2493(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2494(.a(gate64inter0), .b(s_278), .O(gate64inter1));
  and2  gate2495(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2496(.a(s_278), .O(gate64inter3));
  inv1  gate2497(.a(s_279), .O(gate64inter4));
  nand2 gate2498(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2499(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2500(.a(G24), .O(gate64inter7));
  inv1  gate2501(.a(G299), .O(gate64inter8));
  nand2 gate2502(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2503(.a(s_279), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2504(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2505(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2506(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate785(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate786(.a(gate65inter0), .b(s_34), .O(gate65inter1));
  and2  gate787(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate788(.a(s_34), .O(gate65inter3));
  inv1  gate789(.a(s_35), .O(gate65inter4));
  nand2 gate790(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate791(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate792(.a(G25), .O(gate65inter7));
  inv1  gate793(.a(G302), .O(gate65inter8));
  nand2 gate794(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate795(.a(s_35), .b(gate65inter3), .O(gate65inter10));
  nor2  gate796(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate797(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate798(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate967(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate968(.a(gate66inter0), .b(s_60), .O(gate66inter1));
  and2  gate969(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate970(.a(s_60), .O(gate66inter3));
  inv1  gate971(.a(s_61), .O(gate66inter4));
  nand2 gate972(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate973(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate974(.a(G26), .O(gate66inter7));
  inv1  gate975(.a(G302), .O(gate66inter8));
  nand2 gate976(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate977(.a(s_61), .b(gate66inter3), .O(gate66inter10));
  nor2  gate978(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate979(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate980(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2045(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2046(.a(gate68inter0), .b(s_214), .O(gate68inter1));
  and2  gate2047(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2048(.a(s_214), .O(gate68inter3));
  inv1  gate2049(.a(s_215), .O(gate68inter4));
  nand2 gate2050(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2051(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2052(.a(G28), .O(gate68inter7));
  inv1  gate2053(.a(G305), .O(gate68inter8));
  nand2 gate2054(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2055(.a(s_215), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2056(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2057(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2058(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2577(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2578(.a(gate70inter0), .b(s_290), .O(gate70inter1));
  and2  gate2579(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2580(.a(s_290), .O(gate70inter3));
  inv1  gate2581(.a(s_291), .O(gate70inter4));
  nand2 gate2582(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2583(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2584(.a(G30), .O(gate70inter7));
  inv1  gate2585(.a(G308), .O(gate70inter8));
  nand2 gate2586(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2587(.a(s_291), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2588(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2589(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2590(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1667(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1668(.a(gate71inter0), .b(s_160), .O(gate71inter1));
  and2  gate1669(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1670(.a(s_160), .O(gate71inter3));
  inv1  gate1671(.a(s_161), .O(gate71inter4));
  nand2 gate1672(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1673(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1674(.a(G31), .O(gate71inter7));
  inv1  gate1675(.a(G311), .O(gate71inter8));
  nand2 gate1676(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1677(.a(s_161), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1678(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1679(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1680(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate3109(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate3110(.a(gate72inter0), .b(s_366), .O(gate72inter1));
  and2  gate3111(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate3112(.a(s_366), .O(gate72inter3));
  inv1  gate3113(.a(s_367), .O(gate72inter4));
  nand2 gate3114(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate3115(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate3116(.a(G32), .O(gate72inter7));
  inv1  gate3117(.a(G311), .O(gate72inter8));
  nand2 gate3118(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate3119(.a(s_367), .b(gate72inter3), .O(gate72inter10));
  nor2  gate3120(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate3121(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate3122(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate2423(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2424(.a(gate73inter0), .b(s_268), .O(gate73inter1));
  and2  gate2425(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2426(.a(s_268), .O(gate73inter3));
  inv1  gate2427(.a(s_269), .O(gate73inter4));
  nand2 gate2428(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2429(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2430(.a(G1), .O(gate73inter7));
  inv1  gate2431(.a(G314), .O(gate73inter8));
  nand2 gate2432(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2433(.a(s_269), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2434(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2435(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2436(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2605(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2606(.a(gate74inter0), .b(s_294), .O(gate74inter1));
  and2  gate2607(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2608(.a(s_294), .O(gate74inter3));
  inv1  gate2609(.a(s_295), .O(gate74inter4));
  nand2 gate2610(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2611(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2612(.a(G5), .O(gate74inter7));
  inv1  gate2613(.a(G314), .O(gate74inter8));
  nand2 gate2614(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2615(.a(s_295), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2616(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2617(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2618(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1849(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1850(.a(gate76inter0), .b(s_186), .O(gate76inter1));
  and2  gate1851(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1852(.a(s_186), .O(gate76inter3));
  inv1  gate1853(.a(s_187), .O(gate76inter4));
  nand2 gate1854(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1855(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1856(.a(G13), .O(gate76inter7));
  inv1  gate1857(.a(G317), .O(gate76inter8));
  nand2 gate1858(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1859(.a(s_187), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1860(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1861(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1862(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate659(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate660(.a(gate77inter0), .b(s_16), .O(gate77inter1));
  and2  gate661(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate662(.a(s_16), .O(gate77inter3));
  inv1  gate663(.a(s_17), .O(gate77inter4));
  nand2 gate664(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate665(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate666(.a(G2), .O(gate77inter7));
  inv1  gate667(.a(G320), .O(gate77inter8));
  nand2 gate668(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate669(.a(s_17), .b(gate77inter3), .O(gate77inter10));
  nor2  gate670(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate671(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate672(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1205(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1206(.a(gate78inter0), .b(s_94), .O(gate78inter1));
  and2  gate1207(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1208(.a(s_94), .O(gate78inter3));
  inv1  gate1209(.a(s_95), .O(gate78inter4));
  nand2 gate1210(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1211(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1212(.a(G6), .O(gate78inter7));
  inv1  gate1213(.a(G320), .O(gate78inter8));
  nand2 gate1214(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1215(.a(s_95), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1216(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1217(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1218(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1009(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1010(.a(gate82inter0), .b(s_66), .O(gate82inter1));
  and2  gate1011(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1012(.a(s_66), .O(gate82inter3));
  inv1  gate1013(.a(s_67), .O(gate82inter4));
  nand2 gate1014(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1015(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1016(.a(G7), .O(gate82inter7));
  inv1  gate1017(.a(G326), .O(gate82inter8));
  nand2 gate1018(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1019(.a(s_67), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1020(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1021(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1022(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2633(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2634(.a(gate84inter0), .b(s_298), .O(gate84inter1));
  and2  gate2635(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2636(.a(s_298), .O(gate84inter3));
  inv1  gate2637(.a(s_299), .O(gate84inter4));
  nand2 gate2638(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2639(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2640(.a(G15), .O(gate84inter7));
  inv1  gate2641(.a(G329), .O(gate84inter8));
  nand2 gate2642(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2643(.a(s_299), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2644(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2645(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2646(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1541(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1542(.a(gate85inter0), .b(s_142), .O(gate85inter1));
  and2  gate1543(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1544(.a(s_142), .O(gate85inter3));
  inv1  gate1545(.a(s_143), .O(gate85inter4));
  nand2 gate1546(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1547(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1548(.a(G4), .O(gate85inter7));
  inv1  gate1549(.a(G332), .O(gate85inter8));
  nand2 gate1550(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1551(.a(s_143), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1552(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1553(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1554(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1191(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1192(.a(gate86inter0), .b(s_92), .O(gate86inter1));
  and2  gate1193(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1194(.a(s_92), .O(gate86inter3));
  inv1  gate1195(.a(s_93), .O(gate86inter4));
  nand2 gate1196(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1197(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1198(.a(G8), .O(gate86inter7));
  inv1  gate1199(.a(G332), .O(gate86inter8));
  nand2 gate1200(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1201(.a(s_93), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1202(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1203(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1204(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate883(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate884(.a(gate87inter0), .b(s_48), .O(gate87inter1));
  and2  gate885(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate886(.a(s_48), .O(gate87inter3));
  inv1  gate887(.a(s_49), .O(gate87inter4));
  nand2 gate888(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate889(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate890(.a(G12), .O(gate87inter7));
  inv1  gate891(.a(G335), .O(gate87inter8));
  nand2 gate892(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate893(.a(s_49), .b(gate87inter3), .O(gate87inter10));
  nor2  gate894(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate895(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate896(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate2927(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2928(.a(gate88inter0), .b(s_340), .O(gate88inter1));
  and2  gate2929(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2930(.a(s_340), .O(gate88inter3));
  inv1  gate2931(.a(s_341), .O(gate88inter4));
  nand2 gate2932(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2933(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2934(.a(G16), .O(gate88inter7));
  inv1  gate2935(.a(G335), .O(gate88inter8));
  nand2 gate2936(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2937(.a(s_341), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2938(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2939(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2940(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate841(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate842(.a(gate89inter0), .b(s_42), .O(gate89inter1));
  and2  gate843(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate844(.a(s_42), .O(gate89inter3));
  inv1  gate845(.a(s_43), .O(gate89inter4));
  nand2 gate846(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate847(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate848(.a(G17), .O(gate89inter7));
  inv1  gate849(.a(G338), .O(gate89inter8));
  nand2 gate850(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate851(.a(s_43), .b(gate89inter3), .O(gate89inter10));
  nor2  gate852(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate853(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate854(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1331(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1332(.a(gate90inter0), .b(s_112), .O(gate90inter1));
  and2  gate1333(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1334(.a(s_112), .O(gate90inter3));
  inv1  gate1335(.a(s_113), .O(gate90inter4));
  nand2 gate1336(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1337(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1338(.a(G21), .O(gate90inter7));
  inv1  gate1339(.a(G338), .O(gate90inter8));
  nand2 gate1340(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1341(.a(s_113), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1342(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1343(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1344(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2731(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2732(.a(gate94inter0), .b(s_312), .O(gate94inter1));
  and2  gate2733(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2734(.a(s_312), .O(gate94inter3));
  inv1  gate2735(.a(s_313), .O(gate94inter4));
  nand2 gate2736(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2737(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2738(.a(G22), .O(gate94inter7));
  inv1  gate2739(.a(G344), .O(gate94inter8));
  nand2 gate2740(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2741(.a(s_313), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2742(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2743(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2744(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate2647(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2648(.a(gate95inter0), .b(s_300), .O(gate95inter1));
  and2  gate2649(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2650(.a(s_300), .O(gate95inter3));
  inv1  gate2651(.a(s_301), .O(gate95inter4));
  nand2 gate2652(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2653(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2654(.a(G26), .O(gate95inter7));
  inv1  gate2655(.a(G347), .O(gate95inter8));
  nand2 gate2656(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2657(.a(s_301), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2658(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2659(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2660(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate687(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate688(.a(gate97inter0), .b(s_20), .O(gate97inter1));
  and2  gate689(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate690(.a(s_20), .O(gate97inter3));
  inv1  gate691(.a(s_21), .O(gate97inter4));
  nand2 gate692(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate693(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate694(.a(G19), .O(gate97inter7));
  inv1  gate695(.a(G350), .O(gate97inter8));
  nand2 gate696(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate697(.a(s_21), .b(gate97inter3), .O(gate97inter10));
  nor2  gate698(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate699(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate700(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate2227(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2228(.a(gate103inter0), .b(s_240), .O(gate103inter1));
  and2  gate2229(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2230(.a(s_240), .O(gate103inter3));
  inv1  gate2231(.a(s_241), .O(gate103inter4));
  nand2 gate2232(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2233(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2234(.a(G28), .O(gate103inter7));
  inv1  gate2235(.a(G359), .O(gate103inter8));
  nand2 gate2236(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2237(.a(s_241), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2238(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2239(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2240(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2395(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2396(.a(gate104inter0), .b(s_264), .O(gate104inter1));
  and2  gate2397(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2398(.a(s_264), .O(gate104inter3));
  inv1  gate2399(.a(s_265), .O(gate104inter4));
  nand2 gate2400(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2401(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2402(.a(G32), .O(gate104inter7));
  inv1  gate2403(.a(G359), .O(gate104inter8));
  nand2 gate2404(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2405(.a(s_265), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2406(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2407(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2408(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2129(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2130(.a(gate107inter0), .b(s_226), .O(gate107inter1));
  and2  gate2131(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2132(.a(s_226), .O(gate107inter3));
  inv1  gate2133(.a(s_227), .O(gate107inter4));
  nand2 gate2134(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2135(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2136(.a(G366), .O(gate107inter7));
  inv1  gate2137(.a(G367), .O(gate107inter8));
  nand2 gate2138(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2139(.a(s_227), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2140(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2141(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2142(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate743(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate744(.a(gate111inter0), .b(s_28), .O(gate111inter1));
  and2  gate745(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate746(.a(s_28), .O(gate111inter3));
  inv1  gate747(.a(s_29), .O(gate111inter4));
  nand2 gate748(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate749(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate750(.a(G374), .O(gate111inter7));
  inv1  gate751(.a(G375), .O(gate111inter8));
  nand2 gate752(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate753(.a(s_29), .b(gate111inter3), .O(gate111inter10));
  nor2  gate754(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate755(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate756(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate799(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate800(.a(gate114inter0), .b(s_36), .O(gate114inter1));
  and2  gate801(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate802(.a(s_36), .O(gate114inter3));
  inv1  gate803(.a(s_37), .O(gate114inter4));
  nand2 gate804(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate805(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate806(.a(G380), .O(gate114inter7));
  inv1  gate807(.a(G381), .O(gate114inter8));
  nand2 gate808(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate809(.a(s_37), .b(gate114inter3), .O(gate114inter10));
  nor2  gate810(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate811(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate812(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2101(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2102(.a(gate118inter0), .b(s_222), .O(gate118inter1));
  and2  gate2103(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2104(.a(s_222), .O(gate118inter3));
  inv1  gate2105(.a(s_223), .O(gate118inter4));
  nand2 gate2106(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2107(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2108(.a(G388), .O(gate118inter7));
  inv1  gate2109(.a(G389), .O(gate118inter8));
  nand2 gate2110(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2111(.a(s_223), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2112(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2113(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2114(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1079(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1080(.a(gate122inter0), .b(s_76), .O(gate122inter1));
  and2  gate1081(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1082(.a(s_76), .O(gate122inter3));
  inv1  gate1083(.a(s_77), .O(gate122inter4));
  nand2 gate1084(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1085(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1086(.a(G396), .O(gate122inter7));
  inv1  gate1087(.a(G397), .O(gate122inter8));
  nand2 gate1088(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1089(.a(s_77), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1090(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1091(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1092(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate813(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate814(.a(gate123inter0), .b(s_38), .O(gate123inter1));
  and2  gate815(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate816(.a(s_38), .O(gate123inter3));
  inv1  gate817(.a(s_39), .O(gate123inter4));
  nand2 gate818(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate819(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate820(.a(G398), .O(gate123inter7));
  inv1  gate821(.a(G399), .O(gate123inter8));
  nand2 gate822(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate823(.a(s_39), .b(gate123inter3), .O(gate123inter10));
  nor2  gate824(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate825(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate826(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2703(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2704(.a(gate125inter0), .b(s_308), .O(gate125inter1));
  and2  gate2705(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2706(.a(s_308), .O(gate125inter3));
  inv1  gate2707(.a(s_309), .O(gate125inter4));
  nand2 gate2708(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2709(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2710(.a(G402), .O(gate125inter7));
  inv1  gate2711(.a(G403), .O(gate125inter8));
  nand2 gate2712(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2713(.a(s_309), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2714(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2715(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2716(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2115(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2116(.a(gate128inter0), .b(s_224), .O(gate128inter1));
  and2  gate2117(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2118(.a(s_224), .O(gate128inter3));
  inv1  gate2119(.a(s_225), .O(gate128inter4));
  nand2 gate2120(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2121(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2122(.a(G408), .O(gate128inter7));
  inv1  gate2123(.a(G409), .O(gate128inter8));
  nand2 gate2124(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2125(.a(s_225), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2126(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2127(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2128(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1275(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1276(.a(gate132inter0), .b(s_104), .O(gate132inter1));
  and2  gate1277(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1278(.a(s_104), .O(gate132inter3));
  inv1  gate1279(.a(s_105), .O(gate132inter4));
  nand2 gate1280(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1281(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1282(.a(G416), .O(gate132inter7));
  inv1  gate1283(.a(G417), .O(gate132inter8));
  nand2 gate1284(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1285(.a(s_105), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1286(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1287(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1288(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2913(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2914(.a(gate134inter0), .b(s_338), .O(gate134inter1));
  and2  gate2915(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2916(.a(s_338), .O(gate134inter3));
  inv1  gate2917(.a(s_339), .O(gate134inter4));
  nand2 gate2918(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2919(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2920(.a(G420), .O(gate134inter7));
  inv1  gate2921(.a(G421), .O(gate134inter8));
  nand2 gate2922(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2923(.a(s_339), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2924(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2925(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2926(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate1793(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1794(.a(gate135inter0), .b(s_178), .O(gate135inter1));
  and2  gate1795(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1796(.a(s_178), .O(gate135inter3));
  inv1  gate1797(.a(s_179), .O(gate135inter4));
  nand2 gate1798(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1799(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1800(.a(G422), .O(gate135inter7));
  inv1  gate1801(.a(G423), .O(gate135inter8));
  nand2 gate1802(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1803(.a(s_179), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1804(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1805(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1806(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1527(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1528(.a(gate136inter0), .b(s_140), .O(gate136inter1));
  and2  gate1529(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1530(.a(s_140), .O(gate136inter3));
  inv1  gate1531(.a(s_141), .O(gate136inter4));
  nand2 gate1532(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1533(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1534(.a(G424), .O(gate136inter7));
  inv1  gate1535(.a(G425), .O(gate136inter8));
  nand2 gate1536(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1537(.a(s_141), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1538(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1539(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1540(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2857(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2858(.a(gate139inter0), .b(s_330), .O(gate139inter1));
  and2  gate2859(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2860(.a(s_330), .O(gate139inter3));
  inv1  gate2861(.a(s_331), .O(gate139inter4));
  nand2 gate2862(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2863(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2864(.a(G438), .O(gate139inter7));
  inv1  gate2865(.a(G441), .O(gate139inter8));
  nand2 gate2866(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2867(.a(s_331), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2868(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2869(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2870(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1597(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1598(.a(gate142inter0), .b(s_150), .O(gate142inter1));
  and2  gate1599(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1600(.a(s_150), .O(gate142inter3));
  inv1  gate1601(.a(s_151), .O(gate142inter4));
  nand2 gate1602(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1603(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1604(.a(G456), .O(gate142inter7));
  inv1  gate1605(.a(G459), .O(gate142inter8));
  nand2 gate1606(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1607(.a(s_151), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1608(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1609(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1610(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1093(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1094(.a(gate144inter0), .b(s_78), .O(gate144inter1));
  and2  gate1095(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1096(.a(s_78), .O(gate144inter3));
  inv1  gate1097(.a(s_79), .O(gate144inter4));
  nand2 gate1098(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1099(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1100(.a(G468), .O(gate144inter7));
  inv1  gate1101(.a(G471), .O(gate144inter8));
  nand2 gate1102(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1103(.a(s_79), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1104(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1105(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1106(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate3039(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate3040(.a(gate145inter0), .b(s_356), .O(gate145inter1));
  and2  gate3041(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate3042(.a(s_356), .O(gate145inter3));
  inv1  gate3043(.a(s_357), .O(gate145inter4));
  nand2 gate3044(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate3045(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate3046(.a(G474), .O(gate145inter7));
  inv1  gate3047(.a(G477), .O(gate145inter8));
  nand2 gate3048(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate3049(.a(s_357), .b(gate145inter3), .O(gate145inter10));
  nor2  gate3050(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate3051(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate3052(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2759(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2760(.a(gate148inter0), .b(s_316), .O(gate148inter1));
  and2  gate2761(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2762(.a(s_316), .O(gate148inter3));
  inv1  gate2763(.a(s_317), .O(gate148inter4));
  nand2 gate2764(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2765(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2766(.a(G492), .O(gate148inter7));
  inv1  gate2767(.a(G495), .O(gate148inter8));
  nand2 gate2768(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2769(.a(s_317), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2770(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2771(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2772(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2787(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2788(.a(gate150inter0), .b(s_320), .O(gate150inter1));
  and2  gate2789(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2790(.a(s_320), .O(gate150inter3));
  inv1  gate2791(.a(s_321), .O(gate150inter4));
  nand2 gate2792(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2793(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2794(.a(G504), .O(gate150inter7));
  inv1  gate2795(.a(G507), .O(gate150inter8));
  nand2 gate2796(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2797(.a(s_321), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2798(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2799(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2800(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2941(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2942(.a(gate152inter0), .b(s_342), .O(gate152inter1));
  and2  gate2943(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2944(.a(s_342), .O(gate152inter3));
  inv1  gate2945(.a(s_343), .O(gate152inter4));
  nand2 gate2946(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2947(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2948(.a(G516), .O(gate152inter7));
  inv1  gate2949(.a(G519), .O(gate152inter8));
  nand2 gate2950(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2951(.a(s_343), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2952(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2953(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2954(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate855(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate856(.a(gate156inter0), .b(s_44), .O(gate156inter1));
  and2  gate857(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate858(.a(s_44), .O(gate156inter3));
  inv1  gate859(.a(s_45), .O(gate156inter4));
  nand2 gate860(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate861(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate862(.a(G435), .O(gate156inter7));
  inv1  gate863(.a(G525), .O(gate156inter8));
  nand2 gate864(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate865(.a(s_45), .b(gate156inter3), .O(gate156inter10));
  nor2  gate866(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate867(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate868(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1345(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1346(.a(gate159inter0), .b(s_114), .O(gate159inter1));
  and2  gate1347(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1348(.a(s_114), .O(gate159inter3));
  inv1  gate1349(.a(s_115), .O(gate159inter4));
  nand2 gate1350(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1351(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1352(.a(G444), .O(gate159inter7));
  inv1  gate1353(.a(G531), .O(gate159inter8));
  nand2 gate1354(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1355(.a(s_115), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1356(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1357(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1358(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1961(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1962(.a(gate160inter0), .b(s_202), .O(gate160inter1));
  and2  gate1963(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1964(.a(s_202), .O(gate160inter3));
  inv1  gate1965(.a(s_203), .O(gate160inter4));
  nand2 gate1966(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1967(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1968(.a(G447), .O(gate160inter7));
  inv1  gate1969(.a(G531), .O(gate160inter8));
  nand2 gate1970(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1971(.a(s_203), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1972(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1973(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1974(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1933(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1934(.a(gate165inter0), .b(s_198), .O(gate165inter1));
  and2  gate1935(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1936(.a(s_198), .O(gate165inter3));
  inv1  gate1937(.a(s_199), .O(gate165inter4));
  nand2 gate1938(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1939(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1940(.a(G462), .O(gate165inter7));
  inv1  gate1941(.a(G540), .O(gate165inter8));
  nand2 gate1942(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1943(.a(s_199), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1944(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1945(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1946(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate2185(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2186(.a(gate166inter0), .b(s_234), .O(gate166inter1));
  and2  gate2187(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2188(.a(s_234), .O(gate166inter3));
  inv1  gate2189(.a(s_235), .O(gate166inter4));
  nand2 gate2190(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2191(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2192(.a(G465), .O(gate166inter7));
  inv1  gate2193(.a(G540), .O(gate166inter8));
  nand2 gate2194(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2195(.a(s_235), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2196(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2197(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2198(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1289(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1290(.a(gate172inter0), .b(s_106), .O(gate172inter1));
  and2  gate1291(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1292(.a(s_106), .O(gate172inter3));
  inv1  gate1293(.a(s_107), .O(gate172inter4));
  nand2 gate1294(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1295(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1296(.a(G483), .O(gate172inter7));
  inv1  gate1297(.a(G549), .O(gate172inter8));
  nand2 gate1298(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1299(.a(s_107), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1300(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1301(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1302(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2325(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2326(.a(gate173inter0), .b(s_254), .O(gate173inter1));
  and2  gate2327(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2328(.a(s_254), .O(gate173inter3));
  inv1  gate2329(.a(s_255), .O(gate173inter4));
  nand2 gate2330(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2331(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2332(.a(G486), .O(gate173inter7));
  inv1  gate2333(.a(G552), .O(gate173inter8));
  nand2 gate2334(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2335(.a(s_255), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2336(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2337(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2338(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1303(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1304(.a(gate176inter0), .b(s_108), .O(gate176inter1));
  and2  gate1305(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1306(.a(s_108), .O(gate176inter3));
  inv1  gate1307(.a(s_109), .O(gate176inter4));
  nand2 gate1308(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1309(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1310(.a(G495), .O(gate176inter7));
  inv1  gate1311(.a(G555), .O(gate176inter8));
  nand2 gate1312(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1313(.a(s_109), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1314(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1315(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1316(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate897(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate898(.a(gate177inter0), .b(s_50), .O(gate177inter1));
  and2  gate899(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate900(.a(s_50), .O(gate177inter3));
  inv1  gate901(.a(s_51), .O(gate177inter4));
  nand2 gate902(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate903(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate904(.a(G498), .O(gate177inter7));
  inv1  gate905(.a(G558), .O(gate177inter8));
  nand2 gate906(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate907(.a(s_51), .b(gate177inter3), .O(gate177inter10));
  nor2  gate908(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate909(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate910(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1121(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1122(.a(gate180inter0), .b(s_82), .O(gate180inter1));
  and2  gate1123(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1124(.a(s_82), .O(gate180inter3));
  inv1  gate1125(.a(s_83), .O(gate180inter4));
  nand2 gate1126(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1127(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1128(.a(G507), .O(gate180inter7));
  inv1  gate1129(.a(G561), .O(gate180inter8));
  nand2 gate1130(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1131(.a(s_83), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1132(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1133(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1134(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1233(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1234(.a(gate181inter0), .b(s_98), .O(gate181inter1));
  and2  gate1235(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1236(.a(s_98), .O(gate181inter3));
  inv1  gate1237(.a(s_99), .O(gate181inter4));
  nand2 gate1238(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1239(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1240(.a(G510), .O(gate181inter7));
  inv1  gate1241(.a(G564), .O(gate181inter8));
  nand2 gate1242(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1243(.a(s_99), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1244(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1245(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1246(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1401(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1402(.a(gate182inter0), .b(s_122), .O(gate182inter1));
  and2  gate1403(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1404(.a(s_122), .O(gate182inter3));
  inv1  gate1405(.a(s_123), .O(gate182inter4));
  nand2 gate1406(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1407(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1408(.a(G513), .O(gate182inter7));
  inv1  gate1409(.a(G564), .O(gate182inter8));
  nand2 gate1410(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1411(.a(s_123), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1412(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1413(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1414(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1485(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1486(.a(gate183inter0), .b(s_134), .O(gate183inter1));
  and2  gate1487(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1488(.a(s_134), .O(gate183inter3));
  inv1  gate1489(.a(s_135), .O(gate183inter4));
  nand2 gate1490(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1491(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1492(.a(G516), .O(gate183inter7));
  inv1  gate1493(.a(G567), .O(gate183inter8));
  nand2 gate1494(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1495(.a(s_135), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1496(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1497(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1498(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate911(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate912(.a(gate184inter0), .b(s_52), .O(gate184inter1));
  and2  gate913(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate914(.a(s_52), .O(gate184inter3));
  inv1  gate915(.a(s_53), .O(gate184inter4));
  nand2 gate916(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate917(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate918(.a(G519), .O(gate184inter7));
  inv1  gate919(.a(G567), .O(gate184inter8));
  nand2 gate920(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate921(.a(s_53), .b(gate184inter3), .O(gate184inter10));
  nor2  gate922(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate923(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate924(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1807(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1808(.a(gate185inter0), .b(s_180), .O(gate185inter1));
  and2  gate1809(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1810(.a(s_180), .O(gate185inter3));
  inv1  gate1811(.a(s_181), .O(gate185inter4));
  nand2 gate1812(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1813(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1814(.a(G570), .O(gate185inter7));
  inv1  gate1815(.a(G571), .O(gate185inter8));
  nand2 gate1816(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1817(.a(s_181), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1818(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1819(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1820(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate589(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate590(.a(gate186inter0), .b(s_6), .O(gate186inter1));
  and2  gate591(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate592(.a(s_6), .O(gate186inter3));
  inv1  gate593(.a(s_7), .O(gate186inter4));
  nand2 gate594(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate595(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate596(.a(G572), .O(gate186inter7));
  inv1  gate597(.a(G573), .O(gate186inter8));
  nand2 gate598(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate599(.a(s_7), .b(gate186inter3), .O(gate186inter10));
  nor2  gate600(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate601(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate602(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1051(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1052(.a(gate188inter0), .b(s_72), .O(gate188inter1));
  and2  gate1053(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1054(.a(s_72), .O(gate188inter3));
  inv1  gate1055(.a(s_73), .O(gate188inter4));
  nand2 gate1056(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1057(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1058(.a(G576), .O(gate188inter7));
  inv1  gate1059(.a(G577), .O(gate188inter8));
  nand2 gate1060(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1061(.a(s_73), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1062(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1063(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1064(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1989(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1990(.a(gate190inter0), .b(s_206), .O(gate190inter1));
  and2  gate1991(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1992(.a(s_206), .O(gate190inter3));
  inv1  gate1993(.a(s_207), .O(gate190inter4));
  nand2 gate1994(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1995(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1996(.a(G580), .O(gate190inter7));
  inv1  gate1997(.a(G581), .O(gate190inter8));
  nand2 gate1998(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1999(.a(s_207), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2000(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2001(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2002(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2255(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2256(.a(gate192inter0), .b(s_244), .O(gate192inter1));
  and2  gate2257(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2258(.a(s_244), .O(gate192inter3));
  inv1  gate2259(.a(s_245), .O(gate192inter4));
  nand2 gate2260(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2261(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2262(.a(G584), .O(gate192inter7));
  inv1  gate2263(.a(G585), .O(gate192inter8));
  nand2 gate2264(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2265(.a(s_245), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2266(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2267(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2268(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1457(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1458(.a(gate194inter0), .b(s_130), .O(gate194inter1));
  and2  gate1459(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1460(.a(s_130), .O(gate194inter3));
  inv1  gate1461(.a(s_131), .O(gate194inter4));
  nand2 gate1462(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1463(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1464(.a(G588), .O(gate194inter7));
  inv1  gate1465(.a(G589), .O(gate194inter8));
  nand2 gate1466(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1467(.a(s_131), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1468(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1469(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1470(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate3025(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate3026(.a(gate195inter0), .b(s_354), .O(gate195inter1));
  and2  gate3027(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate3028(.a(s_354), .O(gate195inter3));
  inv1  gate3029(.a(s_355), .O(gate195inter4));
  nand2 gate3030(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate3031(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate3032(.a(G590), .O(gate195inter7));
  inv1  gate3033(.a(G591), .O(gate195inter8));
  nand2 gate3034(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate3035(.a(s_355), .b(gate195inter3), .O(gate195inter10));
  nor2  gate3036(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate3037(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate3038(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1247(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1248(.a(gate199inter0), .b(s_100), .O(gate199inter1));
  and2  gate1249(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1250(.a(s_100), .O(gate199inter3));
  inv1  gate1251(.a(s_101), .O(gate199inter4));
  nand2 gate1252(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1253(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1254(.a(G598), .O(gate199inter7));
  inv1  gate1255(.a(G599), .O(gate199inter8));
  nand2 gate1256(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1257(.a(s_101), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1258(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1259(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1260(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate2717(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2718(.a(gate200inter0), .b(s_310), .O(gate200inter1));
  and2  gate2719(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2720(.a(s_310), .O(gate200inter3));
  inv1  gate2721(.a(s_311), .O(gate200inter4));
  nand2 gate2722(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2723(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2724(.a(G600), .O(gate200inter7));
  inv1  gate2725(.a(G601), .O(gate200inter8));
  nand2 gate2726(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2727(.a(s_311), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2728(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2729(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2730(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate771(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate772(.a(gate202inter0), .b(s_32), .O(gate202inter1));
  and2  gate773(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate774(.a(s_32), .O(gate202inter3));
  inv1  gate775(.a(s_33), .O(gate202inter4));
  nand2 gate776(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate777(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate778(.a(G612), .O(gate202inter7));
  inv1  gate779(.a(G617), .O(gate202inter8));
  nand2 gate780(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate781(.a(s_33), .b(gate202inter3), .O(gate202inter10));
  nor2  gate782(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate783(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate784(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1821(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1822(.a(gate204inter0), .b(s_182), .O(gate204inter1));
  and2  gate1823(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1824(.a(s_182), .O(gate204inter3));
  inv1  gate1825(.a(s_183), .O(gate204inter4));
  nand2 gate1826(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1827(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1828(.a(G607), .O(gate204inter7));
  inv1  gate1829(.a(G617), .O(gate204inter8));
  nand2 gate1830(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1831(.a(s_183), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1832(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1833(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1834(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2801(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2802(.a(gate206inter0), .b(s_322), .O(gate206inter1));
  and2  gate2803(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2804(.a(s_322), .O(gate206inter3));
  inv1  gate2805(.a(s_323), .O(gate206inter4));
  nand2 gate2806(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2807(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2808(.a(G632), .O(gate206inter7));
  inv1  gate2809(.a(G637), .O(gate206inter8));
  nand2 gate2810(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2811(.a(s_323), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2812(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2813(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2814(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2745(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2746(.a(gate211inter0), .b(s_314), .O(gate211inter1));
  and2  gate2747(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2748(.a(s_314), .O(gate211inter3));
  inv1  gate2749(.a(s_315), .O(gate211inter4));
  nand2 gate2750(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2751(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2752(.a(G612), .O(gate211inter7));
  inv1  gate2753(.a(G669), .O(gate211inter8));
  nand2 gate2754(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2755(.a(s_315), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2756(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2757(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2758(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate925(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate926(.a(gate217inter0), .b(s_54), .O(gate217inter1));
  and2  gate927(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate928(.a(s_54), .O(gate217inter3));
  inv1  gate929(.a(s_55), .O(gate217inter4));
  nand2 gate930(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate931(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate932(.a(G622), .O(gate217inter7));
  inv1  gate933(.a(G678), .O(gate217inter8));
  nand2 gate934(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate935(.a(s_55), .b(gate217inter3), .O(gate217inter10));
  nor2  gate936(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate937(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate938(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1443(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1444(.a(gate226inter0), .b(s_128), .O(gate226inter1));
  and2  gate1445(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1446(.a(s_128), .O(gate226inter3));
  inv1  gate1447(.a(s_129), .O(gate226inter4));
  nand2 gate1448(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1449(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1450(.a(G692), .O(gate226inter7));
  inv1  gate1451(.a(G693), .O(gate226inter8));
  nand2 gate1452(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1453(.a(s_129), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1454(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1455(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1456(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1065(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1066(.a(gate228inter0), .b(s_74), .O(gate228inter1));
  and2  gate1067(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1068(.a(s_74), .O(gate228inter3));
  inv1  gate1069(.a(s_75), .O(gate228inter4));
  nand2 gate1070(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1071(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1072(.a(G696), .O(gate228inter7));
  inv1  gate1073(.a(G697), .O(gate228inter8));
  nand2 gate1074(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1075(.a(s_75), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1076(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1077(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1078(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1415(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1416(.a(gate230inter0), .b(s_124), .O(gate230inter1));
  and2  gate1417(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1418(.a(s_124), .O(gate230inter3));
  inv1  gate1419(.a(s_125), .O(gate230inter4));
  nand2 gate1420(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1421(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1422(.a(G700), .O(gate230inter7));
  inv1  gate1423(.a(G701), .O(gate230inter8));
  nand2 gate1424(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1425(.a(s_125), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1426(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1427(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1428(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2353(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2354(.a(gate233inter0), .b(s_258), .O(gate233inter1));
  and2  gate2355(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2356(.a(s_258), .O(gate233inter3));
  inv1  gate2357(.a(s_259), .O(gate233inter4));
  nand2 gate2358(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2359(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2360(.a(G242), .O(gate233inter7));
  inv1  gate2361(.a(G718), .O(gate233inter8));
  nand2 gate2362(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2363(.a(s_259), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2364(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2365(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2366(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2563(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2564(.a(gate236inter0), .b(s_288), .O(gate236inter1));
  and2  gate2565(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2566(.a(s_288), .O(gate236inter3));
  inv1  gate2567(.a(s_289), .O(gate236inter4));
  nand2 gate2568(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2569(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2570(.a(G251), .O(gate236inter7));
  inv1  gate2571(.a(G727), .O(gate236inter8));
  nand2 gate2572(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2573(.a(s_289), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2574(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2575(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2576(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2815(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2816(.a(gate240inter0), .b(s_324), .O(gate240inter1));
  and2  gate2817(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2818(.a(s_324), .O(gate240inter3));
  inv1  gate2819(.a(s_325), .O(gate240inter4));
  nand2 gate2820(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2821(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2822(.a(G263), .O(gate240inter7));
  inv1  gate2823(.a(G715), .O(gate240inter8));
  nand2 gate2824(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2825(.a(s_325), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2826(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2827(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2828(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2871(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2872(.a(gate242inter0), .b(s_332), .O(gate242inter1));
  and2  gate2873(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2874(.a(s_332), .O(gate242inter3));
  inv1  gate2875(.a(s_333), .O(gate242inter4));
  nand2 gate2876(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2877(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2878(.a(G718), .O(gate242inter7));
  inv1  gate2879(.a(G730), .O(gate242inter8));
  nand2 gate2880(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2881(.a(s_333), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2882(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2883(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2884(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1219(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1220(.a(gate243inter0), .b(s_96), .O(gate243inter1));
  and2  gate1221(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1222(.a(s_96), .O(gate243inter3));
  inv1  gate1223(.a(s_97), .O(gate243inter4));
  nand2 gate1224(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1225(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1226(.a(G245), .O(gate243inter7));
  inv1  gate1227(.a(G733), .O(gate243inter8));
  nand2 gate1228(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1229(.a(s_97), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1230(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1231(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1232(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2269(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2270(.a(gate245inter0), .b(s_246), .O(gate245inter1));
  and2  gate2271(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2272(.a(s_246), .O(gate245inter3));
  inv1  gate2273(.a(s_247), .O(gate245inter4));
  nand2 gate2274(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2275(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2276(.a(G248), .O(gate245inter7));
  inv1  gate2277(.a(G736), .O(gate245inter8));
  nand2 gate2278(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2279(.a(s_247), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2280(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2281(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2282(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1555(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1556(.a(gate250inter0), .b(s_144), .O(gate250inter1));
  and2  gate1557(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1558(.a(s_144), .O(gate250inter3));
  inv1  gate1559(.a(s_145), .O(gate250inter4));
  nand2 gate1560(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1561(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1562(.a(G706), .O(gate250inter7));
  inv1  gate1563(.a(G742), .O(gate250inter8));
  nand2 gate1564(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1565(.a(s_145), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1566(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1567(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1568(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1765(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1766(.a(gate253inter0), .b(s_174), .O(gate253inter1));
  and2  gate1767(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1768(.a(s_174), .O(gate253inter3));
  inv1  gate1769(.a(s_175), .O(gate253inter4));
  nand2 gate1770(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1771(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1772(.a(G260), .O(gate253inter7));
  inv1  gate1773(.a(G748), .O(gate253inter8));
  nand2 gate1774(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1775(.a(s_175), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1776(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1777(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1778(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2955(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2956(.a(gate256inter0), .b(s_344), .O(gate256inter1));
  and2  gate2957(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2958(.a(s_344), .O(gate256inter3));
  inv1  gate2959(.a(s_345), .O(gate256inter4));
  nand2 gate2960(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2961(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2962(.a(G715), .O(gate256inter7));
  inv1  gate2963(.a(G751), .O(gate256inter8));
  nand2 gate2964(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2965(.a(s_345), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2966(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2967(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2968(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate953(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate954(.a(gate257inter0), .b(s_58), .O(gate257inter1));
  and2  gate955(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate956(.a(s_58), .O(gate257inter3));
  inv1  gate957(.a(s_59), .O(gate257inter4));
  nand2 gate958(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate959(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate960(.a(G754), .O(gate257inter7));
  inv1  gate961(.a(G755), .O(gate257inter8));
  nand2 gate962(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate963(.a(s_59), .b(gate257inter3), .O(gate257inter10));
  nor2  gate964(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate965(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate966(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate2297(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2298(.a(gate258inter0), .b(s_250), .O(gate258inter1));
  and2  gate2299(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2300(.a(s_250), .O(gate258inter3));
  inv1  gate2301(.a(s_251), .O(gate258inter4));
  nand2 gate2302(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2303(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2304(.a(G756), .O(gate258inter7));
  inv1  gate2305(.a(G757), .O(gate258inter8));
  nand2 gate2306(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2307(.a(s_251), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2308(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2309(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2310(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate617(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate618(.a(gate259inter0), .b(s_10), .O(gate259inter1));
  and2  gate619(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate620(.a(s_10), .O(gate259inter3));
  inv1  gate621(.a(s_11), .O(gate259inter4));
  nand2 gate622(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate623(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate624(.a(G758), .O(gate259inter7));
  inv1  gate625(.a(G759), .O(gate259inter8));
  nand2 gate626(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate627(.a(s_11), .b(gate259inter3), .O(gate259inter10));
  nor2  gate628(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate629(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate630(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2451(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2452(.a(gate264inter0), .b(s_272), .O(gate264inter1));
  and2  gate2453(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2454(.a(s_272), .O(gate264inter3));
  inv1  gate2455(.a(s_273), .O(gate264inter4));
  nand2 gate2456(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2457(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2458(.a(G768), .O(gate264inter7));
  inv1  gate2459(.a(G769), .O(gate264inter8));
  nand2 gate2460(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2461(.a(s_273), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2462(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2463(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2464(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2087(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2088(.a(gate267inter0), .b(s_220), .O(gate267inter1));
  and2  gate2089(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2090(.a(s_220), .O(gate267inter3));
  inv1  gate2091(.a(s_221), .O(gate267inter4));
  nand2 gate2092(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2093(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2094(.a(G648), .O(gate267inter7));
  inv1  gate2095(.a(G776), .O(gate267inter8));
  nand2 gate2096(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2097(.a(s_221), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2098(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2099(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2100(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2885(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2886(.a(gate270inter0), .b(s_334), .O(gate270inter1));
  and2  gate2887(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2888(.a(s_334), .O(gate270inter3));
  inv1  gate2889(.a(s_335), .O(gate270inter4));
  nand2 gate2890(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2891(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2892(.a(G657), .O(gate270inter7));
  inv1  gate2893(.a(G785), .O(gate270inter8));
  nand2 gate2894(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2895(.a(s_335), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2896(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2897(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2898(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2003(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2004(.a(gate272inter0), .b(s_208), .O(gate272inter1));
  and2  gate2005(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2006(.a(s_208), .O(gate272inter3));
  inv1  gate2007(.a(s_209), .O(gate272inter4));
  nand2 gate2008(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2009(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2010(.a(G663), .O(gate272inter7));
  inv1  gate2011(.a(G791), .O(gate272inter8));
  nand2 gate2012(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2013(.a(s_209), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2014(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2015(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2016(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1513(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1514(.a(gate280inter0), .b(s_138), .O(gate280inter1));
  and2  gate1515(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1516(.a(s_138), .O(gate280inter3));
  inv1  gate1517(.a(s_139), .O(gate280inter4));
  nand2 gate1518(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1519(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1520(.a(G779), .O(gate280inter7));
  inv1  gate1521(.a(G803), .O(gate280inter8));
  nand2 gate1522(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1523(.a(s_139), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1524(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1525(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1526(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate2535(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2536(.a(gate281inter0), .b(s_284), .O(gate281inter1));
  and2  gate2537(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2538(.a(s_284), .O(gate281inter3));
  inv1  gate2539(.a(s_285), .O(gate281inter4));
  nand2 gate2540(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2541(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2542(.a(G654), .O(gate281inter7));
  inv1  gate2543(.a(G806), .O(gate281inter8));
  nand2 gate2544(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2545(.a(s_285), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2546(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2547(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2548(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2311(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2312(.a(gate283inter0), .b(s_252), .O(gate283inter1));
  and2  gate2313(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2314(.a(s_252), .O(gate283inter3));
  inv1  gate2315(.a(s_253), .O(gate283inter4));
  nand2 gate2316(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2317(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2318(.a(G657), .O(gate283inter7));
  inv1  gate2319(.a(G809), .O(gate283inter8));
  nand2 gate2320(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2321(.a(s_253), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2322(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2323(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2324(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1177(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1178(.a(gate287inter0), .b(s_90), .O(gate287inter1));
  and2  gate1179(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1180(.a(s_90), .O(gate287inter3));
  inv1  gate1181(.a(s_91), .O(gate287inter4));
  nand2 gate1182(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1183(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1184(.a(G663), .O(gate287inter7));
  inv1  gate1185(.a(G815), .O(gate287inter8));
  nand2 gate1186(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1187(.a(s_91), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1188(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1189(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1190(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1639(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1640(.a(gate288inter0), .b(s_156), .O(gate288inter1));
  and2  gate1641(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1642(.a(s_156), .O(gate288inter3));
  inv1  gate1643(.a(s_157), .O(gate288inter4));
  nand2 gate1644(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1645(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1646(.a(G791), .O(gate288inter7));
  inv1  gate1647(.a(G815), .O(gate288inter8));
  nand2 gate1648(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1649(.a(s_157), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1650(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1651(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1652(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1583(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1584(.a(gate289inter0), .b(s_148), .O(gate289inter1));
  and2  gate1585(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1586(.a(s_148), .O(gate289inter3));
  inv1  gate1587(.a(s_149), .O(gate289inter4));
  nand2 gate1588(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1589(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1590(.a(G818), .O(gate289inter7));
  inv1  gate1591(.a(G819), .O(gate289inter8));
  nand2 gate1592(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1593(.a(s_149), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1594(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1595(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1596(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2409(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2410(.a(gate292inter0), .b(s_266), .O(gate292inter1));
  and2  gate2411(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2412(.a(s_266), .O(gate292inter3));
  inv1  gate2413(.a(s_267), .O(gate292inter4));
  nand2 gate2414(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2415(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2416(.a(G824), .O(gate292inter7));
  inv1  gate2417(.a(G825), .O(gate292inter8));
  nand2 gate2418(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2419(.a(s_267), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2420(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2421(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2422(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate995(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate996(.a(gate295inter0), .b(s_64), .O(gate295inter1));
  and2  gate997(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate998(.a(s_64), .O(gate295inter3));
  inv1  gate999(.a(s_65), .O(gate295inter4));
  nand2 gate1000(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1001(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1002(.a(G830), .O(gate295inter7));
  inv1  gate1003(.a(G831), .O(gate295inter8));
  nand2 gate1004(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1005(.a(s_65), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1006(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1007(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1008(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1723(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1724(.a(gate296inter0), .b(s_168), .O(gate296inter1));
  and2  gate1725(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1726(.a(s_168), .O(gate296inter3));
  inv1  gate1727(.a(s_169), .O(gate296inter4));
  nand2 gate1728(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1729(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1730(.a(G826), .O(gate296inter7));
  inv1  gate1731(.a(G827), .O(gate296inter8));
  nand2 gate1732(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1733(.a(s_169), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1734(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1735(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1736(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1359(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1360(.a(gate391inter0), .b(s_116), .O(gate391inter1));
  and2  gate1361(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1362(.a(s_116), .O(gate391inter3));
  inv1  gate1363(.a(s_117), .O(gate391inter4));
  nand2 gate1364(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1365(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1366(.a(G5), .O(gate391inter7));
  inv1  gate1367(.a(G1048), .O(gate391inter8));
  nand2 gate1368(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1369(.a(s_117), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1370(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1371(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1372(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate3137(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate3138(.a(gate393inter0), .b(s_370), .O(gate393inter1));
  and2  gate3139(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate3140(.a(s_370), .O(gate393inter3));
  inv1  gate3141(.a(s_371), .O(gate393inter4));
  nand2 gate3142(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate3143(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate3144(.a(G7), .O(gate393inter7));
  inv1  gate3145(.a(G1054), .O(gate393inter8));
  nand2 gate3146(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate3147(.a(s_371), .b(gate393inter3), .O(gate393inter10));
  nor2  gate3148(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate3149(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate3150(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1107(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1108(.a(gate394inter0), .b(s_80), .O(gate394inter1));
  and2  gate1109(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1110(.a(s_80), .O(gate394inter3));
  inv1  gate1111(.a(s_81), .O(gate394inter4));
  nand2 gate1112(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1113(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1114(.a(G8), .O(gate394inter7));
  inv1  gate1115(.a(G1057), .O(gate394inter8));
  nand2 gate1116(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1117(.a(s_81), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1118(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1119(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1120(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate2339(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2340(.a(gate399inter0), .b(s_256), .O(gate399inter1));
  and2  gate2341(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2342(.a(s_256), .O(gate399inter3));
  inv1  gate2343(.a(s_257), .O(gate399inter4));
  nand2 gate2344(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2345(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2346(.a(G13), .O(gate399inter7));
  inv1  gate2347(.a(G1072), .O(gate399inter8));
  nand2 gate2348(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2349(.a(s_257), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2350(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2351(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2352(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1387(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1388(.a(gate401inter0), .b(s_120), .O(gate401inter1));
  and2  gate1389(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1390(.a(s_120), .O(gate401inter3));
  inv1  gate1391(.a(s_121), .O(gate401inter4));
  nand2 gate1392(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1393(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1394(.a(G15), .O(gate401inter7));
  inv1  gate1395(.a(G1078), .O(gate401inter8));
  nand2 gate1396(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1397(.a(s_121), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1398(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1399(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1400(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1569(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1570(.a(gate405inter0), .b(s_146), .O(gate405inter1));
  and2  gate1571(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1572(.a(s_146), .O(gate405inter3));
  inv1  gate1573(.a(s_147), .O(gate405inter4));
  nand2 gate1574(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1575(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1576(.a(G19), .O(gate405inter7));
  inv1  gate1577(.a(G1090), .O(gate405inter8));
  nand2 gate1578(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1579(.a(s_147), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1580(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1581(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1582(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1835(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1836(.a(gate406inter0), .b(s_184), .O(gate406inter1));
  and2  gate1837(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1838(.a(s_184), .O(gate406inter3));
  inv1  gate1839(.a(s_185), .O(gate406inter4));
  nand2 gate1840(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1841(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1842(.a(G20), .O(gate406inter7));
  inv1  gate1843(.a(G1093), .O(gate406inter8));
  nand2 gate1844(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1845(.a(s_185), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1846(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1847(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1848(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1891(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1892(.a(gate409inter0), .b(s_192), .O(gate409inter1));
  and2  gate1893(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1894(.a(s_192), .O(gate409inter3));
  inv1  gate1895(.a(s_193), .O(gate409inter4));
  nand2 gate1896(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1897(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1898(.a(G23), .O(gate409inter7));
  inv1  gate1899(.a(G1102), .O(gate409inter8));
  nand2 gate1900(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1901(.a(s_193), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1902(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1903(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1904(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate3095(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate3096(.a(gate411inter0), .b(s_364), .O(gate411inter1));
  and2  gate3097(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate3098(.a(s_364), .O(gate411inter3));
  inv1  gate3099(.a(s_365), .O(gate411inter4));
  nand2 gate3100(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate3101(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate3102(.a(G25), .O(gate411inter7));
  inv1  gate3103(.a(G1108), .O(gate411inter8));
  nand2 gate3104(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate3105(.a(s_365), .b(gate411inter3), .O(gate411inter10));
  nor2  gate3106(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate3107(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate3108(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1471(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1472(.a(gate412inter0), .b(s_132), .O(gate412inter1));
  and2  gate1473(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1474(.a(s_132), .O(gate412inter3));
  inv1  gate1475(.a(s_133), .O(gate412inter4));
  nand2 gate1476(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1477(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1478(.a(G26), .O(gate412inter7));
  inv1  gate1479(.a(G1111), .O(gate412inter8));
  nand2 gate1480(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1481(.a(s_133), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1482(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1483(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1484(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2479(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2480(.a(gate415inter0), .b(s_276), .O(gate415inter1));
  and2  gate2481(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2482(.a(s_276), .O(gate415inter3));
  inv1  gate2483(.a(s_277), .O(gate415inter4));
  nand2 gate2484(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2485(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2486(.a(G29), .O(gate415inter7));
  inv1  gate2487(.a(G1120), .O(gate415inter8));
  nand2 gate2488(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2489(.a(s_277), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2490(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2491(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2492(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1317(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1318(.a(gate419inter0), .b(s_110), .O(gate419inter1));
  and2  gate1319(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1320(.a(s_110), .O(gate419inter3));
  inv1  gate1321(.a(s_111), .O(gate419inter4));
  nand2 gate1322(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1323(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1324(.a(G1), .O(gate419inter7));
  inv1  gate1325(.a(G1132), .O(gate419inter8));
  nand2 gate1326(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1327(.a(s_111), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1328(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1329(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1330(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate575(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate576(.a(gate420inter0), .b(s_4), .O(gate420inter1));
  and2  gate577(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate578(.a(s_4), .O(gate420inter3));
  inv1  gate579(.a(s_5), .O(gate420inter4));
  nand2 gate580(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate581(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate582(.a(G1036), .O(gate420inter7));
  inv1  gate583(.a(G1132), .O(gate420inter8));
  nand2 gate584(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate585(.a(s_5), .b(gate420inter3), .O(gate420inter10));
  nor2  gate586(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate587(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate588(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1751(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1752(.a(gate423inter0), .b(s_172), .O(gate423inter1));
  and2  gate1753(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1754(.a(s_172), .O(gate423inter3));
  inv1  gate1755(.a(s_173), .O(gate423inter4));
  nand2 gate1756(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1757(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1758(.a(G3), .O(gate423inter7));
  inv1  gate1759(.a(G1138), .O(gate423inter8));
  nand2 gate1760(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1761(.a(s_173), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1762(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1763(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1764(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2199(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2200(.a(gate425inter0), .b(s_236), .O(gate425inter1));
  and2  gate2201(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2202(.a(s_236), .O(gate425inter3));
  inv1  gate2203(.a(s_237), .O(gate425inter4));
  nand2 gate2204(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2205(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2206(.a(G4), .O(gate425inter7));
  inv1  gate2207(.a(G1141), .O(gate425inter8));
  nand2 gate2208(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2209(.a(s_237), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2210(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2211(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2212(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate939(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate940(.a(gate426inter0), .b(s_56), .O(gate426inter1));
  and2  gate941(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate942(.a(s_56), .O(gate426inter3));
  inv1  gate943(.a(s_57), .O(gate426inter4));
  nand2 gate944(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate945(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate946(.a(G1045), .O(gate426inter7));
  inv1  gate947(.a(G1141), .O(gate426inter8));
  nand2 gate948(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate949(.a(s_57), .b(gate426inter3), .O(gate426inter10));
  nor2  gate950(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate951(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate952(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate729(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate730(.a(gate427inter0), .b(s_26), .O(gate427inter1));
  and2  gate731(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate732(.a(s_26), .O(gate427inter3));
  inv1  gate733(.a(s_27), .O(gate427inter4));
  nand2 gate734(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate735(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate736(.a(G5), .O(gate427inter7));
  inv1  gate737(.a(G1144), .O(gate427inter8));
  nand2 gate738(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate739(.a(s_27), .b(gate427inter3), .O(gate427inter10));
  nor2  gate740(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate741(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate742(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1373(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1374(.a(gate428inter0), .b(s_118), .O(gate428inter1));
  and2  gate1375(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1376(.a(s_118), .O(gate428inter3));
  inv1  gate1377(.a(s_119), .O(gate428inter4));
  nand2 gate1378(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1379(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1380(.a(G1048), .O(gate428inter7));
  inv1  gate1381(.a(G1144), .O(gate428inter8));
  nand2 gate1382(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1383(.a(s_119), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1384(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1385(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1386(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate2675(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2676(.a(gate429inter0), .b(s_304), .O(gate429inter1));
  and2  gate2677(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2678(.a(s_304), .O(gate429inter3));
  inv1  gate2679(.a(s_305), .O(gate429inter4));
  nand2 gate2680(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2681(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2682(.a(G6), .O(gate429inter7));
  inv1  gate2683(.a(G1147), .O(gate429inter8));
  nand2 gate2684(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2685(.a(s_305), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2686(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2687(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2688(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate757(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate758(.a(gate433inter0), .b(s_30), .O(gate433inter1));
  and2  gate759(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate760(.a(s_30), .O(gate433inter3));
  inv1  gate761(.a(s_31), .O(gate433inter4));
  nand2 gate762(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate763(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate764(.a(G8), .O(gate433inter7));
  inv1  gate765(.a(G1153), .O(gate433inter8));
  nand2 gate766(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate767(.a(s_31), .b(gate433inter3), .O(gate433inter10));
  nor2  gate768(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate769(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate770(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate645(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate646(.a(gate434inter0), .b(s_14), .O(gate434inter1));
  and2  gate647(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate648(.a(s_14), .O(gate434inter3));
  inv1  gate649(.a(s_15), .O(gate434inter4));
  nand2 gate650(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate651(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate652(.a(G1057), .O(gate434inter7));
  inv1  gate653(.a(G1153), .O(gate434inter8));
  nand2 gate654(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate655(.a(s_15), .b(gate434inter3), .O(gate434inter10));
  nor2  gate656(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate657(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate658(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate2437(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2438(.a(gate436inter0), .b(s_270), .O(gate436inter1));
  and2  gate2439(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2440(.a(s_270), .O(gate436inter3));
  inv1  gate2441(.a(s_271), .O(gate436inter4));
  nand2 gate2442(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2443(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2444(.a(G1060), .O(gate436inter7));
  inv1  gate2445(.a(G1156), .O(gate436inter8));
  nand2 gate2446(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2447(.a(s_271), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2448(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2449(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2450(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1163(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1164(.a(gate437inter0), .b(s_88), .O(gate437inter1));
  and2  gate1165(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1166(.a(s_88), .O(gate437inter3));
  inv1  gate1167(.a(s_89), .O(gate437inter4));
  nand2 gate1168(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1169(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1170(.a(G10), .O(gate437inter7));
  inv1  gate1171(.a(G1159), .O(gate437inter8));
  nand2 gate1172(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1173(.a(s_89), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1174(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1175(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1176(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2549(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2550(.a(gate438inter0), .b(s_286), .O(gate438inter1));
  and2  gate2551(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2552(.a(s_286), .O(gate438inter3));
  inv1  gate2553(.a(s_287), .O(gate438inter4));
  nand2 gate2554(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2555(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2556(.a(G1063), .O(gate438inter7));
  inv1  gate2557(.a(G1159), .O(gate438inter8));
  nand2 gate2558(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2559(.a(s_287), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2560(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2561(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2562(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate603(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate604(.a(gate443inter0), .b(s_8), .O(gate443inter1));
  and2  gate605(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate606(.a(s_8), .O(gate443inter3));
  inv1  gate607(.a(s_9), .O(gate443inter4));
  nand2 gate608(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate609(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate610(.a(G13), .O(gate443inter7));
  inv1  gate611(.a(G1168), .O(gate443inter8));
  nand2 gate612(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate613(.a(s_9), .b(gate443inter3), .O(gate443inter10));
  nor2  gate614(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate615(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate616(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate3053(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate3054(.a(gate446inter0), .b(s_358), .O(gate446inter1));
  and2  gate3055(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate3056(.a(s_358), .O(gate446inter3));
  inv1  gate3057(.a(s_359), .O(gate446inter4));
  nand2 gate3058(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate3059(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate3060(.a(G1075), .O(gate446inter7));
  inv1  gate3061(.a(G1171), .O(gate446inter8));
  nand2 gate3062(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate3063(.a(s_359), .b(gate446inter3), .O(gate446inter10));
  nor2  gate3064(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate3065(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate3066(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2031(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2032(.a(gate448inter0), .b(s_212), .O(gate448inter1));
  and2  gate2033(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2034(.a(s_212), .O(gate448inter3));
  inv1  gate2035(.a(s_213), .O(gate448inter4));
  nand2 gate2036(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2037(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2038(.a(G1078), .O(gate448inter7));
  inv1  gate2039(.a(G1174), .O(gate448inter8));
  nand2 gate2040(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2041(.a(s_213), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2042(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2043(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2044(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate715(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate716(.a(gate449inter0), .b(s_24), .O(gate449inter1));
  and2  gate717(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate718(.a(s_24), .O(gate449inter3));
  inv1  gate719(.a(s_25), .O(gate449inter4));
  nand2 gate720(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate721(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate722(.a(G16), .O(gate449inter7));
  inv1  gate723(.a(G1177), .O(gate449inter8));
  nand2 gate724(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate725(.a(s_25), .b(gate449inter3), .O(gate449inter10));
  nor2  gate726(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate727(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate728(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2899(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2900(.a(gate452inter0), .b(s_336), .O(gate452inter1));
  and2  gate2901(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2902(.a(s_336), .O(gate452inter3));
  inv1  gate2903(.a(s_337), .O(gate452inter4));
  nand2 gate2904(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2905(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2906(.a(G1084), .O(gate452inter7));
  inv1  gate2907(.a(G1180), .O(gate452inter8));
  nand2 gate2908(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2909(.a(s_337), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2910(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2911(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2912(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate3067(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate3068(.a(gate453inter0), .b(s_360), .O(gate453inter1));
  and2  gate3069(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate3070(.a(s_360), .O(gate453inter3));
  inv1  gate3071(.a(s_361), .O(gate453inter4));
  nand2 gate3072(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate3073(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate3074(.a(G18), .O(gate453inter7));
  inv1  gate3075(.a(G1183), .O(gate453inter8));
  nand2 gate3076(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate3077(.a(s_361), .b(gate453inter3), .O(gate453inter10));
  nor2  gate3078(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate3079(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate3080(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate3123(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate3124(.a(gate457inter0), .b(s_368), .O(gate457inter1));
  and2  gate3125(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate3126(.a(s_368), .O(gate457inter3));
  inv1  gate3127(.a(s_369), .O(gate457inter4));
  nand2 gate3128(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate3129(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate3130(.a(G20), .O(gate457inter7));
  inv1  gate3131(.a(G1189), .O(gate457inter8));
  nand2 gate3132(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate3133(.a(s_369), .b(gate457inter3), .O(gate457inter10));
  nor2  gate3134(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate3135(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate3136(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1037(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1038(.a(gate462inter0), .b(s_70), .O(gate462inter1));
  and2  gate1039(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1040(.a(s_70), .O(gate462inter3));
  inv1  gate1041(.a(s_71), .O(gate462inter4));
  nand2 gate1042(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1043(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1044(.a(G1099), .O(gate462inter7));
  inv1  gate1045(.a(G1195), .O(gate462inter8));
  nand2 gate1046(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1047(.a(s_71), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1048(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1049(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1050(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1737(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1738(.a(gate463inter0), .b(s_170), .O(gate463inter1));
  and2  gate1739(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1740(.a(s_170), .O(gate463inter3));
  inv1  gate1741(.a(s_171), .O(gate463inter4));
  nand2 gate1742(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1743(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1744(.a(G23), .O(gate463inter7));
  inv1  gate1745(.a(G1198), .O(gate463inter8));
  nand2 gate1746(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1747(.a(s_171), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1748(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1749(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1750(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate2507(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2508(.a(gate464inter0), .b(s_280), .O(gate464inter1));
  and2  gate2509(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2510(.a(s_280), .O(gate464inter3));
  inv1  gate2511(.a(s_281), .O(gate464inter4));
  nand2 gate2512(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2513(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2514(.a(G1102), .O(gate464inter7));
  inv1  gate2515(.a(G1198), .O(gate464inter8));
  nand2 gate2516(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2517(.a(s_281), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2518(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2519(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2520(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1653(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1654(.a(gate466inter0), .b(s_158), .O(gate466inter1));
  and2  gate1655(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1656(.a(s_158), .O(gate466inter3));
  inv1  gate1657(.a(s_159), .O(gate466inter4));
  nand2 gate1658(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1659(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1660(.a(G1105), .O(gate466inter7));
  inv1  gate1661(.a(G1201), .O(gate466inter8));
  nand2 gate1662(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1663(.a(s_159), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1664(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1665(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1666(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate2283(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2284(.a(gate468inter0), .b(s_248), .O(gate468inter1));
  and2  gate2285(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2286(.a(s_248), .O(gate468inter3));
  inv1  gate2287(.a(s_249), .O(gate468inter4));
  nand2 gate2288(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2289(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2290(.a(G1108), .O(gate468inter7));
  inv1  gate2291(.a(G1204), .O(gate468inter8));
  nand2 gate2292(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2293(.a(s_249), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2294(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2295(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2296(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate981(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate982(.a(gate469inter0), .b(s_62), .O(gate469inter1));
  and2  gate983(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate984(.a(s_62), .O(gate469inter3));
  inv1  gate985(.a(s_63), .O(gate469inter4));
  nand2 gate986(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate987(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate988(.a(G26), .O(gate469inter7));
  inv1  gate989(.a(G1207), .O(gate469inter8));
  nand2 gate990(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate991(.a(s_63), .b(gate469inter3), .O(gate469inter10));
  nor2  gate992(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate993(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate994(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2843(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2844(.a(gate472inter0), .b(s_328), .O(gate472inter1));
  and2  gate2845(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2846(.a(s_328), .O(gate472inter3));
  inv1  gate2847(.a(s_329), .O(gate472inter4));
  nand2 gate2848(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2849(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2850(.a(G1114), .O(gate472inter7));
  inv1  gate2851(.a(G1210), .O(gate472inter8));
  nand2 gate2852(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2853(.a(s_329), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2854(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2855(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2856(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate2773(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2774(.a(gate473inter0), .b(s_318), .O(gate473inter1));
  and2  gate2775(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2776(.a(s_318), .O(gate473inter3));
  inv1  gate2777(.a(s_319), .O(gate473inter4));
  nand2 gate2778(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2779(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2780(.a(G28), .O(gate473inter7));
  inv1  gate2781(.a(G1213), .O(gate473inter8));
  nand2 gate2782(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2783(.a(s_319), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2784(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2785(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2786(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate3081(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate3082(.a(gate477inter0), .b(s_362), .O(gate477inter1));
  and2  gate3083(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate3084(.a(s_362), .O(gate477inter3));
  inv1  gate3085(.a(s_363), .O(gate477inter4));
  nand2 gate3086(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate3087(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate3088(.a(G30), .O(gate477inter7));
  inv1  gate3089(.a(G1219), .O(gate477inter8));
  nand2 gate3090(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate3091(.a(s_363), .b(gate477inter3), .O(gate477inter10));
  nor2  gate3092(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate3093(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate3094(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1905(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1906(.a(gate481inter0), .b(s_194), .O(gate481inter1));
  and2  gate1907(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1908(.a(s_194), .O(gate481inter3));
  inv1  gate1909(.a(s_195), .O(gate481inter4));
  nand2 gate1910(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1911(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1912(.a(G32), .O(gate481inter7));
  inv1  gate1913(.a(G1225), .O(gate481inter8));
  nand2 gate1914(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1915(.a(s_195), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1916(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1917(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1918(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate673(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate674(.a(gate482inter0), .b(s_18), .O(gate482inter1));
  and2  gate675(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate676(.a(s_18), .O(gate482inter3));
  inv1  gate677(.a(s_19), .O(gate482inter4));
  nand2 gate678(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate679(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate680(.a(G1129), .O(gate482inter7));
  inv1  gate681(.a(G1225), .O(gate482inter8));
  nand2 gate682(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate683(.a(s_19), .b(gate482inter3), .O(gate482inter10));
  nor2  gate684(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate685(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate686(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1429(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1430(.a(gate483inter0), .b(s_126), .O(gate483inter1));
  and2  gate1431(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1432(.a(s_126), .O(gate483inter3));
  inv1  gate1433(.a(s_127), .O(gate483inter4));
  nand2 gate1434(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1435(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1436(.a(G1228), .O(gate483inter7));
  inv1  gate1437(.a(G1229), .O(gate483inter8));
  nand2 gate1438(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1439(.a(s_127), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1440(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1441(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1442(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2157(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2158(.a(gate488inter0), .b(s_230), .O(gate488inter1));
  and2  gate2159(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2160(.a(s_230), .O(gate488inter3));
  inv1  gate2161(.a(s_231), .O(gate488inter4));
  nand2 gate2162(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2163(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2164(.a(G1238), .O(gate488inter7));
  inv1  gate2165(.a(G1239), .O(gate488inter8));
  nand2 gate2166(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2167(.a(s_231), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2168(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2169(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2170(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1695(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1696(.a(gate489inter0), .b(s_164), .O(gate489inter1));
  and2  gate1697(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1698(.a(s_164), .O(gate489inter3));
  inv1  gate1699(.a(s_165), .O(gate489inter4));
  nand2 gate1700(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1701(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1702(.a(G1240), .O(gate489inter7));
  inv1  gate1703(.a(G1241), .O(gate489inter8));
  nand2 gate1704(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1705(.a(s_165), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1706(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1707(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1708(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1499(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1500(.a(gate490inter0), .b(s_136), .O(gate490inter1));
  and2  gate1501(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1502(.a(s_136), .O(gate490inter3));
  inv1  gate1503(.a(s_137), .O(gate490inter4));
  nand2 gate1504(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1505(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1506(.a(G1242), .O(gate490inter7));
  inv1  gate1507(.a(G1243), .O(gate490inter8));
  nand2 gate1508(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1509(.a(s_137), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1510(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1511(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1512(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate827(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate828(.a(gate492inter0), .b(s_40), .O(gate492inter1));
  and2  gate829(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate830(.a(s_40), .O(gate492inter3));
  inv1  gate831(.a(s_41), .O(gate492inter4));
  nand2 gate832(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate833(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate834(.a(G1246), .O(gate492inter7));
  inv1  gate835(.a(G1247), .O(gate492inter8));
  nand2 gate836(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate837(.a(s_41), .b(gate492inter3), .O(gate492inter10));
  nor2  gate838(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate839(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate840(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2521(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2522(.a(gate493inter0), .b(s_282), .O(gate493inter1));
  and2  gate2523(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2524(.a(s_282), .O(gate493inter3));
  inv1  gate2525(.a(s_283), .O(gate493inter4));
  nand2 gate2526(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2527(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2528(.a(G1248), .O(gate493inter7));
  inv1  gate2529(.a(G1249), .O(gate493inter8));
  nand2 gate2530(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2531(.a(s_283), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2532(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2533(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2534(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2591(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2592(.a(gate494inter0), .b(s_292), .O(gate494inter1));
  and2  gate2593(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2594(.a(s_292), .O(gate494inter3));
  inv1  gate2595(.a(s_293), .O(gate494inter4));
  nand2 gate2596(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2597(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2598(.a(G1250), .O(gate494inter7));
  inv1  gate2599(.a(G1251), .O(gate494inter8));
  nand2 gate2600(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2601(.a(s_293), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2602(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2603(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2604(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1947(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1948(.a(gate495inter0), .b(s_200), .O(gate495inter1));
  and2  gate1949(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1950(.a(s_200), .O(gate495inter3));
  inv1  gate1951(.a(s_201), .O(gate495inter4));
  nand2 gate1952(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1953(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1954(.a(G1252), .O(gate495inter7));
  inv1  gate1955(.a(G1253), .O(gate495inter8));
  nand2 gate1956(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1957(.a(s_201), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1958(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1959(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1960(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2171(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2172(.a(gate497inter0), .b(s_232), .O(gate497inter1));
  and2  gate2173(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2174(.a(s_232), .O(gate497inter3));
  inv1  gate2175(.a(s_233), .O(gate497inter4));
  nand2 gate2176(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2177(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2178(.a(G1256), .O(gate497inter7));
  inv1  gate2179(.a(G1257), .O(gate497inter8));
  nand2 gate2180(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2181(.a(s_233), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2182(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2183(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2184(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate701(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate702(.a(gate500inter0), .b(s_22), .O(gate500inter1));
  and2  gate703(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate704(.a(s_22), .O(gate500inter3));
  inv1  gate705(.a(s_23), .O(gate500inter4));
  nand2 gate706(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate707(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate708(.a(G1262), .O(gate500inter7));
  inv1  gate709(.a(G1263), .O(gate500inter8));
  nand2 gate710(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate711(.a(s_23), .b(gate500inter3), .O(gate500inter10));
  nor2  gate712(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate713(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate714(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1877(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1878(.a(gate506inter0), .b(s_190), .O(gate506inter1));
  and2  gate1879(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1880(.a(s_190), .O(gate506inter3));
  inv1  gate1881(.a(s_191), .O(gate506inter4));
  nand2 gate1882(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1883(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1884(.a(G1274), .O(gate506inter7));
  inv1  gate1885(.a(G1275), .O(gate506inter8));
  nand2 gate1886(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1887(.a(s_191), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1888(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1889(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1890(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1709(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1710(.a(gate507inter0), .b(s_166), .O(gate507inter1));
  and2  gate1711(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1712(.a(s_166), .O(gate507inter3));
  inv1  gate1713(.a(s_167), .O(gate507inter4));
  nand2 gate1714(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1715(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1716(.a(G1276), .O(gate507inter7));
  inv1  gate1717(.a(G1277), .O(gate507inter8));
  nand2 gate1718(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1719(.a(s_167), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1720(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1721(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1722(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2213(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2214(.a(gate509inter0), .b(s_238), .O(gate509inter1));
  and2  gate2215(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2216(.a(s_238), .O(gate509inter3));
  inv1  gate2217(.a(s_239), .O(gate509inter4));
  nand2 gate2218(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2219(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2220(.a(G1280), .O(gate509inter7));
  inv1  gate2221(.a(G1281), .O(gate509inter8));
  nand2 gate2222(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2223(.a(s_239), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2224(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2225(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2226(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2689(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2690(.a(gate511inter0), .b(s_306), .O(gate511inter1));
  and2  gate2691(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2692(.a(s_306), .O(gate511inter3));
  inv1  gate2693(.a(s_307), .O(gate511inter4));
  nand2 gate2694(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2695(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2696(.a(G1284), .O(gate511inter7));
  inv1  gate2697(.a(G1285), .O(gate511inter8));
  nand2 gate2698(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2699(.a(s_307), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2700(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2701(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2702(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate2059(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2060(.a(gate512inter0), .b(s_216), .O(gate512inter1));
  and2  gate2061(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2062(.a(s_216), .O(gate512inter3));
  inv1  gate2063(.a(s_217), .O(gate512inter4));
  nand2 gate2064(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2065(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2066(.a(G1286), .O(gate512inter7));
  inv1  gate2067(.a(G1287), .O(gate512inter8));
  nand2 gate2068(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2069(.a(s_217), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2070(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2071(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2072(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate2619(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2620(.a(gate513inter0), .b(s_296), .O(gate513inter1));
  and2  gate2621(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2622(.a(s_296), .O(gate513inter3));
  inv1  gate2623(.a(s_297), .O(gate513inter4));
  nand2 gate2624(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2625(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2626(.a(G1288), .O(gate513inter7));
  inv1  gate2627(.a(G1289), .O(gate513inter8));
  nand2 gate2628(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2629(.a(s_297), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2630(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2631(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2632(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule