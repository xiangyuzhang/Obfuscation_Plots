module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1541(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1542(.a(gate9inter0), .b(s_142), .O(gate9inter1));
  and2  gate1543(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1544(.a(s_142), .O(gate9inter3));
  inv1  gate1545(.a(s_143), .O(gate9inter4));
  nand2 gate1546(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1547(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1548(.a(G1), .O(gate9inter7));
  inv1  gate1549(.a(G2), .O(gate9inter8));
  nand2 gate1550(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1551(.a(s_143), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1552(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1553(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1554(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1345(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1346(.a(gate12inter0), .b(s_114), .O(gate12inter1));
  and2  gate1347(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1348(.a(s_114), .O(gate12inter3));
  inv1  gate1349(.a(s_115), .O(gate12inter4));
  nand2 gate1350(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1351(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1352(.a(G7), .O(gate12inter7));
  inv1  gate1353(.a(G8), .O(gate12inter8));
  nand2 gate1354(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1355(.a(s_115), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1356(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1357(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1358(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate883(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate884(.a(gate13inter0), .b(s_48), .O(gate13inter1));
  and2  gate885(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate886(.a(s_48), .O(gate13inter3));
  inv1  gate887(.a(s_49), .O(gate13inter4));
  nand2 gate888(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate889(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate890(.a(G9), .O(gate13inter7));
  inv1  gate891(.a(G10), .O(gate13inter8));
  nand2 gate892(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate893(.a(s_49), .b(gate13inter3), .O(gate13inter10));
  nor2  gate894(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate895(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate896(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1457(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1458(.a(gate14inter0), .b(s_130), .O(gate14inter1));
  and2  gate1459(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1460(.a(s_130), .O(gate14inter3));
  inv1  gate1461(.a(s_131), .O(gate14inter4));
  nand2 gate1462(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1463(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1464(.a(G11), .O(gate14inter7));
  inv1  gate1465(.a(G12), .O(gate14inter8));
  nand2 gate1466(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1467(.a(s_131), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1468(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1469(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1470(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate841(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate842(.a(gate16inter0), .b(s_42), .O(gate16inter1));
  and2  gate843(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate844(.a(s_42), .O(gate16inter3));
  inv1  gate845(.a(s_43), .O(gate16inter4));
  nand2 gate846(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate847(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate848(.a(G15), .O(gate16inter7));
  inv1  gate849(.a(G16), .O(gate16inter8));
  nand2 gate850(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate851(.a(s_43), .b(gate16inter3), .O(gate16inter10));
  nor2  gate852(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate853(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate854(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1639(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1640(.a(gate18inter0), .b(s_156), .O(gate18inter1));
  and2  gate1641(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1642(.a(s_156), .O(gate18inter3));
  inv1  gate1643(.a(s_157), .O(gate18inter4));
  nand2 gate1644(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1645(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1646(.a(G19), .O(gate18inter7));
  inv1  gate1647(.a(G20), .O(gate18inter8));
  nand2 gate1648(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1649(.a(s_157), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1650(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1651(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1652(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate855(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate856(.a(gate19inter0), .b(s_44), .O(gate19inter1));
  and2  gate857(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate858(.a(s_44), .O(gate19inter3));
  inv1  gate859(.a(s_45), .O(gate19inter4));
  nand2 gate860(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate861(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate862(.a(G21), .O(gate19inter7));
  inv1  gate863(.a(G22), .O(gate19inter8));
  nand2 gate864(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate865(.a(s_45), .b(gate19inter3), .O(gate19inter10));
  nor2  gate866(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate867(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate868(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1513(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1514(.a(gate20inter0), .b(s_138), .O(gate20inter1));
  and2  gate1515(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1516(.a(s_138), .O(gate20inter3));
  inv1  gate1517(.a(s_139), .O(gate20inter4));
  nand2 gate1518(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1519(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1520(.a(G23), .O(gate20inter7));
  inv1  gate1521(.a(G24), .O(gate20inter8));
  nand2 gate1522(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1523(.a(s_139), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1524(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1525(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1526(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1303(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1304(.a(gate22inter0), .b(s_108), .O(gate22inter1));
  and2  gate1305(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1306(.a(s_108), .O(gate22inter3));
  inv1  gate1307(.a(s_109), .O(gate22inter4));
  nand2 gate1308(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1309(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1310(.a(G27), .O(gate22inter7));
  inv1  gate1311(.a(G28), .O(gate22inter8));
  nand2 gate1312(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1313(.a(s_109), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1314(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1315(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1316(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate631(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate632(.a(gate25inter0), .b(s_12), .O(gate25inter1));
  and2  gate633(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate634(.a(s_12), .O(gate25inter3));
  inv1  gate635(.a(s_13), .O(gate25inter4));
  nand2 gate636(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate637(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate638(.a(G1), .O(gate25inter7));
  inv1  gate639(.a(G5), .O(gate25inter8));
  nand2 gate640(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate641(.a(s_13), .b(gate25inter3), .O(gate25inter10));
  nor2  gate642(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate643(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate644(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1065(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1066(.a(gate28inter0), .b(s_74), .O(gate28inter1));
  and2  gate1067(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1068(.a(s_74), .O(gate28inter3));
  inv1  gate1069(.a(s_75), .O(gate28inter4));
  nand2 gate1070(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1071(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1072(.a(G10), .O(gate28inter7));
  inv1  gate1073(.a(G14), .O(gate28inter8));
  nand2 gate1074(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1075(.a(s_75), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1076(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1077(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1078(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1107(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1108(.a(gate33inter0), .b(s_80), .O(gate33inter1));
  and2  gate1109(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1110(.a(s_80), .O(gate33inter3));
  inv1  gate1111(.a(s_81), .O(gate33inter4));
  nand2 gate1112(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1113(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1114(.a(G17), .O(gate33inter7));
  inv1  gate1115(.a(G21), .O(gate33inter8));
  nand2 gate1116(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1117(.a(s_81), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1118(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1119(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1120(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2003(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2004(.a(gate43inter0), .b(s_208), .O(gate43inter1));
  and2  gate2005(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2006(.a(s_208), .O(gate43inter3));
  inv1  gate2007(.a(s_209), .O(gate43inter4));
  nand2 gate2008(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2009(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2010(.a(G3), .O(gate43inter7));
  inv1  gate2011(.a(G269), .O(gate43inter8));
  nand2 gate2012(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2013(.a(s_209), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2014(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2015(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2016(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1723(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1724(.a(gate44inter0), .b(s_168), .O(gate44inter1));
  and2  gate1725(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1726(.a(s_168), .O(gate44inter3));
  inv1  gate1727(.a(s_169), .O(gate44inter4));
  nand2 gate1728(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1729(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1730(.a(G4), .O(gate44inter7));
  inv1  gate1731(.a(G269), .O(gate44inter8));
  nand2 gate1732(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1733(.a(s_169), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1734(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1735(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1736(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1667(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1668(.a(gate46inter0), .b(s_160), .O(gate46inter1));
  and2  gate1669(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1670(.a(s_160), .O(gate46inter3));
  inv1  gate1671(.a(s_161), .O(gate46inter4));
  nand2 gate1672(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1673(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1674(.a(G6), .O(gate46inter7));
  inv1  gate1675(.a(G272), .O(gate46inter8));
  nand2 gate1676(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1677(.a(s_161), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1678(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1679(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1680(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1653(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1654(.a(gate47inter0), .b(s_158), .O(gate47inter1));
  and2  gate1655(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1656(.a(s_158), .O(gate47inter3));
  inv1  gate1657(.a(s_159), .O(gate47inter4));
  nand2 gate1658(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1659(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1660(.a(G7), .O(gate47inter7));
  inv1  gate1661(.a(G275), .O(gate47inter8));
  nand2 gate1662(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1663(.a(s_159), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1664(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1665(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1666(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate603(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate604(.a(gate49inter0), .b(s_8), .O(gate49inter1));
  and2  gate605(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate606(.a(s_8), .O(gate49inter3));
  inv1  gate607(.a(s_9), .O(gate49inter4));
  nand2 gate608(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate609(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate610(.a(G9), .O(gate49inter7));
  inv1  gate611(.a(G278), .O(gate49inter8));
  nand2 gate612(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate613(.a(s_9), .b(gate49inter3), .O(gate49inter10));
  nor2  gate614(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate615(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate616(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1037(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1038(.a(gate51inter0), .b(s_70), .O(gate51inter1));
  and2  gate1039(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1040(.a(s_70), .O(gate51inter3));
  inv1  gate1041(.a(s_71), .O(gate51inter4));
  nand2 gate1042(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1043(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1044(.a(G11), .O(gate51inter7));
  inv1  gate1045(.a(G281), .O(gate51inter8));
  nand2 gate1046(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1047(.a(s_71), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1048(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1049(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1050(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate2031(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2032(.a(gate52inter0), .b(s_212), .O(gate52inter1));
  and2  gate2033(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2034(.a(s_212), .O(gate52inter3));
  inv1  gate2035(.a(s_213), .O(gate52inter4));
  nand2 gate2036(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2037(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2038(.a(G12), .O(gate52inter7));
  inv1  gate2039(.a(G281), .O(gate52inter8));
  nand2 gate2040(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2041(.a(s_213), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2042(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2043(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2044(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2073(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2074(.a(gate55inter0), .b(s_218), .O(gate55inter1));
  and2  gate2075(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2076(.a(s_218), .O(gate55inter3));
  inv1  gate2077(.a(s_219), .O(gate55inter4));
  nand2 gate2078(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2079(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2080(.a(G15), .O(gate55inter7));
  inv1  gate2081(.a(G287), .O(gate55inter8));
  nand2 gate2082(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2083(.a(s_219), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2084(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2085(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2086(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1527(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1528(.a(gate58inter0), .b(s_140), .O(gate58inter1));
  and2  gate1529(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1530(.a(s_140), .O(gate58inter3));
  inv1  gate1531(.a(s_141), .O(gate58inter4));
  nand2 gate1532(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1533(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1534(.a(G18), .O(gate58inter7));
  inv1  gate1535(.a(G290), .O(gate58inter8));
  nand2 gate1536(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1537(.a(s_141), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1538(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1539(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1540(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1681(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1682(.a(gate62inter0), .b(s_162), .O(gate62inter1));
  and2  gate1683(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1684(.a(s_162), .O(gate62inter3));
  inv1  gate1685(.a(s_163), .O(gate62inter4));
  nand2 gate1686(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1687(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1688(.a(G22), .O(gate62inter7));
  inv1  gate1689(.a(G296), .O(gate62inter8));
  nand2 gate1690(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1691(.a(s_163), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1692(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1693(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1694(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1191(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1192(.a(gate64inter0), .b(s_92), .O(gate64inter1));
  and2  gate1193(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1194(.a(s_92), .O(gate64inter3));
  inv1  gate1195(.a(s_93), .O(gate64inter4));
  nand2 gate1196(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1197(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1198(.a(G24), .O(gate64inter7));
  inv1  gate1199(.a(G299), .O(gate64inter8));
  nand2 gate1200(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1201(.a(s_93), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1202(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1203(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1204(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1695(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1696(.a(gate67inter0), .b(s_164), .O(gate67inter1));
  and2  gate1697(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1698(.a(s_164), .O(gate67inter3));
  inv1  gate1699(.a(s_165), .O(gate67inter4));
  nand2 gate1700(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1701(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1702(.a(G27), .O(gate67inter7));
  inv1  gate1703(.a(G305), .O(gate67inter8));
  nand2 gate1704(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1705(.a(s_165), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1706(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1707(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1708(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate967(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate968(.a(gate68inter0), .b(s_60), .O(gate68inter1));
  and2  gate969(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate970(.a(s_60), .O(gate68inter3));
  inv1  gate971(.a(s_61), .O(gate68inter4));
  nand2 gate972(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate973(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate974(.a(G28), .O(gate68inter7));
  inv1  gate975(.a(G305), .O(gate68inter8));
  nand2 gate976(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate977(.a(s_61), .b(gate68inter3), .O(gate68inter10));
  nor2  gate978(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate979(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate980(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate589(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate590(.a(gate71inter0), .b(s_6), .O(gate71inter1));
  and2  gate591(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate592(.a(s_6), .O(gate71inter3));
  inv1  gate593(.a(s_7), .O(gate71inter4));
  nand2 gate594(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate595(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate596(.a(G31), .O(gate71inter7));
  inv1  gate597(.a(G311), .O(gate71inter8));
  nand2 gate598(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate599(.a(s_7), .b(gate71inter3), .O(gate71inter10));
  nor2  gate600(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate601(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate602(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate757(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate758(.a(gate74inter0), .b(s_30), .O(gate74inter1));
  and2  gate759(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate760(.a(s_30), .O(gate74inter3));
  inv1  gate761(.a(s_31), .O(gate74inter4));
  nand2 gate762(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate763(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate764(.a(G5), .O(gate74inter7));
  inv1  gate765(.a(G314), .O(gate74inter8));
  nand2 gate766(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate767(.a(s_31), .b(gate74inter3), .O(gate74inter10));
  nor2  gate768(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate769(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate770(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate827(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate828(.a(gate77inter0), .b(s_40), .O(gate77inter1));
  and2  gate829(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate830(.a(s_40), .O(gate77inter3));
  inv1  gate831(.a(s_41), .O(gate77inter4));
  nand2 gate832(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate833(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate834(.a(G2), .O(gate77inter7));
  inv1  gate835(.a(G320), .O(gate77inter8));
  nand2 gate836(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate837(.a(s_41), .b(gate77inter3), .O(gate77inter10));
  nor2  gate838(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate839(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate840(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1163(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1164(.a(gate79inter0), .b(s_88), .O(gate79inter1));
  and2  gate1165(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1166(.a(s_88), .O(gate79inter3));
  inv1  gate1167(.a(s_89), .O(gate79inter4));
  nand2 gate1168(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1169(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1170(.a(G10), .O(gate79inter7));
  inv1  gate1171(.a(G323), .O(gate79inter8));
  nand2 gate1172(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1173(.a(s_89), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1174(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1175(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1176(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1821(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1822(.a(gate81inter0), .b(s_182), .O(gate81inter1));
  and2  gate1823(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1824(.a(s_182), .O(gate81inter3));
  inv1  gate1825(.a(s_183), .O(gate81inter4));
  nand2 gate1826(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1827(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1828(.a(G3), .O(gate81inter7));
  inv1  gate1829(.a(G326), .O(gate81inter8));
  nand2 gate1830(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1831(.a(s_183), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1832(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1833(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1834(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1387(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1388(.a(gate86inter0), .b(s_120), .O(gate86inter1));
  and2  gate1389(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1390(.a(s_120), .O(gate86inter3));
  inv1  gate1391(.a(s_121), .O(gate86inter4));
  nand2 gate1392(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1393(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1394(.a(G8), .O(gate86inter7));
  inv1  gate1395(.a(G332), .O(gate86inter8));
  nand2 gate1396(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1397(.a(s_121), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1398(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1399(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1400(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1009(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1010(.a(gate91inter0), .b(s_66), .O(gate91inter1));
  and2  gate1011(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1012(.a(s_66), .O(gate91inter3));
  inv1  gate1013(.a(s_67), .O(gate91inter4));
  nand2 gate1014(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1015(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1016(.a(G25), .O(gate91inter7));
  inv1  gate1017(.a(G341), .O(gate91inter8));
  nand2 gate1018(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1019(.a(s_67), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1020(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1021(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1022(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2017(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2018(.a(gate94inter0), .b(s_210), .O(gate94inter1));
  and2  gate2019(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2020(.a(s_210), .O(gate94inter3));
  inv1  gate2021(.a(s_211), .O(gate94inter4));
  nand2 gate2022(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2023(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2024(.a(G22), .O(gate94inter7));
  inv1  gate2025(.a(G344), .O(gate94inter8));
  nand2 gate2026(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2027(.a(s_211), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2028(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2029(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2030(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1429(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1430(.a(gate95inter0), .b(s_126), .O(gate95inter1));
  and2  gate1431(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1432(.a(s_126), .O(gate95inter3));
  inv1  gate1433(.a(s_127), .O(gate95inter4));
  nand2 gate1434(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1435(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1436(.a(G26), .O(gate95inter7));
  inv1  gate1437(.a(G347), .O(gate95inter8));
  nand2 gate1438(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1439(.a(s_127), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1440(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1441(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1442(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1135(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1136(.a(gate99inter0), .b(s_84), .O(gate99inter1));
  and2  gate1137(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1138(.a(s_84), .O(gate99inter3));
  inv1  gate1139(.a(s_85), .O(gate99inter4));
  nand2 gate1140(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1141(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1142(.a(G27), .O(gate99inter7));
  inv1  gate1143(.a(G353), .O(gate99inter8));
  nand2 gate1144(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1145(.a(s_85), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1146(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1147(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1148(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate729(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate730(.a(gate101inter0), .b(s_26), .O(gate101inter1));
  and2  gate731(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate732(.a(s_26), .O(gate101inter3));
  inv1  gate733(.a(s_27), .O(gate101inter4));
  nand2 gate734(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate735(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate736(.a(G20), .O(gate101inter7));
  inv1  gate737(.a(G356), .O(gate101inter8));
  nand2 gate738(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate739(.a(s_27), .b(gate101inter3), .O(gate101inter10));
  nor2  gate740(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate741(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate742(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate715(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate716(.a(gate110inter0), .b(s_24), .O(gate110inter1));
  and2  gate717(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate718(.a(s_24), .O(gate110inter3));
  inv1  gate719(.a(s_25), .O(gate110inter4));
  nand2 gate720(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate721(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate722(.a(G372), .O(gate110inter7));
  inv1  gate723(.a(G373), .O(gate110inter8));
  nand2 gate724(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate725(.a(s_25), .b(gate110inter3), .O(gate110inter10));
  nor2  gate726(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate727(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate728(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate925(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate926(.a(gate112inter0), .b(s_54), .O(gate112inter1));
  and2  gate927(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate928(.a(s_54), .O(gate112inter3));
  inv1  gate929(.a(s_55), .O(gate112inter4));
  nand2 gate930(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate931(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate932(.a(G376), .O(gate112inter7));
  inv1  gate933(.a(G377), .O(gate112inter8));
  nand2 gate934(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate935(.a(s_55), .b(gate112inter3), .O(gate112inter10));
  nor2  gate936(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate937(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate938(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1023(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1024(.a(gate115inter0), .b(s_68), .O(gate115inter1));
  and2  gate1025(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1026(.a(s_68), .O(gate115inter3));
  inv1  gate1027(.a(s_69), .O(gate115inter4));
  nand2 gate1028(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1029(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1030(.a(G382), .O(gate115inter7));
  inv1  gate1031(.a(G383), .O(gate115inter8));
  nand2 gate1032(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1033(.a(s_69), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1034(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1035(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1036(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate701(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate702(.a(gate119inter0), .b(s_22), .O(gate119inter1));
  and2  gate703(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate704(.a(s_22), .O(gate119inter3));
  inv1  gate705(.a(s_23), .O(gate119inter4));
  nand2 gate706(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate707(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate708(.a(G390), .O(gate119inter7));
  inv1  gate709(.a(G391), .O(gate119inter8));
  nand2 gate710(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate711(.a(s_23), .b(gate119inter3), .O(gate119inter10));
  nor2  gate712(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate713(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate714(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1121(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1122(.a(gate128inter0), .b(s_82), .O(gate128inter1));
  and2  gate1123(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1124(.a(s_82), .O(gate128inter3));
  inv1  gate1125(.a(s_83), .O(gate128inter4));
  nand2 gate1126(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1127(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1128(.a(G408), .O(gate128inter7));
  inv1  gate1129(.a(G409), .O(gate128inter8));
  nand2 gate1130(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1131(.a(s_83), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1132(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1133(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1134(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1975(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1976(.a(gate129inter0), .b(s_204), .O(gate129inter1));
  and2  gate1977(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1978(.a(s_204), .O(gate129inter3));
  inv1  gate1979(.a(s_205), .O(gate129inter4));
  nand2 gate1980(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1981(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1982(.a(G410), .O(gate129inter7));
  inv1  gate1983(.a(G411), .O(gate129inter8));
  nand2 gate1984(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1985(.a(s_205), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1986(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1987(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1988(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate799(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate800(.a(gate131inter0), .b(s_36), .O(gate131inter1));
  and2  gate801(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate802(.a(s_36), .O(gate131inter3));
  inv1  gate803(.a(s_37), .O(gate131inter4));
  nand2 gate804(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate805(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate806(.a(G414), .O(gate131inter7));
  inv1  gate807(.a(G415), .O(gate131inter8));
  nand2 gate808(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate809(.a(s_37), .b(gate131inter3), .O(gate131inter10));
  nor2  gate810(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate811(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate812(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate911(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate912(.a(gate133inter0), .b(s_52), .O(gate133inter1));
  and2  gate913(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate914(.a(s_52), .O(gate133inter3));
  inv1  gate915(.a(s_53), .O(gate133inter4));
  nand2 gate916(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate917(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate918(.a(G418), .O(gate133inter7));
  inv1  gate919(.a(G419), .O(gate133inter8));
  nand2 gate920(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate921(.a(s_53), .b(gate133inter3), .O(gate133inter10));
  nor2  gate922(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate923(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate924(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1611(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1612(.a(gate136inter0), .b(s_152), .O(gate136inter1));
  and2  gate1613(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1614(.a(s_152), .O(gate136inter3));
  inv1  gate1615(.a(s_153), .O(gate136inter4));
  nand2 gate1616(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1617(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1618(.a(G424), .O(gate136inter7));
  inv1  gate1619(.a(G425), .O(gate136inter8));
  nand2 gate1620(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1621(.a(s_153), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1622(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1623(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1624(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate547(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate548(.a(gate141inter0), .b(s_0), .O(gate141inter1));
  and2  gate549(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate550(.a(s_0), .O(gate141inter3));
  inv1  gate551(.a(s_1), .O(gate141inter4));
  nand2 gate552(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate553(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate554(.a(G450), .O(gate141inter7));
  inv1  gate555(.a(G453), .O(gate141inter8));
  nand2 gate556(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate557(.a(s_1), .b(gate141inter3), .O(gate141inter10));
  nor2  gate558(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate559(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate560(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1079(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1080(.a(gate144inter0), .b(s_76), .O(gate144inter1));
  and2  gate1081(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1082(.a(s_76), .O(gate144inter3));
  inv1  gate1083(.a(s_77), .O(gate144inter4));
  nand2 gate1084(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1085(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1086(.a(G468), .O(gate144inter7));
  inv1  gate1087(.a(G471), .O(gate144inter8));
  nand2 gate1088(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1089(.a(s_77), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1090(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1091(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1092(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1919(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1920(.a(gate147inter0), .b(s_196), .O(gate147inter1));
  and2  gate1921(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1922(.a(s_196), .O(gate147inter3));
  inv1  gate1923(.a(s_197), .O(gate147inter4));
  nand2 gate1924(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1925(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1926(.a(G486), .O(gate147inter7));
  inv1  gate1927(.a(G489), .O(gate147inter8));
  nand2 gate1928(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1929(.a(s_197), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1930(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1931(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1932(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1737(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1738(.a(gate153inter0), .b(s_170), .O(gate153inter1));
  and2  gate1739(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1740(.a(s_170), .O(gate153inter3));
  inv1  gate1741(.a(s_171), .O(gate153inter4));
  nand2 gate1742(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1743(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1744(.a(G426), .O(gate153inter7));
  inv1  gate1745(.a(G522), .O(gate153inter8));
  nand2 gate1746(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1747(.a(s_171), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1748(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1749(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1750(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1359(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1360(.a(gate154inter0), .b(s_116), .O(gate154inter1));
  and2  gate1361(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1362(.a(s_116), .O(gate154inter3));
  inv1  gate1363(.a(s_117), .O(gate154inter4));
  nand2 gate1364(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1365(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1366(.a(G429), .O(gate154inter7));
  inv1  gate1367(.a(G522), .O(gate154inter8));
  nand2 gate1368(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1369(.a(s_117), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1370(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1371(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1372(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate687(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate688(.a(gate156inter0), .b(s_20), .O(gate156inter1));
  and2  gate689(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate690(.a(s_20), .O(gate156inter3));
  inv1  gate691(.a(s_21), .O(gate156inter4));
  nand2 gate692(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate693(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate694(.a(G435), .O(gate156inter7));
  inv1  gate695(.a(G525), .O(gate156inter8));
  nand2 gate696(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate697(.a(s_21), .b(gate156inter3), .O(gate156inter10));
  nor2  gate698(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate699(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate700(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2087(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2088(.a(gate165inter0), .b(s_220), .O(gate165inter1));
  and2  gate2089(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2090(.a(s_220), .O(gate165inter3));
  inv1  gate2091(.a(s_221), .O(gate165inter4));
  nand2 gate2092(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2093(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2094(.a(G462), .O(gate165inter7));
  inv1  gate2095(.a(G540), .O(gate165inter8));
  nand2 gate2096(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2097(.a(s_221), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2098(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2099(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2100(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1779(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1780(.a(gate167inter0), .b(s_176), .O(gate167inter1));
  and2  gate1781(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1782(.a(s_176), .O(gate167inter3));
  inv1  gate1783(.a(s_177), .O(gate167inter4));
  nand2 gate1784(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1785(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1786(.a(G468), .O(gate167inter7));
  inv1  gate1787(.a(G543), .O(gate167inter8));
  nand2 gate1788(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1789(.a(s_177), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1790(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1791(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1792(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate617(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate618(.a(gate174inter0), .b(s_10), .O(gate174inter1));
  and2  gate619(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate620(.a(s_10), .O(gate174inter3));
  inv1  gate621(.a(s_11), .O(gate174inter4));
  nand2 gate622(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate623(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate624(.a(G489), .O(gate174inter7));
  inv1  gate625(.a(G552), .O(gate174inter8));
  nand2 gate626(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate627(.a(s_11), .b(gate174inter3), .O(gate174inter10));
  nor2  gate628(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate629(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate630(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1569(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1570(.a(gate175inter0), .b(s_146), .O(gate175inter1));
  and2  gate1571(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1572(.a(s_146), .O(gate175inter3));
  inv1  gate1573(.a(s_147), .O(gate175inter4));
  nand2 gate1574(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1575(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1576(.a(G492), .O(gate175inter7));
  inv1  gate1577(.a(G555), .O(gate175inter8));
  nand2 gate1578(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1579(.a(s_147), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1580(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1581(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1582(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1471(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1472(.a(gate177inter0), .b(s_132), .O(gate177inter1));
  and2  gate1473(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1474(.a(s_132), .O(gate177inter3));
  inv1  gate1475(.a(s_133), .O(gate177inter4));
  nand2 gate1476(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1477(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1478(.a(G498), .O(gate177inter7));
  inv1  gate1479(.a(G558), .O(gate177inter8));
  nand2 gate1480(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1481(.a(s_133), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1482(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1483(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1484(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1947(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1948(.a(gate180inter0), .b(s_200), .O(gate180inter1));
  and2  gate1949(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1950(.a(s_200), .O(gate180inter3));
  inv1  gate1951(.a(s_201), .O(gate180inter4));
  nand2 gate1952(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1953(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1954(.a(G507), .O(gate180inter7));
  inv1  gate1955(.a(G561), .O(gate180inter8));
  nand2 gate1956(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1957(.a(s_201), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1958(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1959(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1960(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate939(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate940(.a(gate181inter0), .b(s_56), .O(gate181inter1));
  and2  gate941(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate942(.a(s_56), .O(gate181inter3));
  inv1  gate943(.a(s_57), .O(gate181inter4));
  nand2 gate944(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate945(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate946(.a(G510), .O(gate181inter7));
  inv1  gate947(.a(G564), .O(gate181inter8));
  nand2 gate948(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate949(.a(s_57), .b(gate181inter3), .O(gate181inter10));
  nor2  gate950(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate951(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate952(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1905(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1906(.a(gate185inter0), .b(s_194), .O(gate185inter1));
  and2  gate1907(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1908(.a(s_194), .O(gate185inter3));
  inv1  gate1909(.a(s_195), .O(gate185inter4));
  nand2 gate1910(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1911(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1912(.a(G570), .O(gate185inter7));
  inv1  gate1913(.a(G571), .O(gate185inter8));
  nand2 gate1914(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1915(.a(s_195), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1916(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1917(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1918(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1051(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1052(.a(gate189inter0), .b(s_72), .O(gate189inter1));
  and2  gate1053(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1054(.a(s_72), .O(gate189inter3));
  inv1  gate1055(.a(s_73), .O(gate189inter4));
  nand2 gate1056(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1057(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1058(.a(G578), .O(gate189inter7));
  inv1  gate1059(.a(G579), .O(gate189inter8));
  nand2 gate1060(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1061(.a(s_73), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1062(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1063(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1064(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1331(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1332(.a(gate191inter0), .b(s_112), .O(gate191inter1));
  and2  gate1333(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1334(.a(s_112), .O(gate191inter3));
  inv1  gate1335(.a(s_113), .O(gate191inter4));
  nand2 gate1336(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1337(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1338(.a(G582), .O(gate191inter7));
  inv1  gate1339(.a(G583), .O(gate191inter8));
  nand2 gate1340(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1341(.a(s_113), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1342(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1343(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1344(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1793(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1794(.a(gate194inter0), .b(s_178), .O(gate194inter1));
  and2  gate1795(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1796(.a(s_178), .O(gate194inter3));
  inv1  gate1797(.a(s_179), .O(gate194inter4));
  nand2 gate1798(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1799(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1800(.a(G588), .O(gate194inter7));
  inv1  gate1801(.a(G589), .O(gate194inter8));
  nand2 gate1802(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1803(.a(s_179), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1804(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1805(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1806(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1261(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1262(.a(gate196inter0), .b(s_102), .O(gate196inter1));
  and2  gate1263(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1264(.a(s_102), .O(gate196inter3));
  inv1  gate1265(.a(s_103), .O(gate196inter4));
  nand2 gate1266(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1267(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1268(.a(G592), .O(gate196inter7));
  inv1  gate1269(.a(G593), .O(gate196inter8));
  nand2 gate1270(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1271(.a(s_103), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1272(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1273(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1274(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1485(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1486(.a(gate209inter0), .b(s_134), .O(gate209inter1));
  and2  gate1487(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1488(.a(s_134), .O(gate209inter3));
  inv1  gate1489(.a(s_135), .O(gate209inter4));
  nand2 gate1490(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1491(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1492(.a(G602), .O(gate209inter7));
  inv1  gate1493(.a(G666), .O(gate209inter8));
  nand2 gate1494(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1495(.a(s_135), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1496(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1497(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1498(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate981(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate982(.a(gate212inter0), .b(s_62), .O(gate212inter1));
  and2  gate983(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate984(.a(s_62), .O(gate212inter3));
  inv1  gate985(.a(s_63), .O(gate212inter4));
  nand2 gate986(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate987(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate988(.a(G617), .O(gate212inter7));
  inv1  gate989(.a(G669), .O(gate212inter8));
  nand2 gate990(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate991(.a(s_63), .b(gate212inter3), .O(gate212inter10));
  nor2  gate992(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate993(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate994(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1093(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1094(.a(gate213inter0), .b(s_78), .O(gate213inter1));
  and2  gate1095(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1096(.a(s_78), .O(gate213inter3));
  inv1  gate1097(.a(s_79), .O(gate213inter4));
  nand2 gate1098(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1099(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1100(.a(G602), .O(gate213inter7));
  inv1  gate1101(.a(G672), .O(gate213inter8));
  nand2 gate1102(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1103(.a(s_79), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1104(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1105(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1106(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1401(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1402(.a(gate223inter0), .b(s_122), .O(gate223inter1));
  and2  gate1403(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1404(.a(s_122), .O(gate223inter3));
  inv1  gate1405(.a(s_123), .O(gate223inter4));
  nand2 gate1406(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1407(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1408(.a(G627), .O(gate223inter7));
  inv1  gate1409(.a(G687), .O(gate223inter8));
  nand2 gate1410(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1411(.a(s_123), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1412(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1413(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1414(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate673(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate674(.a(gate225inter0), .b(s_18), .O(gate225inter1));
  and2  gate675(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate676(.a(s_18), .O(gate225inter3));
  inv1  gate677(.a(s_19), .O(gate225inter4));
  nand2 gate678(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate679(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate680(.a(G690), .O(gate225inter7));
  inv1  gate681(.a(G691), .O(gate225inter8));
  nand2 gate682(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate683(.a(s_19), .b(gate225inter3), .O(gate225inter10));
  nor2  gate684(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate685(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate686(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1219(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1220(.a(gate227inter0), .b(s_96), .O(gate227inter1));
  and2  gate1221(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1222(.a(s_96), .O(gate227inter3));
  inv1  gate1223(.a(s_97), .O(gate227inter4));
  nand2 gate1224(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1225(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1226(.a(G694), .O(gate227inter7));
  inv1  gate1227(.a(G695), .O(gate227inter8));
  nand2 gate1228(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1229(.a(s_97), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1230(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1231(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1232(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate645(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate646(.a(gate233inter0), .b(s_14), .O(gate233inter1));
  and2  gate647(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate648(.a(s_14), .O(gate233inter3));
  inv1  gate649(.a(s_15), .O(gate233inter4));
  nand2 gate650(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate651(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate652(.a(G242), .O(gate233inter7));
  inv1  gate653(.a(G718), .O(gate233inter8));
  nand2 gate654(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate655(.a(s_15), .b(gate233inter3), .O(gate233inter10));
  nor2  gate656(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate657(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate658(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1933(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1934(.a(gate234inter0), .b(s_198), .O(gate234inter1));
  and2  gate1935(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1936(.a(s_198), .O(gate234inter3));
  inv1  gate1937(.a(s_199), .O(gate234inter4));
  nand2 gate1938(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1939(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1940(.a(G245), .O(gate234inter7));
  inv1  gate1941(.a(G721), .O(gate234inter8));
  nand2 gate1942(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1943(.a(s_199), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1944(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1945(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1946(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate785(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate786(.a(gate235inter0), .b(s_34), .O(gate235inter1));
  and2  gate787(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate788(.a(s_34), .O(gate235inter3));
  inv1  gate789(.a(s_35), .O(gate235inter4));
  nand2 gate790(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate791(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate792(.a(G248), .O(gate235inter7));
  inv1  gate793(.a(G724), .O(gate235inter8));
  nand2 gate794(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate795(.a(s_35), .b(gate235inter3), .O(gate235inter10));
  nor2  gate796(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate797(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate798(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate813(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate814(.a(gate236inter0), .b(s_38), .O(gate236inter1));
  and2  gate815(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate816(.a(s_38), .O(gate236inter3));
  inv1  gate817(.a(s_39), .O(gate236inter4));
  nand2 gate818(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate819(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate820(.a(G251), .O(gate236inter7));
  inv1  gate821(.a(G727), .O(gate236inter8));
  nand2 gate822(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate823(.a(s_39), .b(gate236inter3), .O(gate236inter10));
  nor2  gate824(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate825(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate826(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1961(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1962(.a(gate242inter0), .b(s_202), .O(gate242inter1));
  and2  gate1963(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1964(.a(s_202), .O(gate242inter3));
  inv1  gate1965(.a(s_203), .O(gate242inter4));
  nand2 gate1966(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1967(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1968(.a(G718), .O(gate242inter7));
  inv1  gate1969(.a(G730), .O(gate242inter8));
  nand2 gate1970(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1971(.a(s_203), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1972(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1973(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1974(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate897(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate898(.a(gate245inter0), .b(s_50), .O(gate245inter1));
  and2  gate899(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate900(.a(s_50), .O(gate245inter3));
  inv1  gate901(.a(s_51), .O(gate245inter4));
  nand2 gate902(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate903(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate904(.a(G248), .O(gate245inter7));
  inv1  gate905(.a(G736), .O(gate245inter8));
  nand2 gate906(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate907(.a(s_51), .b(gate245inter3), .O(gate245inter10));
  nor2  gate908(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate909(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate910(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate953(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate954(.a(gate248inter0), .b(s_58), .O(gate248inter1));
  and2  gate955(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate956(.a(s_58), .O(gate248inter3));
  inv1  gate957(.a(s_59), .O(gate248inter4));
  nand2 gate958(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate959(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate960(.a(G727), .O(gate248inter7));
  inv1  gate961(.a(G739), .O(gate248inter8));
  nand2 gate962(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate963(.a(s_59), .b(gate248inter3), .O(gate248inter10));
  nor2  gate964(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate965(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate966(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1989(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1990(.a(gate258inter0), .b(s_206), .O(gate258inter1));
  and2  gate1991(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1992(.a(s_206), .O(gate258inter3));
  inv1  gate1993(.a(s_207), .O(gate258inter4));
  nand2 gate1994(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1995(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1996(.a(G756), .O(gate258inter7));
  inv1  gate1997(.a(G757), .O(gate258inter8));
  nand2 gate1998(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1999(.a(s_207), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2000(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2001(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2002(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1373(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1374(.a(gate261inter0), .b(s_118), .O(gate261inter1));
  and2  gate1375(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1376(.a(s_118), .O(gate261inter3));
  inv1  gate1377(.a(s_119), .O(gate261inter4));
  nand2 gate1378(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1379(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1380(.a(G762), .O(gate261inter7));
  inv1  gate1381(.a(G763), .O(gate261inter8));
  nand2 gate1382(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1383(.a(s_119), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1384(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1385(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1386(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1247(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1248(.a(gate280inter0), .b(s_100), .O(gate280inter1));
  and2  gate1249(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1250(.a(s_100), .O(gate280inter3));
  inv1  gate1251(.a(s_101), .O(gate280inter4));
  nand2 gate1252(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1253(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1254(.a(G779), .O(gate280inter7));
  inv1  gate1255(.a(G803), .O(gate280inter8));
  nand2 gate1256(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1257(.a(s_101), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1258(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1259(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1260(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1149(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1150(.a(gate285inter0), .b(s_86), .O(gate285inter1));
  and2  gate1151(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1152(.a(s_86), .O(gate285inter3));
  inv1  gate1153(.a(s_87), .O(gate285inter4));
  nand2 gate1154(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1155(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1156(.a(G660), .O(gate285inter7));
  inv1  gate1157(.a(G812), .O(gate285inter8));
  nand2 gate1158(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1159(.a(s_87), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1160(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1161(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1162(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1751(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1752(.a(gate295inter0), .b(s_172), .O(gate295inter1));
  and2  gate1753(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1754(.a(s_172), .O(gate295inter3));
  inv1  gate1755(.a(s_173), .O(gate295inter4));
  nand2 gate1756(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1757(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1758(.a(G830), .O(gate295inter7));
  inv1  gate1759(.a(G831), .O(gate295inter8));
  nand2 gate1760(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1761(.a(s_173), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1762(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1763(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1764(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1177(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1178(.a(gate296inter0), .b(s_90), .O(gate296inter1));
  and2  gate1179(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1180(.a(s_90), .O(gate296inter3));
  inv1  gate1181(.a(s_91), .O(gate296inter4));
  nand2 gate1182(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1183(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1184(.a(G826), .O(gate296inter7));
  inv1  gate1185(.a(G827), .O(gate296inter8));
  nand2 gate1186(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1187(.a(s_91), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1188(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1189(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1190(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate575(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate576(.a(gate392inter0), .b(s_4), .O(gate392inter1));
  and2  gate577(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate578(.a(s_4), .O(gate392inter3));
  inv1  gate579(.a(s_5), .O(gate392inter4));
  nand2 gate580(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate581(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate582(.a(G6), .O(gate392inter7));
  inv1  gate583(.a(G1051), .O(gate392inter8));
  nand2 gate584(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate585(.a(s_5), .b(gate392inter3), .O(gate392inter10));
  nor2  gate586(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate587(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate588(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate659(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate660(.a(gate395inter0), .b(s_16), .O(gate395inter1));
  and2  gate661(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate662(.a(s_16), .O(gate395inter3));
  inv1  gate663(.a(s_17), .O(gate395inter4));
  nand2 gate664(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate665(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate666(.a(G9), .O(gate395inter7));
  inv1  gate667(.a(G1060), .O(gate395inter8));
  nand2 gate668(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate669(.a(s_17), .b(gate395inter3), .O(gate395inter10));
  nor2  gate670(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate671(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate672(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate869(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate870(.a(gate396inter0), .b(s_46), .O(gate396inter1));
  and2  gate871(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate872(.a(s_46), .O(gate396inter3));
  inv1  gate873(.a(s_47), .O(gate396inter4));
  nand2 gate874(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate875(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate876(.a(G10), .O(gate396inter7));
  inv1  gate877(.a(G1063), .O(gate396inter8));
  nand2 gate878(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate879(.a(s_47), .b(gate396inter3), .O(gate396inter10));
  nor2  gate880(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate881(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate882(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1555(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1556(.a(gate397inter0), .b(s_144), .O(gate397inter1));
  and2  gate1557(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1558(.a(s_144), .O(gate397inter3));
  inv1  gate1559(.a(s_145), .O(gate397inter4));
  nand2 gate1560(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1561(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1562(.a(G11), .O(gate397inter7));
  inv1  gate1563(.a(G1066), .O(gate397inter8));
  nand2 gate1564(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1565(.a(s_145), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1566(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1567(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1568(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1835(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1836(.a(gate400inter0), .b(s_184), .O(gate400inter1));
  and2  gate1837(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1838(.a(s_184), .O(gate400inter3));
  inv1  gate1839(.a(s_185), .O(gate400inter4));
  nand2 gate1840(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1841(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1842(.a(G14), .O(gate400inter7));
  inv1  gate1843(.a(G1075), .O(gate400inter8));
  nand2 gate1844(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1845(.a(s_185), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1846(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1847(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1848(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate561(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate562(.a(gate402inter0), .b(s_2), .O(gate402inter1));
  and2  gate563(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate564(.a(s_2), .O(gate402inter3));
  inv1  gate565(.a(s_3), .O(gate402inter4));
  nand2 gate566(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate567(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate568(.a(G16), .O(gate402inter7));
  inv1  gate569(.a(G1081), .O(gate402inter8));
  nand2 gate570(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate571(.a(s_3), .b(gate402inter3), .O(gate402inter10));
  nor2  gate572(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate573(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate574(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1765(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1766(.a(gate403inter0), .b(s_174), .O(gate403inter1));
  and2  gate1767(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1768(.a(s_174), .O(gate403inter3));
  inv1  gate1769(.a(s_175), .O(gate403inter4));
  nand2 gate1770(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1771(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1772(.a(G17), .O(gate403inter7));
  inv1  gate1773(.a(G1084), .O(gate403inter8));
  nand2 gate1774(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1775(.a(s_175), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1776(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1777(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1778(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2059(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2060(.a(gate414inter0), .b(s_216), .O(gate414inter1));
  and2  gate2061(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2062(.a(s_216), .O(gate414inter3));
  inv1  gate2063(.a(s_217), .O(gate414inter4));
  nand2 gate2064(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2065(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2066(.a(G28), .O(gate414inter7));
  inv1  gate2067(.a(G1117), .O(gate414inter8));
  nand2 gate2068(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2069(.a(s_217), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2070(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2071(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2072(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1317(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1318(.a(gate420inter0), .b(s_110), .O(gate420inter1));
  and2  gate1319(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1320(.a(s_110), .O(gate420inter3));
  inv1  gate1321(.a(s_111), .O(gate420inter4));
  nand2 gate1322(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1323(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1324(.a(G1036), .O(gate420inter7));
  inv1  gate1325(.a(G1132), .O(gate420inter8));
  nand2 gate1326(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1327(.a(s_111), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1328(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1329(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1330(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1205(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1206(.a(gate422inter0), .b(s_94), .O(gate422inter1));
  and2  gate1207(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1208(.a(s_94), .O(gate422inter3));
  inv1  gate1209(.a(s_95), .O(gate422inter4));
  nand2 gate1210(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1211(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1212(.a(G1039), .O(gate422inter7));
  inv1  gate1213(.a(G1135), .O(gate422inter8));
  nand2 gate1214(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1215(.a(s_95), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1216(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1217(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1218(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1877(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1878(.a(gate427inter0), .b(s_190), .O(gate427inter1));
  and2  gate1879(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1880(.a(s_190), .O(gate427inter3));
  inv1  gate1881(.a(s_191), .O(gate427inter4));
  nand2 gate1882(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1883(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1884(.a(G5), .O(gate427inter7));
  inv1  gate1885(.a(G1144), .O(gate427inter8));
  nand2 gate1886(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1887(.a(s_191), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1888(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1889(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1890(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1891(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1892(.a(gate429inter0), .b(s_192), .O(gate429inter1));
  and2  gate1893(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1894(.a(s_192), .O(gate429inter3));
  inv1  gate1895(.a(s_193), .O(gate429inter4));
  nand2 gate1896(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1897(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1898(.a(G6), .O(gate429inter7));
  inv1  gate1899(.a(G1147), .O(gate429inter8));
  nand2 gate1900(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1901(.a(s_193), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1902(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1903(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1904(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1415(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1416(.a(gate430inter0), .b(s_124), .O(gate430inter1));
  and2  gate1417(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1418(.a(s_124), .O(gate430inter3));
  inv1  gate1419(.a(s_125), .O(gate430inter4));
  nand2 gate1420(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1421(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1422(.a(G1051), .O(gate430inter7));
  inv1  gate1423(.a(G1147), .O(gate430inter8));
  nand2 gate1424(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1425(.a(s_125), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1426(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1427(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1428(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1289(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1290(.a(gate434inter0), .b(s_106), .O(gate434inter1));
  and2  gate1291(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1292(.a(s_106), .O(gate434inter3));
  inv1  gate1293(.a(s_107), .O(gate434inter4));
  nand2 gate1294(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1295(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1296(.a(G1057), .O(gate434inter7));
  inv1  gate1297(.a(G1153), .O(gate434inter8));
  nand2 gate1298(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1299(.a(s_107), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1300(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1301(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1302(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1275(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1276(.a(gate436inter0), .b(s_104), .O(gate436inter1));
  and2  gate1277(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1278(.a(s_104), .O(gate436inter3));
  inv1  gate1279(.a(s_105), .O(gate436inter4));
  nand2 gate1280(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1281(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1282(.a(G1060), .O(gate436inter7));
  inv1  gate1283(.a(G1156), .O(gate436inter8));
  nand2 gate1284(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1285(.a(s_105), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1286(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1287(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1288(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1597(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1598(.a(gate438inter0), .b(s_150), .O(gate438inter1));
  and2  gate1599(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1600(.a(s_150), .O(gate438inter3));
  inv1  gate1601(.a(s_151), .O(gate438inter4));
  nand2 gate1602(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1603(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1604(.a(G1063), .O(gate438inter7));
  inv1  gate1605(.a(G1159), .O(gate438inter8));
  nand2 gate1606(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1607(.a(s_151), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1608(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1609(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1610(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1443(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1444(.a(gate442inter0), .b(s_128), .O(gate442inter1));
  and2  gate1445(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1446(.a(s_128), .O(gate442inter3));
  inv1  gate1447(.a(s_129), .O(gate442inter4));
  nand2 gate1448(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1449(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1450(.a(G1069), .O(gate442inter7));
  inv1  gate1451(.a(G1165), .O(gate442inter8));
  nand2 gate1452(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1453(.a(s_129), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1454(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1455(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1456(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1499(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1500(.a(gate445inter0), .b(s_136), .O(gate445inter1));
  and2  gate1501(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1502(.a(s_136), .O(gate445inter3));
  inv1  gate1503(.a(s_137), .O(gate445inter4));
  nand2 gate1504(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1505(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1506(.a(G14), .O(gate445inter7));
  inv1  gate1507(.a(G1171), .O(gate445inter8));
  nand2 gate1508(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1509(.a(s_137), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1510(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1511(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1512(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1849(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1850(.a(gate450inter0), .b(s_186), .O(gate450inter1));
  and2  gate1851(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1852(.a(s_186), .O(gate450inter3));
  inv1  gate1853(.a(s_187), .O(gate450inter4));
  nand2 gate1854(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1855(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1856(.a(G1081), .O(gate450inter7));
  inv1  gate1857(.a(G1177), .O(gate450inter8));
  nand2 gate1858(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1859(.a(s_187), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1860(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1861(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1862(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1625(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1626(.a(gate459inter0), .b(s_154), .O(gate459inter1));
  and2  gate1627(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1628(.a(s_154), .O(gate459inter3));
  inv1  gate1629(.a(s_155), .O(gate459inter4));
  nand2 gate1630(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1631(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1632(.a(G21), .O(gate459inter7));
  inv1  gate1633(.a(G1192), .O(gate459inter8));
  nand2 gate1634(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1635(.a(s_155), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1636(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1637(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1638(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1233(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1234(.a(gate466inter0), .b(s_98), .O(gate466inter1));
  and2  gate1235(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1236(.a(s_98), .O(gate466inter3));
  inv1  gate1237(.a(s_99), .O(gate466inter4));
  nand2 gate1238(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1239(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1240(.a(G1105), .O(gate466inter7));
  inv1  gate1241(.a(G1201), .O(gate466inter8));
  nand2 gate1242(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1243(.a(s_99), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1244(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1245(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1246(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1709(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1710(.a(gate467inter0), .b(s_166), .O(gate467inter1));
  and2  gate1711(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1712(.a(s_166), .O(gate467inter3));
  inv1  gate1713(.a(s_167), .O(gate467inter4));
  nand2 gate1714(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1715(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1716(.a(G25), .O(gate467inter7));
  inv1  gate1717(.a(G1204), .O(gate467inter8));
  nand2 gate1718(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1719(.a(s_167), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1720(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1721(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1722(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate771(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate772(.a(gate468inter0), .b(s_32), .O(gate468inter1));
  and2  gate773(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate774(.a(s_32), .O(gate468inter3));
  inv1  gate775(.a(s_33), .O(gate468inter4));
  nand2 gate776(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate777(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate778(.a(G1108), .O(gate468inter7));
  inv1  gate779(.a(G1204), .O(gate468inter8));
  nand2 gate780(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate781(.a(s_33), .b(gate468inter3), .O(gate468inter10));
  nor2  gate782(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate783(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate784(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate743(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate744(.a(gate474inter0), .b(s_28), .O(gate474inter1));
  and2  gate745(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate746(.a(s_28), .O(gate474inter3));
  inv1  gate747(.a(s_29), .O(gate474inter4));
  nand2 gate748(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate749(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate750(.a(G1117), .O(gate474inter7));
  inv1  gate751(.a(G1213), .O(gate474inter8));
  nand2 gate752(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate753(.a(s_29), .b(gate474inter3), .O(gate474inter10));
  nor2  gate754(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate755(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate756(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1807(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1808(.a(gate481inter0), .b(s_180), .O(gate481inter1));
  and2  gate1809(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1810(.a(s_180), .O(gate481inter3));
  inv1  gate1811(.a(s_181), .O(gate481inter4));
  nand2 gate1812(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1813(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1814(.a(G32), .O(gate481inter7));
  inv1  gate1815(.a(G1225), .O(gate481inter8));
  nand2 gate1816(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1817(.a(s_181), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1818(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1819(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1820(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate995(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate996(.a(gate493inter0), .b(s_64), .O(gate493inter1));
  and2  gate997(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate998(.a(s_64), .O(gate493inter3));
  inv1  gate999(.a(s_65), .O(gate493inter4));
  nand2 gate1000(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1001(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1002(.a(G1248), .O(gate493inter7));
  inv1  gate1003(.a(G1249), .O(gate493inter8));
  nand2 gate1004(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1005(.a(s_65), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1006(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1007(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1008(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2045(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2046(.a(gate502inter0), .b(s_214), .O(gate502inter1));
  and2  gate2047(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2048(.a(s_214), .O(gate502inter3));
  inv1  gate2049(.a(s_215), .O(gate502inter4));
  nand2 gate2050(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2051(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2052(.a(G1266), .O(gate502inter7));
  inv1  gate2053(.a(G1267), .O(gate502inter8));
  nand2 gate2054(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2055(.a(s_215), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2056(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2057(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2058(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1863(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1864(.a(gate508inter0), .b(s_188), .O(gate508inter1));
  and2  gate1865(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1866(.a(s_188), .O(gate508inter3));
  inv1  gate1867(.a(s_189), .O(gate508inter4));
  nand2 gate1868(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1869(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1870(.a(G1278), .O(gate508inter7));
  inv1  gate1871(.a(G1279), .O(gate508inter8));
  nand2 gate1872(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1873(.a(s_189), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1874(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1875(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1876(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1583(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1584(.a(gate509inter0), .b(s_148), .O(gate509inter1));
  and2  gate1585(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1586(.a(s_148), .O(gate509inter3));
  inv1  gate1587(.a(s_149), .O(gate509inter4));
  nand2 gate1588(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1589(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1590(.a(G1280), .O(gate509inter7));
  inv1  gate1591(.a(G1281), .O(gate509inter8));
  nand2 gate1592(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1593(.a(s_149), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1594(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1595(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1596(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule