module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1443(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1444(.a(gate14inter0), .b(s_128), .O(gate14inter1));
  and2  gate1445(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1446(.a(s_128), .O(gate14inter3));
  inv1  gate1447(.a(s_129), .O(gate14inter4));
  nand2 gate1448(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1449(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1450(.a(G11), .O(gate14inter7));
  inv1  gate1451(.a(G12), .O(gate14inter8));
  nand2 gate1452(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1453(.a(s_129), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1454(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1455(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1456(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate757(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate758(.a(gate15inter0), .b(s_30), .O(gate15inter1));
  and2  gate759(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate760(.a(s_30), .O(gate15inter3));
  inv1  gate761(.a(s_31), .O(gate15inter4));
  nand2 gate762(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate763(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate764(.a(G13), .O(gate15inter7));
  inv1  gate765(.a(G14), .O(gate15inter8));
  nand2 gate766(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate767(.a(s_31), .b(gate15inter3), .O(gate15inter10));
  nor2  gate768(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate769(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate770(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate967(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate968(.a(gate17inter0), .b(s_60), .O(gate17inter1));
  and2  gate969(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate970(.a(s_60), .O(gate17inter3));
  inv1  gate971(.a(s_61), .O(gate17inter4));
  nand2 gate972(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate973(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate974(.a(G17), .O(gate17inter7));
  inv1  gate975(.a(G18), .O(gate17inter8));
  nand2 gate976(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate977(.a(s_61), .b(gate17inter3), .O(gate17inter10));
  nor2  gate978(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate979(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate980(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1093(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1094(.a(gate18inter0), .b(s_78), .O(gate18inter1));
  and2  gate1095(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1096(.a(s_78), .O(gate18inter3));
  inv1  gate1097(.a(s_79), .O(gate18inter4));
  nand2 gate1098(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1099(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1100(.a(G19), .O(gate18inter7));
  inv1  gate1101(.a(G20), .O(gate18inter8));
  nand2 gate1102(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1103(.a(s_79), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1104(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1105(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1106(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1471(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1472(.a(gate19inter0), .b(s_132), .O(gate19inter1));
  and2  gate1473(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1474(.a(s_132), .O(gate19inter3));
  inv1  gate1475(.a(s_133), .O(gate19inter4));
  nand2 gate1476(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1477(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1478(.a(G21), .O(gate19inter7));
  inv1  gate1479(.a(G22), .O(gate19inter8));
  nand2 gate1480(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1481(.a(s_133), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1482(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1483(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1484(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2241(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2242(.a(gate20inter0), .b(s_242), .O(gate20inter1));
  and2  gate2243(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2244(.a(s_242), .O(gate20inter3));
  inv1  gate2245(.a(s_243), .O(gate20inter4));
  nand2 gate2246(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2247(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2248(.a(G23), .O(gate20inter7));
  inv1  gate2249(.a(G24), .O(gate20inter8));
  nand2 gate2250(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2251(.a(s_243), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2252(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2253(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2254(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2395(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2396(.a(gate24inter0), .b(s_264), .O(gate24inter1));
  and2  gate2397(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2398(.a(s_264), .O(gate24inter3));
  inv1  gate2399(.a(s_265), .O(gate24inter4));
  nand2 gate2400(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2401(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2402(.a(G31), .O(gate24inter7));
  inv1  gate2403(.a(G32), .O(gate24inter8));
  nand2 gate2404(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2405(.a(s_265), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2406(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2407(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2408(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate2465(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2466(.a(gate25inter0), .b(s_274), .O(gate25inter1));
  and2  gate2467(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2468(.a(s_274), .O(gate25inter3));
  inv1  gate2469(.a(s_275), .O(gate25inter4));
  nand2 gate2470(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2471(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2472(.a(G1), .O(gate25inter7));
  inv1  gate2473(.a(G5), .O(gate25inter8));
  nand2 gate2474(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2475(.a(s_275), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2476(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2477(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2478(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1975(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1976(.a(gate27inter0), .b(s_204), .O(gate27inter1));
  and2  gate1977(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1978(.a(s_204), .O(gate27inter3));
  inv1  gate1979(.a(s_205), .O(gate27inter4));
  nand2 gate1980(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1981(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1982(.a(G2), .O(gate27inter7));
  inv1  gate1983(.a(G6), .O(gate27inter8));
  nand2 gate1984(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1985(.a(s_205), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1986(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1987(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1988(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate2423(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2424(.a(gate28inter0), .b(s_268), .O(gate28inter1));
  and2  gate2425(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2426(.a(s_268), .O(gate28inter3));
  inv1  gate2427(.a(s_269), .O(gate28inter4));
  nand2 gate2428(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2429(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2430(.a(G10), .O(gate28inter7));
  inv1  gate2431(.a(G14), .O(gate28inter8));
  nand2 gate2432(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2433(.a(s_269), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2434(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2435(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2436(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate701(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate702(.a(gate29inter0), .b(s_22), .O(gate29inter1));
  and2  gate703(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate704(.a(s_22), .O(gate29inter3));
  inv1  gate705(.a(s_23), .O(gate29inter4));
  nand2 gate706(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate707(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate708(.a(G3), .O(gate29inter7));
  inv1  gate709(.a(G7), .O(gate29inter8));
  nand2 gate710(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate711(.a(s_23), .b(gate29inter3), .O(gate29inter10));
  nor2  gate712(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate713(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate714(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1401(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1402(.a(gate30inter0), .b(s_122), .O(gate30inter1));
  and2  gate1403(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1404(.a(s_122), .O(gate30inter3));
  inv1  gate1405(.a(s_123), .O(gate30inter4));
  nand2 gate1406(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1407(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1408(.a(G11), .O(gate30inter7));
  inv1  gate1409(.a(G15), .O(gate30inter8));
  nand2 gate1410(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1411(.a(s_123), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1412(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1413(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1414(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1793(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1794(.a(gate33inter0), .b(s_178), .O(gate33inter1));
  and2  gate1795(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1796(.a(s_178), .O(gate33inter3));
  inv1  gate1797(.a(s_179), .O(gate33inter4));
  nand2 gate1798(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1799(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1800(.a(G17), .O(gate33inter7));
  inv1  gate1801(.a(G21), .O(gate33inter8));
  nand2 gate1802(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1803(.a(s_179), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1804(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1805(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1806(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1751(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1752(.a(gate34inter0), .b(s_172), .O(gate34inter1));
  and2  gate1753(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1754(.a(s_172), .O(gate34inter3));
  inv1  gate1755(.a(s_173), .O(gate34inter4));
  nand2 gate1756(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1757(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1758(.a(G25), .O(gate34inter7));
  inv1  gate1759(.a(G29), .O(gate34inter8));
  nand2 gate1760(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1761(.a(s_173), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1762(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1763(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1764(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2745(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2746(.a(gate38inter0), .b(s_314), .O(gate38inter1));
  and2  gate2747(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2748(.a(s_314), .O(gate38inter3));
  inv1  gate2749(.a(s_315), .O(gate38inter4));
  nand2 gate2750(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2751(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2752(.a(G27), .O(gate38inter7));
  inv1  gate2753(.a(G31), .O(gate38inter8));
  nand2 gate2754(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2755(.a(s_315), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2756(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2757(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2758(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2311(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2312(.a(gate41inter0), .b(s_252), .O(gate41inter1));
  and2  gate2313(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2314(.a(s_252), .O(gate41inter3));
  inv1  gate2315(.a(s_253), .O(gate41inter4));
  nand2 gate2316(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2317(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2318(.a(G1), .O(gate41inter7));
  inv1  gate2319(.a(G266), .O(gate41inter8));
  nand2 gate2320(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2321(.a(s_253), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2322(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2323(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2324(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2913(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2914(.a(gate42inter0), .b(s_338), .O(gate42inter1));
  and2  gate2915(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2916(.a(s_338), .O(gate42inter3));
  inv1  gate2917(.a(s_339), .O(gate42inter4));
  nand2 gate2918(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2919(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2920(.a(G2), .O(gate42inter7));
  inv1  gate2921(.a(G266), .O(gate42inter8));
  nand2 gate2922(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2923(.a(s_339), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2924(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2925(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2926(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2017(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2018(.a(gate44inter0), .b(s_210), .O(gate44inter1));
  and2  gate2019(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2020(.a(s_210), .O(gate44inter3));
  inv1  gate2021(.a(s_211), .O(gate44inter4));
  nand2 gate2022(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2023(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2024(.a(G4), .O(gate44inter7));
  inv1  gate2025(.a(G269), .O(gate44inter8));
  nand2 gate2026(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2027(.a(s_211), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2028(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2029(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2030(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate911(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate912(.a(gate48inter0), .b(s_52), .O(gate48inter1));
  and2  gate913(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate914(.a(s_52), .O(gate48inter3));
  inv1  gate915(.a(s_53), .O(gate48inter4));
  nand2 gate916(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate917(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate918(.a(G8), .O(gate48inter7));
  inv1  gate919(.a(G275), .O(gate48inter8));
  nand2 gate920(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate921(.a(s_53), .b(gate48inter3), .O(gate48inter10));
  nor2  gate922(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate923(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate924(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2199(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2200(.a(gate49inter0), .b(s_236), .O(gate49inter1));
  and2  gate2201(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2202(.a(s_236), .O(gate49inter3));
  inv1  gate2203(.a(s_237), .O(gate49inter4));
  nand2 gate2204(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2205(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2206(.a(G9), .O(gate49inter7));
  inv1  gate2207(.a(G278), .O(gate49inter8));
  nand2 gate2208(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2209(.a(s_237), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2210(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2211(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2212(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1135(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1136(.a(gate50inter0), .b(s_84), .O(gate50inter1));
  and2  gate1137(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1138(.a(s_84), .O(gate50inter3));
  inv1  gate1139(.a(s_85), .O(gate50inter4));
  nand2 gate1140(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1141(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1142(.a(G10), .O(gate50inter7));
  inv1  gate1143(.a(G278), .O(gate50inter8));
  nand2 gate1144(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1145(.a(s_85), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1146(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1147(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1148(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1219(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1220(.a(gate54inter0), .b(s_96), .O(gate54inter1));
  and2  gate1221(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1222(.a(s_96), .O(gate54inter3));
  inv1  gate1223(.a(s_97), .O(gate54inter4));
  nand2 gate1224(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1225(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1226(.a(G14), .O(gate54inter7));
  inv1  gate1227(.a(G284), .O(gate54inter8));
  nand2 gate1228(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1229(.a(s_97), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1230(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1231(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1232(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate2941(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2942(.a(gate55inter0), .b(s_342), .O(gate55inter1));
  and2  gate2943(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2944(.a(s_342), .O(gate55inter3));
  inv1  gate2945(.a(s_343), .O(gate55inter4));
  nand2 gate2946(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2947(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2948(.a(G15), .O(gate55inter7));
  inv1  gate2949(.a(G287), .O(gate55inter8));
  nand2 gate2950(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2951(.a(s_343), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2952(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2953(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2954(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2507(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2508(.a(gate56inter0), .b(s_280), .O(gate56inter1));
  and2  gate2509(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2510(.a(s_280), .O(gate56inter3));
  inv1  gate2511(.a(s_281), .O(gate56inter4));
  nand2 gate2512(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2513(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2514(.a(G16), .O(gate56inter7));
  inv1  gate2515(.a(G287), .O(gate56inter8));
  nand2 gate2516(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2517(.a(s_281), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2518(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2519(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2520(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1457(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1458(.a(gate60inter0), .b(s_130), .O(gate60inter1));
  and2  gate1459(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1460(.a(s_130), .O(gate60inter3));
  inv1  gate1461(.a(s_131), .O(gate60inter4));
  nand2 gate1462(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1463(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1464(.a(G20), .O(gate60inter7));
  inv1  gate1465(.a(G293), .O(gate60inter8));
  nand2 gate1466(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1467(.a(s_131), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1468(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1469(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1470(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate2983(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2984(.a(gate63inter0), .b(s_348), .O(gate63inter1));
  and2  gate2985(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2986(.a(s_348), .O(gate63inter3));
  inv1  gate2987(.a(s_349), .O(gate63inter4));
  nand2 gate2988(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2989(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2990(.a(G23), .O(gate63inter7));
  inv1  gate2991(.a(G299), .O(gate63inter8));
  nand2 gate2992(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2993(.a(s_349), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2994(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2995(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2996(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2857(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2858(.a(gate67inter0), .b(s_330), .O(gate67inter1));
  and2  gate2859(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2860(.a(s_330), .O(gate67inter3));
  inv1  gate2861(.a(s_331), .O(gate67inter4));
  nand2 gate2862(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2863(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2864(.a(G27), .O(gate67inter7));
  inv1  gate2865(.a(G305), .O(gate67inter8));
  nand2 gate2866(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2867(.a(s_331), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2868(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2869(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2870(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2633(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2634(.a(gate69inter0), .b(s_298), .O(gate69inter1));
  and2  gate2635(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2636(.a(s_298), .O(gate69inter3));
  inv1  gate2637(.a(s_299), .O(gate69inter4));
  nand2 gate2638(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2639(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2640(.a(G29), .O(gate69inter7));
  inv1  gate2641(.a(G308), .O(gate69inter8));
  nand2 gate2642(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2643(.a(s_299), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2644(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2645(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2646(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1821(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1822(.a(gate70inter0), .b(s_182), .O(gate70inter1));
  and2  gate1823(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1824(.a(s_182), .O(gate70inter3));
  inv1  gate1825(.a(s_183), .O(gate70inter4));
  nand2 gate1826(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1827(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1828(.a(G30), .O(gate70inter7));
  inv1  gate1829(.a(G308), .O(gate70inter8));
  nand2 gate1830(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1831(.a(s_183), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1832(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1833(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1834(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1737(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1738(.a(gate73inter0), .b(s_170), .O(gate73inter1));
  and2  gate1739(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1740(.a(s_170), .O(gate73inter3));
  inv1  gate1741(.a(s_171), .O(gate73inter4));
  nand2 gate1742(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1743(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1744(.a(G1), .O(gate73inter7));
  inv1  gate1745(.a(G314), .O(gate73inter8));
  nand2 gate1746(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1747(.a(s_171), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1748(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1749(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1750(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate883(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate884(.a(gate77inter0), .b(s_48), .O(gate77inter1));
  and2  gate885(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate886(.a(s_48), .O(gate77inter3));
  inv1  gate887(.a(s_49), .O(gate77inter4));
  nand2 gate888(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate889(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate890(.a(G2), .O(gate77inter7));
  inv1  gate891(.a(G320), .O(gate77inter8));
  nand2 gate892(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate893(.a(s_49), .b(gate77inter3), .O(gate77inter10));
  nor2  gate894(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate895(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate896(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1653(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1654(.a(gate78inter0), .b(s_158), .O(gate78inter1));
  and2  gate1655(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1656(.a(s_158), .O(gate78inter3));
  inv1  gate1657(.a(s_159), .O(gate78inter4));
  nand2 gate1658(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1659(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1660(.a(G6), .O(gate78inter7));
  inv1  gate1661(.a(G320), .O(gate78inter8));
  nand2 gate1662(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1663(.a(s_159), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1664(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1665(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1666(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2521(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2522(.a(gate79inter0), .b(s_282), .O(gate79inter1));
  and2  gate2523(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2524(.a(s_282), .O(gate79inter3));
  inv1  gate2525(.a(s_283), .O(gate79inter4));
  nand2 gate2526(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2527(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2528(.a(G10), .O(gate79inter7));
  inv1  gate2529(.a(G323), .O(gate79inter8));
  nand2 gate2530(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2531(.a(s_283), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2532(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2533(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2534(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1289(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1290(.a(gate80inter0), .b(s_106), .O(gate80inter1));
  and2  gate1291(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1292(.a(s_106), .O(gate80inter3));
  inv1  gate1293(.a(s_107), .O(gate80inter4));
  nand2 gate1294(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1295(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1296(.a(G14), .O(gate80inter7));
  inv1  gate1297(.a(G323), .O(gate80inter8));
  nand2 gate1298(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1299(.a(s_107), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1300(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1301(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1302(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1527(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1528(.a(gate84inter0), .b(s_140), .O(gate84inter1));
  and2  gate1529(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1530(.a(s_140), .O(gate84inter3));
  inv1  gate1531(.a(s_141), .O(gate84inter4));
  nand2 gate1532(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1533(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1534(.a(G15), .O(gate84inter7));
  inv1  gate1535(.a(G329), .O(gate84inter8));
  nand2 gate1536(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1537(.a(s_141), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1538(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1539(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1540(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate981(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate982(.a(gate85inter0), .b(s_62), .O(gate85inter1));
  and2  gate983(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate984(.a(s_62), .O(gate85inter3));
  inv1  gate985(.a(s_63), .O(gate85inter4));
  nand2 gate986(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate987(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate988(.a(G4), .O(gate85inter7));
  inv1  gate989(.a(G332), .O(gate85inter8));
  nand2 gate990(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate991(.a(s_63), .b(gate85inter3), .O(gate85inter10));
  nor2  gate992(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate993(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate994(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2759(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2760(.a(gate87inter0), .b(s_316), .O(gate87inter1));
  and2  gate2761(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2762(.a(s_316), .O(gate87inter3));
  inv1  gate2763(.a(s_317), .O(gate87inter4));
  nand2 gate2764(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2765(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2766(.a(G12), .O(gate87inter7));
  inv1  gate2767(.a(G335), .O(gate87inter8));
  nand2 gate2768(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2769(.a(s_317), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2770(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2771(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2772(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate2059(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2060(.a(gate88inter0), .b(s_216), .O(gate88inter1));
  and2  gate2061(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2062(.a(s_216), .O(gate88inter3));
  inv1  gate2063(.a(s_217), .O(gate88inter4));
  nand2 gate2064(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2065(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2066(.a(G16), .O(gate88inter7));
  inv1  gate2067(.a(G335), .O(gate88inter8));
  nand2 gate2068(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2069(.a(s_217), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2070(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2071(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2072(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2619(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2620(.a(gate90inter0), .b(s_296), .O(gate90inter1));
  and2  gate2621(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2622(.a(s_296), .O(gate90inter3));
  inv1  gate2623(.a(s_297), .O(gate90inter4));
  nand2 gate2624(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2625(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2626(.a(G21), .O(gate90inter7));
  inv1  gate2627(.a(G338), .O(gate90inter8));
  nand2 gate2628(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2629(.a(s_297), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2630(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2631(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2632(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2185(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2186(.a(gate91inter0), .b(s_234), .O(gate91inter1));
  and2  gate2187(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2188(.a(s_234), .O(gate91inter3));
  inv1  gate2189(.a(s_235), .O(gate91inter4));
  nand2 gate2190(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2191(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2192(.a(G25), .O(gate91inter7));
  inv1  gate2193(.a(G341), .O(gate91inter8));
  nand2 gate2194(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2195(.a(s_235), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2196(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2197(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2198(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1079(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1080(.a(gate94inter0), .b(s_76), .O(gate94inter1));
  and2  gate1081(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1082(.a(s_76), .O(gate94inter3));
  inv1  gate1083(.a(s_77), .O(gate94inter4));
  nand2 gate1084(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1085(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1086(.a(G22), .O(gate94inter7));
  inv1  gate1087(.a(G344), .O(gate94inter8));
  nand2 gate1088(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1089(.a(s_77), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1090(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1091(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1092(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2787(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2788(.a(gate96inter0), .b(s_320), .O(gate96inter1));
  and2  gate2789(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2790(.a(s_320), .O(gate96inter3));
  inv1  gate2791(.a(s_321), .O(gate96inter4));
  nand2 gate2792(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2793(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2794(.a(G30), .O(gate96inter7));
  inv1  gate2795(.a(G347), .O(gate96inter8));
  nand2 gate2796(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2797(.a(s_321), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2798(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2799(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2800(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2997(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2998(.a(gate97inter0), .b(s_350), .O(gate97inter1));
  and2  gate2999(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate3000(.a(s_350), .O(gate97inter3));
  inv1  gate3001(.a(s_351), .O(gate97inter4));
  nand2 gate3002(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate3003(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate3004(.a(G19), .O(gate97inter7));
  inv1  gate3005(.a(G350), .O(gate97inter8));
  nand2 gate3006(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate3007(.a(s_351), .b(gate97inter3), .O(gate97inter10));
  nor2  gate3008(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate3009(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate3010(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate645(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate646(.a(gate98inter0), .b(s_14), .O(gate98inter1));
  and2  gate647(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate648(.a(s_14), .O(gate98inter3));
  inv1  gate649(.a(s_15), .O(gate98inter4));
  nand2 gate650(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate651(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate652(.a(G23), .O(gate98inter7));
  inv1  gate653(.a(G350), .O(gate98inter8));
  nand2 gate654(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate655(.a(s_15), .b(gate98inter3), .O(gate98inter10));
  nor2  gate656(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate657(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate658(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate575(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate576(.a(gate100inter0), .b(s_4), .O(gate100inter1));
  and2  gate577(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate578(.a(s_4), .O(gate100inter3));
  inv1  gate579(.a(s_5), .O(gate100inter4));
  nand2 gate580(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate581(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate582(.a(G31), .O(gate100inter7));
  inv1  gate583(.a(G353), .O(gate100inter8));
  nand2 gate584(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate585(.a(s_5), .b(gate100inter3), .O(gate100inter10));
  nor2  gate586(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate587(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate588(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1891(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1892(.a(gate102inter0), .b(s_192), .O(gate102inter1));
  and2  gate1893(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1894(.a(s_192), .O(gate102inter3));
  inv1  gate1895(.a(s_193), .O(gate102inter4));
  nand2 gate1896(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1897(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1898(.a(G24), .O(gate102inter7));
  inv1  gate1899(.a(G356), .O(gate102inter8));
  nand2 gate1900(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1901(.a(s_193), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1902(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1903(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1904(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1695(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1696(.a(gate103inter0), .b(s_164), .O(gate103inter1));
  and2  gate1697(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1698(.a(s_164), .O(gate103inter3));
  inv1  gate1699(.a(s_165), .O(gate103inter4));
  nand2 gate1700(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1701(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1702(.a(G28), .O(gate103inter7));
  inv1  gate1703(.a(G359), .O(gate103inter8));
  nand2 gate1704(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1705(.a(s_165), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1706(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1707(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1708(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1849(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1850(.a(gate104inter0), .b(s_186), .O(gate104inter1));
  and2  gate1851(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1852(.a(s_186), .O(gate104inter3));
  inv1  gate1853(.a(s_187), .O(gate104inter4));
  nand2 gate1854(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1855(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1856(.a(G32), .O(gate104inter7));
  inv1  gate1857(.a(G359), .O(gate104inter8));
  nand2 gate1858(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1859(.a(s_187), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1860(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1861(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1862(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1807(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1808(.a(gate107inter0), .b(s_180), .O(gate107inter1));
  and2  gate1809(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1810(.a(s_180), .O(gate107inter3));
  inv1  gate1811(.a(s_181), .O(gate107inter4));
  nand2 gate1812(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1813(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1814(.a(G366), .O(gate107inter7));
  inv1  gate1815(.a(G367), .O(gate107inter8));
  nand2 gate1816(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1817(.a(s_181), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1818(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1819(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1820(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2773(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2774(.a(gate110inter0), .b(s_318), .O(gate110inter1));
  and2  gate2775(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2776(.a(s_318), .O(gate110inter3));
  inv1  gate2777(.a(s_319), .O(gate110inter4));
  nand2 gate2778(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2779(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2780(.a(G372), .O(gate110inter7));
  inv1  gate2781(.a(G373), .O(gate110inter8));
  nand2 gate2782(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2783(.a(s_319), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2784(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2785(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2786(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1247(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1248(.a(gate113inter0), .b(s_100), .O(gate113inter1));
  and2  gate1249(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1250(.a(s_100), .O(gate113inter3));
  inv1  gate1251(.a(s_101), .O(gate113inter4));
  nand2 gate1252(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1253(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1254(.a(G378), .O(gate113inter7));
  inv1  gate1255(.a(G379), .O(gate113inter8));
  nand2 gate1256(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1257(.a(s_101), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1258(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1259(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1260(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2493(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2494(.a(gate116inter0), .b(s_278), .O(gate116inter1));
  and2  gate2495(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2496(.a(s_278), .O(gate116inter3));
  inv1  gate2497(.a(s_279), .O(gate116inter4));
  nand2 gate2498(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2499(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2500(.a(G384), .O(gate116inter7));
  inv1  gate2501(.a(G385), .O(gate116inter8));
  nand2 gate2502(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2503(.a(s_279), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2504(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2505(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2506(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate897(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate898(.a(gate118inter0), .b(s_50), .O(gate118inter1));
  and2  gate899(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate900(.a(s_50), .O(gate118inter3));
  inv1  gate901(.a(s_51), .O(gate118inter4));
  nand2 gate902(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate903(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate904(.a(G388), .O(gate118inter7));
  inv1  gate905(.a(G389), .O(gate118inter8));
  nand2 gate906(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate907(.a(s_51), .b(gate118inter3), .O(gate118inter10));
  nor2  gate908(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate909(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate910(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2955(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2956(.a(gate119inter0), .b(s_344), .O(gate119inter1));
  and2  gate2957(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2958(.a(s_344), .O(gate119inter3));
  inv1  gate2959(.a(s_345), .O(gate119inter4));
  nand2 gate2960(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2961(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2962(.a(G390), .O(gate119inter7));
  inv1  gate2963(.a(G391), .O(gate119inter8));
  nand2 gate2964(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2965(.a(s_345), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2966(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2967(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2968(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2801(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2802(.a(gate123inter0), .b(s_322), .O(gate123inter1));
  and2  gate2803(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2804(.a(s_322), .O(gate123inter3));
  inv1  gate2805(.a(s_323), .O(gate123inter4));
  nand2 gate2806(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2807(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2808(.a(G398), .O(gate123inter7));
  inv1  gate2809(.a(G399), .O(gate123inter8));
  nand2 gate2810(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2811(.a(s_323), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2812(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2813(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2814(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2899(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2900(.a(gate125inter0), .b(s_336), .O(gate125inter1));
  and2  gate2901(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2902(.a(s_336), .O(gate125inter3));
  inv1  gate2903(.a(s_337), .O(gate125inter4));
  nand2 gate2904(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2905(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2906(.a(G402), .O(gate125inter7));
  inv1  gate2907(.a(G403), .O(gate125inter8));
  nand2 gate2908(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2909(.a(s_337), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2910(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2911(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2912(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1275(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1276(.a(gate131inter0), .b(s_104), .O(gate131inter1));
  and2  gate1277(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1278(.a(s_104), .O(gate131inter3));
  inv1  gate1279(.a(s_105), .O(gate131inter4));
  nand2 gate1280(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1281(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1282(.a(G414), .O(gate131inter7));
  inv1  gate1283(.a(G415), .O(gate131inter8));
  nand2 gate1284(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1285(.a(s_105), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1286(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1287(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1288(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate785(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate786(.a(gate132inter0), .b(s_34), .O(gate132inter1));
  and2  gate787(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate788(.a(s_34), .O(gate132inter3));
  inv1  gate789(.a(s_35), .O(gate132inter4));
  nand2 gate790(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate791(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate792(.a(G416), .O(gate132inter7));
  inv1  gate793(.a(G417), .O(gate132inter8));
  nand2 gate794(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate795(.a(s_35), .b(gate132inter3), .O(gate132inter10));
  nor2  gate796(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate797(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate798(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2255(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2256(.a(gate133inter0), .b(s_244), .O(gate133inter1));
  and2  gate2257(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2258(.a(s_244), .O(gate133inter3));
  inv1  gate2259(.a(s_245), .O(gate133inter4));
  nand2 gate2260(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2261(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2262(.a(G418), .O(gate133inter7));
  inv1  gate2263(.a(G419), .O(gate133inter8));
  nand2 gate2264(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2265(.a(s_245), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2266(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2267(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2268(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1051(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1052(.a(gate136inter0), .b(s_72), .O(gate136inter1));
  and2  gate1053(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1054(.a(s_72), .O(gate136inter3));
  inv1  gate1055(.a(s_73), .O(gate136inter4));
  nand2 gate1056(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1057(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1058(.a(G424), .O(gate136inter7));
  inv1  gate1059(.a(G425), .O(gate136inter8));
  nand2 gate1060(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1061(.a(s_73), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1062(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1063(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1064(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1345(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1346(.a(gate137inter0), .b(s_114), .O(gate137inter1));
  and2  gate1347(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1348(.a(s_114), .O(gate137inter3));
  inv1  gate1349(.a(s_115), .O(gate137inter4));
  nand2 gate1350(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1351(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1352(.a(G426), .O(gate137inter7));
  inv1  gate1353(.a(G429), .O(gate137inter8));
  nand2 gate1354(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1355(.a(s_115), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1356(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1357(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1358(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1485(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1486(.a(gate138inter0), .b(s_134), .O(gate138inter1));
  and2  gate1487(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1488(.a(s_134), .O(gate138inter3));
  inv1  gate1489(.a(s_135), .O(gate138inter4));
  nand2 gate1490(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1491(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1492(.a(G432), .O(gate138inter7));
  inv1  gate1493(.a(G435), .O(gate138inter8));
  nand2 gate1494(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1495(.a(s_135), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1496(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1497(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1498(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2367(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2368(.a(gate141inter0), .b(s_260), .O(gate141inter1));
  and2  gate2369(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2370(.a(s_260), .O(gate141inter3));
  inv1  gate2371(.a(s_261), .O(gate141inter4));
  nand2 gate2372(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2373(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2374(.a(G450), .O(gate141inter7));
  inv1  gate2375(.a(G453), .O(gate141inter8));
  nand2 gate2376(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2377(.a(s_261), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2378(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2379(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2380(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate2563(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2564(.a(gate145inter0), .b(s_288), .O(gate145inter1));
  and2  gate2565(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2566(.a(s_288), .O(gate145inter3));
  inv1  gate2567(.a(s_289), .O(gate145inter4));
  nand2 gate2568(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2569(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2570(.a(G474), .O(gate145inter7));
  inv1  gate2571(.a(G477), .O(gate145inter8));
  nand2 gate2572(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2573(.a(s_289), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2574(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2575(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2576(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1359(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1360(.a(gate146inter0), .b(s_116), .O(gate146inter1));
  and2  gate1361(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1362(.a(s_116), .O(gate146inter3));
  inv1  gate1363(.a(s_117), .O(gate146inter4));
  nand2 gate1364(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1365(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1366(.a(G480), .O(gate146inter7));
  inv1  gate1367(.a(G483), .O(gate146inter8));
  nand2 gate1368(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1369(.a(s_117), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1370(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1371(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1372(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2213(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2214(.a(gate147inter0), .b(s_238), .O(gate147inter1));
  and2  gate2215(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2216(.a(s_238), .O(gate147inter3));
  inv1  gate2217(.a(s_239), .O(gate147inter4));
  nand2 gate2218(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2219(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2220(.a(G486), .O(gate147inter7));
  inv1  gate2221(.a(G489), .O(gate147inter8));
  nand2 gate2222(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2223(.a(s_239), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2224(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2225(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2226(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate2073(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2074(.a(gate148inter0), .b(s_218), .O(gate148inter1));
  and2  gate2075(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2076(.a(s_218), .O(gate148inter3));
  inv1  gate2077(.a(s_219), .O(gate148inter4));
  nand2 gate2078(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2079(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2080(.a(G492), .O(gate148inter7));
  inv1  gate2081(.a(G495), .O(gate148inter8));
  nand2 gate2082(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2083(.a(s_219), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2084(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2085(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2086(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1065(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1066(.a(gate151inter0), .b(s_74), .O(gate151inter1));
  and2  gate1067(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1068(.a(s_74), .O(gate151inter3));
  inv1  gate1069(.a(s_75), .O(gate151inter4));
  nand2 gate1070(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1071(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1072(.a(G510), .O(gate151inter7));
  inv1  gate1073(.a(G513), .O(gate151inter8));
  nand2 gate1074(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1075(.a(s_75), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1076(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1077(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1078(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1429(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1430(.a(gate156inter0), .b(s_126), .O(gate156inter1));
  and2  gate1431(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1432(.a(s_126), .O(gate156inter3));
  inv1  gate1433(.a(s_127), .O(gate156inter4));
  nand2 gate1434(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1435(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1436(.a(G435), .O(gate156inter7));
  inv1  gate1437(.a(G525), .O(gate156inter8));
  nand2 gate1438(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1439(.a(s_127), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1440(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1441(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1442(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate743(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate744(.a(gate157inter0), .b(s_28), .O(gate157inter1));
  and2  gate745(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate746(.a(s_28), .O(gate157inter3));
  inv1  gate747(.a(s_29), .O(gate157inter4));
  nand2 gate748(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate749(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate750(.a(G438), .O(gate157inter7));
  inv1  gate751(.a(G528), .O(gate157inter8));
  nand2 gate752(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate753(.a(s_29), .b(gate157inter3), .O(gate157inter10));
  nor2  gate754(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate755(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate756(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1541(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1542(.a(gate159inter0), .b(s_142), .O(gate159inter1));
  and2  gate1543(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1544(.a(s_142), .O(gate159inter3));
  inv1  gate1545(.a(s_143), .O(gate159inter4));
  nand2 gate1546(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1547(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1548(.a(G444), .O(gate159inter7));
  inv1  gate1549(.a(G531), .O(gate159inter8));
  nand2 gate1550(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1551(.a(s_143), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1552(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1553(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1554(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2689(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2690(.a(gate160inter0), .b(s_306), .O(gate160inter1));
  and2  gate2691(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2692(.a(s_306), .O(gate160inter3));
  inv1  gate2693(.a(s_307), .O(gate160inter4));
  nand2 gate2694(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2695(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2696(.a(G447), .O(gate160inter7));
  inv1  gate2697(.a(G531), .O(gate160inter8));
  nand2 gate2698(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2699(.a(s_307), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2700(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2701(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2702(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1835(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1836(.a(gate167inter0), .b(s_184), .O(gate167inter1));
  and2  gate1837(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1838(.a(s_184), .O(gate167inter3));
  inv1  gate1839(.a(s_185), .O(gate167inter4));
  nand2 gate1840(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1841(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1842(.a(G468), .O(gate167inter7));
  inv1  gate1843(.a(G543), .O(gate167inter8));
  nand2 gate1844(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1845(.a(s_185), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1846(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1847(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1848(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2171(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2172(.a(gate169inter0), .b(s_232), .O(gate169inter1));
  and2  gate2173(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2174(.a(s_232), .O(gate169inter3));
  inv1  gate2175(.a(s_233), .O(gate169inter4));
  nand2 gate2176(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2177(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2178(.a(G474), .O(gate169inter7));
  inv1  gate2179(.a(G546), .O(gate169inter8));
  nand2 gate2180(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2181(.a(s_233), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2182(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2183(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2184(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1163(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1164(.a(gate170inter0), .b(s_88), .O(gate170inter1));
  and2  gate1165(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1166(.a(s_88), .O(gate170inter3));
  inv1  gate1167(.a(s_89), .O(gate170inter4));
  nand2 gate1168(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1169(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1170(.a(G477), .O(gate170inter7));
  inv1  gate1171(.a(G546), .O(gate170inter8));
  nand2 gate1172(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1173(.a(s_89), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1174(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1175(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1176(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate2843(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2844(.a(gate171inter0), .b(s_328), .O(gate171inter1));
  and2  gate2845(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2846(.a(s_328), .O(gate171inter3));
  inv1  gate2847(.a(s_329), .O(gate171inter4));
  nand2 gate2848(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2849(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2850(.a(G480), .O(gate171inter7));
  inv1  gate2851(.a(G549), .O(gate171inter8));
  nand2 gate2852(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2853(.a(s_329), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2854(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2855(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2856(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2045(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2046(.a(gate172inter0), .b(s_214), .O(gate172inter1));
  and2  gate2047(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2048(.a(s_214), .O(gate172inter3));
  inv1  gate2049(.a(s_215), .O(gate172inter4));
  nand2 gate2050(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2051(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2052(.a(G483), .O(gate172inter7));
  inv1  gate2053(.a(G549), .O(gate172inter8));
  nand2 gate2054(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2055(.a(s_215), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2056(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2057(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2058(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1555(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1556(.a(gate175inter0), .b(s_144), .O(gate175inter1));
  and2  gate1557(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1558(.a(s_144), .O(gate175inter3));
  inv1  gate1559(.a(s_145), .O(gate175inter4));
  nand2 gate1560(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1561(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1562(.a(G492), .O(gate175inter7));
  inv1  gate1563(.a(G555), .O(gate175inter8));
  nand2 gate1564(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1565(.a(s_145), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1566(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1567(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1568(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1681(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1682(.a(gate176inter0), .b(s_162), .O(gate176inter1));
  and2  gate1683(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1684(.a(s_162), .O(gate176inter3));
  inv1  gate1685(.a(s_163), .O(gate176inter4));
  nand2 gate1686(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1687(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1688(.a(G495), .O(gate176inter7));
  inv1  gate1689(.a(G555), .O(gate176inter8));
  nand2 gate1690(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1691(.a(s_163), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1692(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1693(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1694(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate2969(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2970(.a(gate177inter0), .b(s_346), .O(gate177inter1));
  and2  gate2971(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2972(.a(s_346), .O(gate177inter3));
  inv1  gate2973(.a(s_347), .O(gate177inter4));
  nand2 gate2974(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2975(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2976(.a(G498), .O(gate177inter7));
  inv1  gate2977(.a(G558), .O(gate177inter8));
  nand2 gate2978(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2979(.a(s_347), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2980(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2981(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2982(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1121(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1122(.a(gate182inter0), .b(s_82), .O(gate182inter1));
  and2  gate1123(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1124(.a(s_82), .O(gate182inter3));
  inv1  gate1125(.a(s_83), .O(gate182inter4));
  nand2 gate1126(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1127(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1128(.a(G513), .O(gate182inter7));
  inv1  gate1129(.a(G564), .O(gate182inter8));
  nand2 gate1130(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1131(.a(s_83), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1132(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1133(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1134(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate2283(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2284(.a(gate183inter0), .b(s_248), .O(gate183inter1));
  and2  gate2285(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2286(.a(s_248), .O(gate183inter3));
  inv1  gate2287(.a(s_249), .O(gate183inter4));
  nand2 gate2288(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2289(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2290(.a(G516), .O(gate183inter7));
  inv1  gate2291(.a(G567), .O(gate183inter8));
  nand2 gate2292(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2293(.a(s_249), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2294(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2295(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2296(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1989(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1990(.a(gate185inter0), .b(s_206), .O(gate185inter1));
  and2  gate1991(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1992(.a(s_206), .O(gate185inter3));
  inv1  gate1993(.a(s_207), .O(gate185inter4));
  nand2 gate1994(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1995(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1996(.a(G570), .O(gate185inter7));
  inv1  gate1997(.a(G571), .O(gate185inter8));
  nand2 gate1998(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1999(.a(s_207), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2000(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2001(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2002(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate799(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate800(.a(gate199inter0), .b(s_36), .O(gate199inter1));
  and2  gate801(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate802(.a(s_36), .O(gate199inter3));
  inv1  gate803(.a(s_37), .O(gate199inter4));
  nand2 gate804(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate805(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate806(.a(G598), .O(gate199inter7));
  inv1  gate807(.a(G599), .O(gate199inter8));
  nand2 gate808(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate809(.a(s_37), .b(gate199inter3), .O(gate199inter10));
  nor2  gate810(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate811(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate812(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1933(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1934(.a(gate203inter0), .b(s_198), .O(gate203inter1));
  and2  gate1935(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1936(.a(s_198), .O(gate203inter3));
  inv1  gate1937(.a(s_199), .O(gate203inter4));
  nand2 gate1938(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1939(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1940(.a(G602), .O(gate203inter7));
  inv1  gate1941(.a(G612), .O(gate203inter8));
  nand2 gate1942(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1943(.a(s_199), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1944(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1945(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1946(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate603(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate604(.a(gate205inter0), .b(s_8), .O(gate205inter1));
  and2  gate605(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate606(.a(s_8), .O(gate205inter3));
  inv1  gate607(.a(s_9), .O(gate205inter4));
  nand2 gate608(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate609(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate610(.a(G622), .O(gate205inter7));
  inv1  gate611(.a(G627), .O(gate205inter8));
  nand2 gate612(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate613(.a(s_9), .b(gate205inter3), .O(gate205inter10));
  nor2  gate614(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate615(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate616(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1373(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1374(.a(gate207inter0), .b(s_118), .O(gate207inter1));
  and2  gate1375(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1376(.a(s_118), .O(gate207inter3));
  inv1  gate1377(.a(s_119), .O(gate207inter4));
  nand2 gate1378(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1379(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1380(.a(G622), .O(gate207inter7));
  inv1  gate1381(.a(G632), .O(gate207inter8));
  nand2 gate1382(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1383(.a(s_119), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1384(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1385(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1386(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2325(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2326(.a(gate208inter0), .b(s_254), .O(gate208inter1));
  and2  gate2327(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2328(.a(s_254), .O(gate208inter3));
  inv1  gate2329(.a(s_255), .O(gate208inter4));
  nand2 gate2330(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2331(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2332(.a(G627), .O(gate208inter7));
  inv1  gate2333(.a(G637), .O(gate208inter8));
  nand2 gate2334(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2335(.a(s_255), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2336(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2337(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2338(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1709(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1710(.a(gate209inter0), .b(s_166), .O(gate209inter1));
  and2  gate1711(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1712(.a(s_166), .O(gate209inter3));
  inv1  gate1713(.a(s_167), .O(gate209inter4));
  nand2 gate1714(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1715(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1716(.a(G602), .O(gate209inter7));
  inv1  gate1717(.a(G666), .O(gate209inter8));
  nand2 gate1718(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1719(.a(s_167), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1720(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1721(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1722(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1919(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1920(.a(gate213inter0), .b(s_196), .O(gate213inter1));
  and2  gate1921(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1922(.a(s_196), .O(gate213inter3));
  inv1  gate1923(.a(s_197), .O(gate213inter4));
  nand2 gate1924(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1925(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1926(.a(G602), .O(gate213inter7));
  inv1  gate1927(.a(G672), .O(gate213inter8));
  nand2 gate1928(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1929(.a(s_197), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1930(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1931(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1932(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2605(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2606(.a(gate215inter0), .b(s_294), .O(gate215inter1));
  and2  gate2607(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2608(.a(s_294), .O(gate215inter3));
  inv1  gate2609(.a(s_295), .O(gate215inter4));
  nand2 gate2610(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2611(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2612(.a(G607), .O(gate215inter7));
  inv1  gate2613(.a(G675), .O(gate215inter8));
  nand2 gate2614(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2615(.a(s_295), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2616(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2617(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2618(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1261(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1262(.a(gate216inter0), .b(s_102), .O(gate216inter1));
  and2  gate1263(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1264(.a(s_102), .O(gate216inter3));
  inv1  gate1265(.a(s_103), .O(gate216inter4));
  nand2 gate1266(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1267(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1268(.a(G617), .O(gate216inter7));
  inv1  gate1269(.a(G675), .O(gate216inter8));
  nand2 gate1270(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1271(.a(s_103), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1272(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1273(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1274(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate617(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate618(.a(gate218inter0), .b(s_10), .O(gate218inter1));
  and2  gate619(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate620(.a(s_10), .O(gate218inter3));
  inv1  gate621(.a(s_11), .O(gate218inter4));
  nand2 gate622(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate623(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate624(.a(G627), .O(gate218inter7));
  inv1  gate625(.a(G678), .O(gate218inter8));
  nand2 gate626(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate627(.a(s_11), .b(gate218inter3), .O(gate218inter10));
  nor2  gate628(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate629(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate630(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate659(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate660(.a(gate220inter0), .b(s_16), .O(gate220inter1));
  and2  gate661(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate662(.a(s_16), .O(gate220inter3));
  inv1  gate663(.a(s_17), .O(gate220inter4));
  nand2 gate664(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate665(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate666(.a(G637), .O(gate220inter7));
  inv1  gate667(.a(G681), .O(gate220inter8));
  nand2 gate668(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate669(.a(s_17), .b(gate220inter3), .O(gate220inter10));
  nor2  gate670(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate671(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate672(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate2675(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2676(.a(gate221inter0), .b(s_304), .O(gate221inter1));
  and2  gate2677(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2678(.a(s_304), .O(gate221inter3));
  inv1  gate2679(.a(s_305), .O(gate221inter4));
  nand2 gate2680(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2681(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2682(.a(G622), .O(gate221inter7));
  inv1  gate2683(.a(G684), .O(gate221inter8));
  nand2 gate2684(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2685(.a(s_305), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2686(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2687(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2688(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate953(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate954(.a(gate226inter0), .b(s_58), .O(gate226inter1));
  and2  gate955(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate956(.a(s_58), .O(gate226inter3));
  inv1  gate957(.a(s_59), .O(gate226inter4));
  nand2 gate958(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate959(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate960(.a(G692), .O(gate226inter7));
  inv1  gate961(.a(G693), .O(gate226inter8));
  nand2 gate962(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate963(.a(s_59), .b(gate226inter3), .O(gate226inter10));
  nor2  gate964(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate965(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate966(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2409(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2410(.a(gate228inter0), .b(s_266), .O(gate228inter1));
  and2  gate2411(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2412(.a(s_266), .O(gate228inter3));
  inv1  gate2413(.a(s_267), .O(gate228inter4));
  nand2 gate2414(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2415(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2416(.a(G696), .O(gate228inter7));
  inv1  gate2417(.a(G697), .O(gate228inter8));
  nand2 gate2418(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2419(.a(s_267), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2420(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2421(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2422(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2339(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2340(.a(gate230inter0), .b(s_256), .O(gate230inter1));
  and2  gate2341(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2342(.a(s_256), .O(gate230inter3));
  inv1  gate2343(.a(s_257), .O(gate230inter4));
  nand2 gate2344(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2345(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2346(.a(G700), .O(gate230inter7));
  inv1  gate2347(.a(G701), .O(gate230inter8));
  nand2 gate2348(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2349(.a(s_257), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2350(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2351(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2352(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2227(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2228(.a(gate231inter0), .b(s_240), .O(gate231inter1));
  and2  gate2229(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2230(.a(s_240), .O(gate231inter3));
  inv1  gate2231(.a(s_241), .O(gate231inter4));
  nand2 gate2232(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2233(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2234(.a(G702), .O(gate231inter7));
  inv1  gate2235(.a(G703), .O(gate231inter8));
  nand2 gate2236(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2237(.a(s_241), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2238(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2239(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2240(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2087(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2088(.a(gate232inter0), .b(s_220), .O(gate232inter1));
  and2  gate2089(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2090(.a(s_220), .O(gate232inter3));
  inv1  gate2091(.a(s_221), .O(gate232inter4));
  nand2 gate2092(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2093(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2094(.a(G704), .O(gate232inter7));
  inv1  gate2095(.a(G705), .O(gate232inter8));
  nand2 gate2096(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2097(.a(s_221), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2098(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2099(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2100(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate547(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate548(.a(gate234inter0), .b(s_0), .O(gate234inter1));
  and2  gate549(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate550(.a(s_0), .O(gate234inter3));
  inv1  gate551(.a(s_1), .O(gate234inter4));
  nand2 gate552(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate553(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate554(.a(G245), .O(gate234inter7));
  inv1  gate555(.a(G721), .O(gate234inter8));
  nand2 gate556(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate557(.a(s_1), .b(gate234inter3), .O(gate234inter10));
  nor2  gate558(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate559(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate560(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1233(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1234(.a(gate235inter0), .b(s_98), .O(gate235inter1));
  and2  gate1235(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1236(.a(s_98), .O(gate235inter3));
  inv1  gate1237(.a(s_99), .O(gate235inter4));
  nand2 gate1238(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1239(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1240(.a(G248), .O(gate235inter7));
  inv1  gate1241(.a(G724), .O(gate235inter8));
  nand2 gate1242(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1243(.a(s_99), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1244(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1245(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1246(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1625(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1626(.a(gate237inter0), .b(s_154), .O(gate237inter1));
  and2  gate1627(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1628(.a(s_154), .O(gate237inter3));
  inv1  gate1629(.a(s_155), .O(gate237inter4));
  nand2 gate1630(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1631(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1632(.a(G254), .O(gate237inter7));
  inv1  gate1633(.a(G706), .O(gate237inter8));
  nand2 gate1634(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1635(.a(s_155), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1636(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1637(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1638(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1863(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1864(.a(gate239inter0), .b(s_188), .O(gate239inter1));
  and2  gate1865(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1866(.a(s_188), .O(gate239inter3));
  inv1  gate1867(.a(s_189), .O(gate239inter4));
  nand2 gate1868(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1869(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1870(.a(G260), .O(gate239inter7));
  inv1  gate1871(.a(G712), .O(gate239inter8));
  nand2 gate1872(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1873(.a(s_189), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1874(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1875(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1876(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2871(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2872(.a(gate242inter0), .b(s_332), .O(gate242inter1));
  and2  gate2873(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2874(.a(s_332), .O(gate242inter3));
  inv1  gate2875(.a(s_333), .O(gate242inter4));
  nand2 gate2876(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2877(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2878(.a(G718), .O(gate242inter7));
  inv1  gate2879(.a(G730), .O(gate242inter8));
  nand2 gate2880(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2881(.a(s_333), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2882(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2883(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2884(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1947(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1948(.a(gate243inter0), .b(s_200), .O(gate243inter1));
  and2  gate1949(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1950(.a(s_200), .O(gate243inter3));
  inv1  gate1951(.a(s_201), .O(gate243inter4));
  nand2 gate1952(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1953(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1954(.a(G245), .O(gate243inter7));
  inv1  gate1955(.a(G733), .O(gate243inter8));
  nand2 gate1956(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1957(.a(s_201), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1958(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1959(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1960(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1723(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1724(.a(gate248inter0), .b(s_168), .O(gate248inter1));
  and2  gate1725(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1726(.a(s_168), .O(gate248inter3));
  inv1  gate1727(.a(s_169), .O(gate248inter4));
  nand2 gate1728(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1729(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1730(.a(G727), .O(gate248inter7));
  inv1  gate1731(.a(G739), .O(gate248inter8));
  nand2 gate1732(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1733(.a(s_169), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1734(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1735(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1736(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate869(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate870(.a(gate249inter0), .b(s_46), .O(gate249inter1));
  and2  gate871(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate872(.a(s_46), .O(gate249inter3));
  inv1  gate873(.a(s_47), .O(gate249inter4));
  nand2 gate874(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate875(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate876(.a(G254), .O(gate249inter7));
  inv1  gate877(.a(G742), .O(gate249inter8));
  nand2 gate878(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate879(.a(s_47), .b(gate249inter3), .O(gate249inter10));
  nor2  gate880(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate881(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate882(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2829(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2830(.a(gate252inter0), .b(s_326), .O(gate252inter1));
  and2  gate2831(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2832(.a(s_326), .O(gate252inter3));
  inv1  gate2833(.a(s_327), .O(gate252inter4));
  nand2 gate2834(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2835(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2836(.a(G709), .O(gate252inter7));
  inv1  gate2837(.a(G745), .O(gate252inter8));
  nand2 gate2838(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2839(.a(s_327), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2840(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2841(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2842(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2577(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2578(.a(gate255inter0), .b(s_290), .O(gate255inter1));
  and2  gate2579(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2580(.a(s_290), .O(gate255inter3));
  inv1  gate2581(.a(s_291), .O(gate255inter4));
  nand2 gate2582(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2583(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2584(.a(G263), .O(gate255inter7));
  inv1  gate2585(.a(G751), .O(gate255inter8));
  nand2 gate2586(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2587(.a(s_291), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2588(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2589(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2590(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate715(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate716(.a(gate257inter0), .b(s_24), .O(gate257inter1));
  and2  gate717(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate718(.a(s_24), .O(gate257inter3));
  inv1  gate719(.a(s_25), .O(gate257inter4));
  nand2 gate720(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate721(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate722(.a(G754), .O(gate257inter7));
  inv1  gate723(.a(G755), .O(gate257inter8));
  nand2 gate724(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate725(.a(s_25), .b(gate257inter3), .O(gate257inter10));
  nor2  gate726(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate727(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate728(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate813(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate814(.a(gate268inter0), .b(s_38), .O(gate268inter1));
  and2  gate815(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate816(.a(s_38), .O(gate268inter3));
  inv1  gate817(.a(s_39), .O(gate268inter4));
  nand2 gate818(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate819(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate820(.a(G651), .O(gate268inter7));
  inv1  gate821(.a(G779), .O(gate268inter8));
  nand2 gate822(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate823(.a(s_39), .b(gate268inter3), .O(gate268inter10));
  nor2  gate824(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate825(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate826(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate2269(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2270(.a(gate269inter0), .b(s_246), .O(gate269inter1));
  and2  gate2271(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2272(.a(s_246), .O(gate269inter3));
  inv1  gate2273(.a(s_247), .O(gate269inter4));
  nand2 gate2274(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2275(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2276(.a(G654), .O(gate269inter7));
  inv1  gate2277(.a(G782), .O(gate269inter8));
  nand2 gate2278(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2279(.a(s_247), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2280(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2281(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2282(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2549(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2550(.a(gate277inter0), .b(s_286), .O(gate277inter1));
  and2  gate2551(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2552(.a(s_286), .O(gate277inter3));
  inv1  gate2553(.a(s_287), .O(gate277inter4));
  nand2 gate2554(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2555(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2556(.a(G648), .O(gate277inter7));
  inv1  gate2557(.a(G800), .O(gate277inter8));
  nand2 gate2558(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2559(.a(s_287), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2560(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2561(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2562(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1611(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1612(.a(gate278inter0), .b(s_152), .O(gate278inter1));
  and2  gate1613(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1614(.a(s_152), .O(gate278inter3));
  inv1  gate1615(.a(s_153), .O(gate278inter4));
  nand2 gate1616(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1617(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1618(.a(G776), .O(gate278inter7));
  inv1  gate1619(.a(G800), .O(gate278inter8));
  nand2 gate1620(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1621(.a(s_153), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1622(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1623(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1624(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2591(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2592(.a(gate281inter0), .b(s_292), .O(gate281inter1));
  and2  gate2593(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2594(.a(s_292), .O(gate281inter3));
  inv1  gate2595(.a(s_293), .O(gate281inter4));
  nand2 gate2596(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2597(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2598(.a(G654), .O(gate281inter7));
  inv1  gate2599(.a(G806), .O(gate281inter8));
  nand2 gate2600(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2601(.a(s_293), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2602(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2603(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2604(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1667(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1668(.a(gate282inter0), .b(s_160), .O(gate282inter1));
  and2  gate1669(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1670(.a(s_160), .O(gate282inter3));
  inv1  gate1671(.a(s_161), .O(gate282inter4));
  nand2 gate1672(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1673(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1674(.a(G782), .O(gate282inter7));
  inv1  gate1675(.a(G806), .O(gate282inter8));
  nand2 gate1676(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1677(.a(s_161), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1678(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1679(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1680(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2143(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2144(.a(gate283inter0), .b(s_228), .O(gate283inter1));
  and2  gate2145(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2146(.a(s_228), .O(gate283inter3));
  inv1  gate2147(.a(s_229), .O(gate283inter4));
  nand2 gate2148(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2149(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2150(.a(G657), .O(gate283inter7));
  inv1  gate2151(.a(G809), .O(gate283inter8));
  nand2 gate2152(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2153(.a(s_229), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2154(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2155(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2156(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1877(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1878(.a(gate284inter0), .b(s_190), .O(gate284inter1));
  and2  gate1879(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1880(.a(s_190), .O(gate284inter3));
  inv1  gate1881(.a(s_191), .O(gate284inter4));
  nand2 gate1882(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1883(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1884(.a(G785), .O(gate284inter7));
  inv1  gate1885(.a(G809), .O(gate284inter8));
  nand2 gate1886(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1887(.a(s_191), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1888(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1889(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1890(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2451(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2452(.a(gate285inter0), .b(s_272), .O(gate285inter1));
  and2  gate2453(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2454(.a(s_272), .O(gate285inter3));
  inv1  gate2455(.a(s_273), .O(gate285inter4));
  nand2 gate2456(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2457(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2458(.a(G660), .O(gate285inter7));
  inv1  gate2459(.a(G812), .O(gate285inter8));
  nand2 gate2460(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2461(.a(s_273), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2462(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2463(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2464(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2353(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2354(.a(gate288inter0), .b(s_258), .O(gate288inter1));
  and2  gate2355(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2356(.a(s_258), .O(gate288inter3));
  inv1  gate2357(.a(s_259), .O(gate288inter4));
  nand2 gate2358(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2359(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2360(.a(G791), .O(gate288inter7));
  inv1  gate2361(.a(G815), .O(gate288inter8));
  nand2 gate2362(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2363(.a(s_259), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2364(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2365(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2366(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate995(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate996(.a(gate289inter0), .b(s_64), .O(gate289inter1));
  and2  gate997(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate998(.a(s_64), .O(gate289inter3));
  inv1  gate999(.a(s_65), .O(gate289inter4));
  nand2 gate1000(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1001(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1002(.a(G818), .O(gate289inter7));
  inv1  gate1003(.a(G819), .O(gate289inter8));
  nand2 gate1004(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1005(.a(s_65), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1006(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1007(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1008(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate2535(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2536(.a(gate290inter0), .b(s_284), .O(gate290inter1));
  and2  gate2537(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2538(.a(s_284), .O(gate290inter3));
  inv1  gate2539(.a(s_285), .O(gate290inter4));
  nand2 gate2540(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2541(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2542(.a(G820), .O(gate290inter7));
  inv1  gate2543(.a(G821), .O(gate290inter8));
  nand2 gate2544(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2545(.a(s_285), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2546(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2547(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2548(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1177(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1178(.a(gate294inter0), .b(s_90), .O(gate294inter1));
  and2  gate1179(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1180(.a(s_90), .O(gate294inter3));
  inv1  gate1181(.a(s_91), .O(gate294inter4));
  nand2 gate1182(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1183(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1184(.a(G832), .O(gate294inter7));
  inv1  gate1185(.a(G833), .O(gate294inter8));
  nand2 gate1186(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1187(.a(s_91), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1188(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1189(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1190(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2479(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2480(.a(gate295inter0), .b(s_276), .O(gate295inter1));
  and2  gate2481(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2482(.a(s_276), .O(gate295inter3));
  inv1  gate2483(.a(s_277), .O(gate295inter4));
  nand2 gate2484(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2485(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2486(.a(G830), .O(gate295inter7));
  inv1  gate2487(.a(G831), .O(gate295inter8));
  nand2 gate2488(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2489(.a(s_277), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2490(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2491(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2492(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2129(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2130(.a(gate387inter0), .b(s_226), .O(gate387inter1));
  and2  gate2131(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2132(.a(s_226), .O(gate387inter3));
  inv1  gate2133(.a(s_227), .O(gate387inter4));
  nand2 gate2134(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2135(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2136(.a(G1), .O(gate387inter7));
  inv1  gate2137(.a(G1036), .O(gate387inter8));
  nand2 gate2138(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2139(.a(s_227), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2140(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2141(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2142(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate2731(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2732(.a(gate390inter0), .b(s_312), .O(gate390inter1));
  and2  gate2733(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2734(.a(s_312), .O(gate390inter3));
  inv1  gate2735(.a(s_313), .O(gate390inter4));
  nand2 gate2736(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2737(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2738(.a(G4), .O(gate390inter7));
  inv1  gate2739(.a(G1045), .O(gate390inter8));
  nand2 gate2740(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2741(.a(s_313), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2742(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2743(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2744(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate2927(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2928(.a(gate391inter0), .b(s_340), .O(gate391inter1));
  and2  gate2929(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2930(.a(s_340), .O(gate391inter3));
  inv1  gate2931(.a(s_341), .O(gate391inter4));
  nand2 gate2932(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2933(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2934(.a(G5), .O(gate391inter7));
  inv1  gate2935(.a(G1048), .O(gate391inter8));
  nand2 gate2936(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2937(.a(s_341), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2938(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2939(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2940(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1597(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1598(.a(gate393inter0), .b(s_150), .O(gate393inter1));
  and2  gate1599(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1600(.a(s_150), .O(gate393inter3));
  inv1  gate1601(.a(s_151), .O(gate393inter4));
  nand2 gate1602(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1603(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1604(.a(G7), .O(gate393inter7));
  inv1  gate1605(.a(G1054), .O(gate393inter8));
  nand2 gate1606(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1607(.a(s_151), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1608(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1609(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1610(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate771(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate772(.a(gate394inter0), .b(s_32), .O(gate394inter1));
  and2  gate773(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate774(.a(s_32), .O(gate394inter3));
  inv1  gate775(.a(s_33), .O(gate394inter4));
  nand2 gate776(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate777(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate778(.a(G8), .O(gate394inter7));
  inv1  gate779(.a(G1057), .O(gate394inter8));
  nand2 gate780(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate781(.a(s_33), .b(gate394inter3), .O(gate394inter10));
  nor2  gate782(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate783(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate784(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1905(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1906(.a(gate400inter0), .b(s_194), .O(gate400inter1));
  and2  gate1907(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1908(.a(s_194), .O(gate400inter3));
  inv1  gate1909(.a(s_195), .O(gate400inter4));
  nand2 gate1910(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1911(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1912(.a(G14), .O(gate400inter7));
  inv1  gate1913(.a(G1075), .O(gate400inter8));
  nand2 gate1914(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1915(.a(s_195), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1916(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1917(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1918(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate925(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate926(.a(gate406inter0), .b(s_54), .O(gate406inter1));
  and2  gate927(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate928(.a(s_54), .O(gate406inter3));
  inv1  gate929(.a(s_55), .O(gate406inter4));
  nand2 gate930(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate931(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate932(.a(G20), .O(gate406inter7));
  inv1  gate933(.a(G1093), .O(gate406inter8));
  nand2 gate934(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate935(.a(s_55), .b(gate406inter3), .O(gate406inter10));
  nor2  gate936(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate937(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate938(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1331(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1332(.a(gate409inter0), .b(s_112), .O(gate409inter1));
  and2  gate1333(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1334(.a(s_112), .O(gate409inter3));
  inv1  gate1335(.a(s_113), .O(gate409inter4));
  nand2 gate1336(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1337(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1338(.a(G23), .O(gate409inter7));
  inv1  gate1339(.a(G1102), .O(gate409inter8));
  nand2 gate1340(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1341(.a(s_113), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1342(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1343(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1344(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2381(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2382(.a(gate410inter0), .b(s_262), .O(gate410inter1));
  and2  gate2383(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2384(.a(s_262), .O(gate410inter3));
  inv1  gate2385(.a(s_263), .O(gate410inter4));
  nand2 gate2386(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2387(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2388(.a(G24), .O(gate410inter7));
  inv1  gate2389(.a(G1105), .O(gate410inter8));
  nand2 gate2390(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2391(.a(s_263), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2392(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2393(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2394(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1513(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1514(.a(gate412inter0), .b(s_138), .O(gate412inter1));
  and2  gate1515(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1516(.a(s_138), .O(gate412inter3));
  inv1  gate1517(.a(s_139), .O(gate412inter4));
  nand2 gate1518(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1519(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1520(.a(G26), .O(gate412inter7));
  inv1  gate1521(.a(G1111), .O(gate412inter8));
  nand2 gate1522(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1523(.a(s_139), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1524(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1525(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1526(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1149(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1150(.a(gate417inter0), .b(s_86), .O(gate417inter1));
  and2  gate1151(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1152(.a(s_86), .O(gate417inter3));
  inv1  gate1153(.a(s_87), .O(gate417inter4));
  nand2 gate1154(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1155(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1156(.a(G31), .O(gate417inter7));
  inv1  gate1157(.a(G1126), .O(gate417inter8));
  nand2 gate1158(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1159(.a(s_87), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1160(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1161(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1162(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2703(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2704(.a(gate418inter0), .b(s_308), .O(gate418inter1));
  and2  gate2705(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2706(.a(s_308), .O(gate418inter3));
  inv1  gate2707(.a(s_309), .O(gate418inter4));
  nand2 gate2708(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2709(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2710(.a(G32), .O(gate418inter7));
  inv1  gate2711(.a(G1129), .O(gate418inter8));
  nand2 gate2712(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2713(.a(s_309), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2714(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2715(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2716(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1765(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1766(.a(gate419inter0), .b(s_174), .O(gate419inter1));
  and2  gate1767(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1768(.a(s_174), .O(gate419inter3));
  inv1  gate1769(.a(s_175), .O(gate419inter4));
  nand2 gate1770(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1771(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1772(.a(G1), .O(gate419inter7));
  inv1  gate1773(.a(G1132), .O(gate419inter8));
  nand2 gate1774(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1775(.a(s_175), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1776(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1777(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1778(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1107(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1108(.a(gate421inter0), .b(s_80), .O(gate421inter1));
  and2  gate1109(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1110(.a(s_80), .O(gate421inter3));
  inv1  gate1111(.a(s_81), .O(gate421inter4));
  nand2 gate1112(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1113(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1114(.a(G2), .O(gate421inter7));
  inv1  gate1115(.a(G1135), .O(gate421inter8));
  nand2 gate1116(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1117(.a(s_81), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1118(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1119(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1120(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1303(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1304(.a(gate422inter0), .b(s_108), .O(gate422inter1));
  and2  gate1305(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1306(.a(s_108), .O(gate422inter3));
  inv1  gate1307(.a(s_109), .O(gate422inter4));
  nand2 gate1308(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1309(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1310(.a(G1039), .O(gate422inter7));
  inv1  gate1311(.a(G1135), .O(gate422inter8));
  nand2 gate1312(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1313(.a(s_109), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1314(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1315(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1316(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate2031(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2032(.a(gate423inter0), .b(s_212), .O(gate423inter1));
  and2  gate2033(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2034(.a(s_212), .O(gate423inter3));
  inv1  gate2035(.a(s_213), .O(gate423inter4));
  nand2 gate2036(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2037(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2038(.a(G3), .O(gate423inter7));
  inv1  gate2039(.a(G1138), .O(gate423inter8));
  nand2 gate2040(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2041(.a(s_213), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2042(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2043(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2044(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2661(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2662(.a(gate424inter0), .b(s_302), .O(gate424inter1));
  and2  gate2663(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2664(.a(s_302), .O(gate424inter3));
  inv1  gate2665(.a(s_303), .O(gate424inter4));
  nand2 gate2666(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2667(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2668(.a(G1042), .O(gate424inter7));
  inv1  gate2669(.a(G1138), .O(gate424inter8));
  nand2 gate2670(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2671(.a(s_303), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2672(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2673(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2674(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate841(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate842(.a(gate426inter0), .b(s_42), .O(gate426inter1));
  and2  gate843(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate844(.a(s_42), .O(gate426inter3));
  inv1  gate845(.a(s_43), .O(gate426inter4));
  nand2 gate846(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate847(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate848(.a(G1045), .O(gate426inter7));
  inv1  gate849(.a(G1141), .O(gate426inter8));
  nand2 gate850(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate851(.a(s_43), .b(gate426inter3), .O(gate426inter10));
  nor2  gate852(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate853(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate854(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2003(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2004(.a(gate428inter0), .b(s_208), .O(gate428inter1));
  and2  gate2005(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2006(.a(s_208), .O(gate428inter3));
  inv1  gate2007(.a(s_209), .O(gate428inter4));
  nand2 gate2008(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2009(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2010(.a(G1048), .O(gate428inter7));
  inv1  gate2011(.a(G1144), .O(gate428inter8));
  nand2 gate2012(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2013(.a(s_209), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2014(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2015(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2016(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate827(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate828(.a(gate436inter0), .b(s_40), .O(gate436inter1));
  and2  gate829(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate830(.a(s_40), .O(gate436inter3));
  inv1  gate831(.a(s_41), .O(gate436inter4));
  nand2 gate832(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate833(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate834(.a(G1060), .O(gate436inter7));
  inv1  gate835(.a(G1156), .O(gate436inter8));
  nand2 gate836(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate837(.a(s_41), .b(gate436inter3), .O(gate436inter10));
  nor2  gate838(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate839(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate840(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1779(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1780(.a(gate437inter0), .b(s_176), .O(gate437inter1));
  and2  gate1781(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1782(.a(s_176), .O(gate437inter3));
  inv1  gate1783(.a(s_177), .O(gate437inter4));
  nand2 gate1784(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1785(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1786(.a(G10), .O(gate437inter7));
  inv1  gate1787(.a(G1159), .O(gate437inter8));
  nand2 gate1788(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1789(.a(s_177), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1790(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1791(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1792(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1317(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1318(.a(gate438inter0), .b(s_110), .O(gate438inter1));
  and2  gate1319(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1320(.a(s_110), .O(gate438inter3));
  inv1  gate1321(.a(s_111), .O(gate438inter4));
  nand2 gate1322(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1323(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1324(.a(G1063), .O(gate438inter7));
  inv1  gate1325(.a(G1159), .O(gate438inter8));
  nand2 gate1326(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1327(.a(s_111), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1328(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1329(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1330(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1415(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1416(.a(gate439inter0), .b(s_124), .O(gate439inter1));
  and2  gate1417(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1418(.a(s_124), .O(gate439inter3));
  inv1  gate1419(.a(s_125), .O(gate439inter4));
  nand2 gate1420(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1421(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1422(.a(G11), .O(gate439inter7));
  inv1  gate1423(.a(G1162), .O(gate439inter8));
  nand2 gate1424(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1425(.a(s_125), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1426(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1427(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1428(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1961(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1962(.a(gate440inter0), .b(s_202), .O(gate440inter1));
  and2  gate1963(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1964(.a(s_202), .O(gate440inter3));
  inv1  gate1965(.a(s_203), .O(gate440inter4));
  nand2 gate1966(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1967(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1968(.a(G1066), .O(gate440inter7));
  inv1  gate1969(.a(G1162), .O(gate440inter8));
  nand2 gate1970(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1971(.a(s_203), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1972(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1973(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1974(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1639(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1640(.a(gate445inter0), .b(s_156), .O(gate445inter1));
  and2  gate1641(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1642(.a(s_156), .O(gate445inter3));
  inv1  gate1643(.a(s_157), .O(gate445inter4));
  nand2 gate1644(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1645(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1646(.a(G14), .O(gate445inter7));
  inv1  gate1647(.a(G1171), .O(gate445inter8));
  nand2 gate1648(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1649(.a(s_157), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1650(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1651(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1652(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate673(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate674(.a(gate448inter0), .b(s_18), .O(gate448inter1));
  and2  gate675(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate676(.a(s_18), .O(gate448inter3));
  inv1  gate677(.a(s_19), .O(gate448inter4));
  nand2 gate678(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate679(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate680(.a(G1078), .O(gate448inter7));
  inv1  gate681(.a(G1174), .O(gate448inter8));
  nand2 gate682(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate683(.a(s_19), .b(gate448inter3), .O(gate448inter10));
  nor2  gate684(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate685(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate686(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2717(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2718(.a(gate451inter0), .b(s_310), .O(gate451inter1));
  and2  gate2719(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2720(.a(s_310), .O(gate451inter3));
  inv1  gate2721(.a(s_311), .O(gate451inter4));
  nand2 gate2722(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2723(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2724(.a(G17), .O(gate451inter7));
  inv1  gate2725(.a(G1180), .O(gate451inter8));
  nand2 gate2726(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2727(.a(s_311), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2728(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2729(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2730(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2157(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2158(.a(gate453inter0), .b(s_230), .O(gate453inter1));
  and2  gate2159(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2160(.a(s_230), .O(gate453inter3));
  inv1  gate2161(.a(s_231), .O(gate453inter4));
  nand2 gate2162(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2163(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2164(.a(G18), .O(gate453inter7));
  inv1  gate2165(.a(G1183), .O(gate453inter8));
  nand2 gate2166(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2167(.a(s_231), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2168(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2169(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2170(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1569(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1570(.a(gate455inter0), .b(s_146), .O(gate455inter1));
  and2  gate1571(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1572(.a(s_146), .O(gate455inter3));
  inv1  gate1573(.a(s_147), .O(gate455inter4));
  nand2 gate1574(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1575(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1576(.a(G19), .O(gate455inter7));
  inv1  gate1577(.a(G1186), .O(gate455inter8));
  nand2 gate1578(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1579(.a(s_147), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1580(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1581(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1582(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate855(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate856(.a(gate458inter0), .b(s_44), .O(gate458inter1));
  and2  gate857(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate858(.a(s_44), .O(gate458inter3));
  inv1  gate859(.a(s_45), .O(gate458inter4));
  nand2 gate860(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate861(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate862(.a(G1093), .O(gate458inter7));
  inv1  gate863(.a(G1189), .O(gate458inter8));
  nand2 gate864(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate865(.a(s_45), .b(gate458inter3), .O(gate458inter10));
  nor2  gate866(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate867(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate868(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1205(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1206(.a(gate460inter0), .b(s_94), .O(gate460inter1));
  and2  gate1207(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1208(.a(s_94), .O(gate460inter3));
  inv1  gate1209(.a(s_95), .O(gate460inter4));
  nand2 gate1210(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1211(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1212(.a(G1096), .O(gate460inter7));
  inv1  gate1213(.a(G1192), .O(gate460inter8));
  nand2 gate1214(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1215(.a(s_95), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1216(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1217(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1218(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2885(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2886(.a(gate462inter0), .b(s_334), .O(gate462inter1));
  and2  gate2887(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2888(.a(s_334), .O(gate462inter3));
  inv1  gate2889(.a(s_335), .O(gate462inter4));
  nand2 gate2890(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2891(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2892(.a(G1099), .O(gate462inter7));
  inv1  gate2893(.a(G1195), .O(gate462inter8));
  nand2 gate2894(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2895(.a(s_335), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2896(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2897(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2898(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1037(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1038(.a(gate469inter0), .b(s_70), .O(gate469inter1));
  and2  gate1039(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1040(.a(s_70), .O(gate469inter3));
  inv1  gate1041(.a(s_71), .O(gate469inter4));
  nand2 gate1042(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1043(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1044(.a(G26), .O(gate469inter7));
  inv1  gate1045(.a(G1207), .O(gate469inter8));
  nand2 gate1046(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1047(.a(s_71), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1048(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1049(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1050(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2437(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2438(.a(gate471inter0), .b(s_270), .O(gate471inter1));
  and2  gate2439(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2440(.a(s_270), .O(gate471inter3));
  inv1  gate2441(.a(s_271), .O(gate471inter4));
  nand2 gate2442(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2443(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2444(.a(G27), .O(gate471inter7));
  inv1  gate2445(.a(G1210), .O(gate471inter8));
  nand2 gate2446(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2447(.a(s_271), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2448(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2449(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2450(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2815(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2816(.a(gate472inter0), .b(s_324), .O(gate472inter1));
  and2  gate2817(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2818(.a(s_324), .O(gate472inter3));
  inv1  gate2819(.a(s_325), .O(gate472inter4));
  nand2 gate2820(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2821(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2822(.a(G1114), .O(gate472inter7));
  inv1  gate2823(.a(G1210), .O(gate472inter8));
  nand2 gate2824(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2825(.a(s_325), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2826(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2827(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2828(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1023(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1024(.a(gate475inter0), .b(s_68), .O(gate475inter1));
  and2  gate1025(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1026(.a(s_68), .O(gate475inter3));
  inv1  gate1027(.a(s_69), .O(gate475inter4));
  nand2 gate1028(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1029(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1030(.a(G29), .O(gate475inter7));
  inv1  gate1031(.a(G1216), .O(gate475inter8));
  nand2 gate1032(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1033(.a(s_69), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1034(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1035(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1036(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate939(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate940(.a(gate476inter0), .b(s_56), .O(gate476inter1));
  and2  gate941(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate942(.a(s_56), .O(gate476inter3));
  inv1  gate943(.a(s_57), .O(gate476inter4));
  nand2 gate944(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate945(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate946(.a(G1120), .O(gate476inter7));
  inv1  gate947(.a(G1216), .O(gate476inter8));
  nand2 gate948(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate949(.a(s_57), .b(gate476inter3), .O(gate476inter10));
  nor2  gate950(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate951(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate952(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1009(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1010(.a(gate478inter0), .b(s_66), .O(gate478inter1));
  and2  gate1011(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1012(.a(s_66), .O(gate478inter3));
  inv1  gate1013(.a(s_67), .O(gate478inter4));
  nand2 gate1014(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1015(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1016(.a(G1123), .O(gate478inter7));
  inv1  gate1017(.a(G1219), .O(gate478inter8));
  nand2 gate1018(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1019(.a(s_67), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1020(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1021(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1022(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2297(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2298(.a(gate479inter0), .b(s_250), .O(gate479inter1));
  and2  gate2299(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2300(.a(s_250), .O(gate479inter3));
  inv1  gate2301(.a(s_251), .O(gate479inter4));
  nand2 gate2302(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2303(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2304(.a(G31), .O(gate479inter7));
  inv1  gate2305(.a(G1222), .O(gate479inter8));
  nand2 gate2306(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2307(.a(s_251), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2308(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2309(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2310(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2101(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2102(.a(gate482inter0), .b(s_222), .O(gate482inter1));
  and2  gate2103(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2104(.a(s_222), .O(gate482inter3));
  inv1  gate2105(.a(s_223), .O(gate482inter4));
  nand2 gate2106(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2107(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2108(.a(G1129), .O(gate482inter7));
  inv1  gate2109(.a(G1225), .O(gate482inter8));
  nand2 gate2110(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2111(.a(s_223), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2112(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2113(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2114(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate2115(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2116(.a(gate484inter0), .b(s_224), .O(gate484inter1));
  and2  gate2117(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2118(.a(s_224), .O(gate484inter3));
  inv1  gate2119(.a(s_225), .O(gate484inter4));
  nand2 gate2120(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2121(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2122(.a(G1230), .O(gate484inter7));
  inv1  gate2123(.a(G1231), .O(gate484inter8));
  nand2 gate2124(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2125(.a(s_225), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2126(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2127(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2128(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate561(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate562(.a(gate489inter0), .b(s_2), .O(gate489inter1));
  and2  gate563(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate564(.a(s_2), .O(gate489inter3));
  inv1  gate565(.a(s_3), .O(gate489inter4));
  nand2 gate566(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate567(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate568(.a(G1240), .O(gate489inter7));
  inv1  gate569(.a(G1241), .O(gate489inter8));
  nand2 gate570(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate571(.a(s_3), .b(gate489inter3), .O(gate489inter10));
  nor2  gate572(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate573(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate574(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate687(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate688(.a(gate491inter0), .b(s_20), .O(gate491inter1));
  and2  gate689(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate690(.a(s_20), .O(gate491inter3));
  inv1  gate691(.a(s_21), .O(gate491inter4));
  nand2 gate692(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate693(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate694(.a(G1244), .O(gate491inter7));
  inv1  gate695(.a(G1245), .O(gate491inter8));
  nand2 gate696(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate697(.a(s_21), .b(gate491inter3), .O(gate491inter10));
  nor2  gate698(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate699(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate700(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1499(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1500(.a(gate495inter0), .b(s_136), .O(gate495inter1));
  and2  gate1501(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1502(.a(s_136), .O(gate495inter3));
  inv1  gate1503(.a(s_137), .O(gate495inter4));
  nand2 gate1504(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1505(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1506(.a(G1252), .O(gate495inter7));
  inv1  gate1507(.a(G1253), .O(gate495inter8));
  nand2 gate1508(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1509(.a(s_137), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1510(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1511(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1512(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate2647(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2648(.a(gate498inter0), .b(s_300), .O(gate498inter1));
  and2  gate2649(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2650(.a(s_300), .O(gate498inter3));
  inv1  gate2651(.a(s_301), .O(gate498inter4));
  nand2 gate2652(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2653(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2654(.a(G1258), .O(gate498inter7));
  inv1  gate2655(.a(G1259), .O(gate498inter8));
  nand2 gate2656(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2657(.a(s_301), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2658(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2659(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2660(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate631(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate632(.a(gate500inter0), .b(s_12), .O(gate500inter1));
  and2  gate633(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate634(.a(s_12), .O(gate500inter3));
  inv1  gate635(.a(s_13), .O(gate500inter4));
  nand2 gate636(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate637(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate638(.a(G1262), .O(gate500inter7));
  inv1  gate639(.a(G1263), .O(gate500inter8));
  nand2 gate640(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate641(.a(s_13), .b(gate500inter3), .O(gate500inter10));
  nor2  gate642(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate643(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate644(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate589(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate590(.a(gate502inter0), .b(s_6), .O(gate502inter1));
  and2  gate591(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate592(.a(s_6), .O(gate502inter3));
  inv1  gate593(.a(s_7), .O(gate502inter4));
  nand2 gate594(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate595(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate596(.a(G1266), .O(gate502inter7));
  inv1  gate597(.a(G1267), .O(gate502inter8));
  nand2 gate598(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate599(.a(s_7), .b(gate502inter3), .O(gate502inter10));
  nor2  gate600(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate601(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate602(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1387(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1388(.a(gate506inter0), .b(s_120), .O(gate506inter1));
  and2  gate1389(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1390(.a(s_120), .O(gate506inter3));
  inv1  gate1391(.a(s_121), .O(gate506inter4));
  nand2 gate1392(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1393(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1394(.a(G1274), .O(gate506inter7));
  inv1  gate1395(.a(G1275), .O(gate506inter8));
  nand2 gate1396(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1397(.a(s_121), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1398(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1399(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1400(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1583(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1584(.a(gate510inter0), .b(s_148), .O(gate510inter1));
  and2  gate1585(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1586(.a(s_148), .O(gate510inter3));
  inv1  gate1587(.a(s_149), .O(gate510inter4));
  nand2 gate1588(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1589(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1590(.a(G1282), .O(gate510inter7));
  inv1  gate1591(.a(G1283), .O(gate510inter8));
  nand2 gate1592(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1593(.a(s_149), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1594(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1595(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1596(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1191(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1192(.a(gate511inter0), .b(s_92), .O(gate511inter1));
  and2  gate1193(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1194(.a(s_92), .O(gate511inter3));
  inv1  gate1195(.a(s_93), .O(gate511inter4));
  nand2 gate1196(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1197(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1198(.a(G1284), .O(gate511inter7));
  inv1  gate1199(.a(G1285), .O(gate511inter8));
  nand2 gate1200(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1201(.a(s_93), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1202(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1203(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1204(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate729(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate730(.a(gate514inter0), .b(s_26), .O(gate514inter1));
  and2  gate731(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate732(.a(s_26), .O(gate514inter3));
  inv1  gate733(.a(s_27), .O(gate514inter4));
  nand2 gate734(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate735(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate736(.a(G1290), .O(gate514inter7));
  inv1  gate737(.a(G1291), .O(gate514inter8));
  nand2 gate738(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate739(.a(s_27), .b(gate514inter3), .O(gate514inter10));
  nor2  gate740(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate741(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate742(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule