module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate7inter0, gate7inter1, gate7inter2, gate7inter3, gate7inter4, gate7inter5, gate7inter6, gate7inter7, gate7inter8, gate7inter9, gate7inter10, gate7inter11, gate7inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );

  xor2  gate567(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate568(.a(gate5inter0), .b(s_52), .O(gate5inter1));
  and2  gate569(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate570(.a(s_52), .O(gate5inter3));
  inv1  gate571(.a(s_53), .O(gate5inter4));
  nand2 gate572(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate573(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate574(.a(N33), .O(gate5inter7));
  inv1  gate575(.a(N37), .O(gate5inter8));
  nand2 gate576(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate577(.a(s_53), .b(gate5inter3), .O(gate5inter10));
  nor2  gate578(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate579(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate580(.a(gate5inter12), .b(gate5inter1), .O(N254));
xor2 gate6( .a(N41), .b(N45), .O(N255) );

  xor2  gate301(.a(N53), .b(N49), .O(gate7inter0));
  nand2 gate302(.a(gate7inter0), .b(s_14), .O(gate7inter1));
  and2  gate303(.a(N53), .b(N49), .O(gate7inter2));
  inv1  gate304(.a(s_14), .O(gate7inter3));
  inv1  gate305(.a(s_15), .O(gate7inter4));
  nand2 gate306(.a(gate7inter4), .b(gate7inter3), .O(gate7inter5));
  nor2  gate307(.a(gate7inter5), .b(gate7inter2), .O(gate7inter6));
  inv1  gate308(.a(N49), .O(gate7inter7));
  inv1  gate309(.a(N53), .O(gate7inter8));
  nand2 gate310(.a(gate7inter8), .b(gate7inter7), .O(gate7inter9));
  nand2 gate311(.a(s_15), .b(gate7inter3), .O(gate7inter10));
  nor2  gate312(.a(gate7inter10), .b(gate7inter9), .O(gate7inter11));
  nor2  gate313(.a(gate7inter11), .b(gate7inter6), .O(gate7inter12));
  nand2 gate314(.a(gate7inter12), .b(gate7inter1), .O(N256));
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );

  xor2  gate329(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate330(.a(gate15inter0), .b(s_18), .O(gate15inter1));
  and2  gate331(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate332(.a(s_18), .O(gate15inter3));
  inv1  gate333(.a(s_19), .O(gate15inter4));
  nand2 gate334(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate335(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate336(.a(N113), .O(gate15inter7));
  inv1  gate337(.a(N117), .O(gate15inter8));
  nand2 gate338(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate339(.a(s_19), .b(gate15inter3), .O(gate15inter10));
  nor2  gate340(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate341(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate342(.a(gate15inter12), .b(gate15inter1), .O(N264));
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );

  xor2  gate497(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate498(.a(gate32inter0), .b(s_42), .O(gate32inter1));
  and2  gate499(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate500(.a(s_42), .O(gate32inter3));
  inv1  gate501(.a(s_43), .O(gate32inter4));
  nand2 gate502(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate503(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate504(.a(N45), .O(gate32inter7));
  inv1  gate505(.a(N61), .O(gate32inter8));
  nand2 gate506(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate507(.a(s_43), .b(gate32inter3), .O(gate32inter10));
  nor2  gate508(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate509(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate510(.a(gate32inter12), .b(gate32inter1), .O(N281));
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );

  xor2  gate553(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate554(.a(gate36inter0), .b(s_50), .O(gate36inter1));
  and2  gate555(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate556(.a(s_50), .O(gate36inter3));
  inv1  gate557(.a(s_51), .O(gate36inter4));
  nand2 gate558(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate559(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate560(.a(N101), .O(gate36inter7));
  inv1  gate561(.a(N117), .O(gate36inter8));
  nand2 gate562(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate563(.a(s_51), .b(gate36inter3), .O(gate36inter10));
  nor2  gate564(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate565(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate566(.a(gate36inter12), .b(gate36inter1), .O(N285));
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );

  xor2  gate595(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate596(.a(gate40inter0), .b(s_56), .O(gate40inter1));
  and2  gate597(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate598(.a(s_56), .O(gate40inter3));
  inv1  gate599(.a(s_57), .O(gate40inter4));
  nand2 gate600(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate601(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate602(.a(N109), .O(gate40inter7));
  inv1  gate603(.a(N125), .O(gate40inter8));
  nand2 gate604(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate605(.a(s_57), .b(gate40inter3), .O(gate40inter10));
  nor2  gate606(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate607(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate608(.a(gate40inter12), .b(gate40inter1), .O(N289));

  xor2  gate483(.a(N251), .b(N250), .O(gate41inter0));
  nand2 gate484(.a(gate41inter0), .b(s_40), .O(gate41inter1));
  and2  gate485(.a(N251), .b(N250), .O(gate41inter2));
  inv1  gate486(.a(s_40), .O(gate41inter3));
  inv1  gate487(.a(s_41), .O(gate41inter4));
  nand2 gate488(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate489(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate490(.a(N250), .O(gate41inter7));
  inv1  gate491(.a(N251), .O(gate41inter8));
  nand2 gate492(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate493(.a(s_41), .b(gate41inter3), .O(gate41inter10));
  nor2  gate494(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate495(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate496(.a(gate41inter12), .b(gate41inter1), .O(N290));

  xor2  gate371(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate372(.a(gate42inter0), .b(s_24), .O(gate42inter1));
  and2  gate373(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate374(.a(s_24), .O(gate42inter3));
  inv1  gate375(.a(s_25), .O(gate42inter4));
  nand2 gate376(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate377(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate378(.a(N252), .O(gate42inter7));
  inv1  gate379(.a(N253), .O(gate42inter8));
  nand2 gate380(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate381(.a(s_25), .b(gate42inter3), .O(gate42inter10));
  nor2  gate382(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate383(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate384(.a(gate42inter12), .b(gate42inter1), .O(N293));
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );

  xor2  gate357(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate358(.a(gate54inter0), .b(s_22), .O(gate54inter1));
  and2  gate359(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate360(.a(s_22), .O(gate54inter3));
  inv1  gate361(.a(s_23), .O(gate54inter4));
  nand2 gate362(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate363(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate364(.a(N284), .O(gate54inter7));
  inv1  gate365(.a(N285), .O(gate54inter8));
  nand2 gate366(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate367(.a(s_23), .b(gate54inter3), .O(gate54inter10));
  nor2  gate368(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate369(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate370(.a(gate54inter12), .b(gate54inter1), .O(N319));
xor2 gate55( .a(N286), .b(N287), .O(N320) );

  xor2  gate511(.a(N289), .b(N288), .O(gate56inter0));
  nand2 gate512(.a(gate56inter0), .b(s_44), .O(gate56inter1));
  and2  gate513(.a(N289), .b(N288), .O(gate56inter2));
  inv1  gate514(.a(s_44), .O(gate56inter3));
  inv1  gate515(.a(s_45), .O(gate56inter4));
  nand2 gate516(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate517(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate518(.a(N288), .O(gate56inter7));
  inv1  gate519(.a(N289), .O(gate56inter8));
  nand2 gate520(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate521(.a(s_45), .b(gate56inter3), .O(gate56inter10));
  nor2  gate522(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate523(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate524(.a(gate56inter12), .b(gate56inter1), .O(N321));
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate203(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate204(.a(gate59inter0), .b(s_0), .O(gate59inter1));
  and2  gate205(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate206(.a(s_0), .O(gate59inter3));
  inv1  gate207(.a(s_1), .O(gate59inter4));
  nand2 gate208(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate209(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate210(.a(N290), .O(gate59inter7));
  inv1  gate211(.a(N296), .O(gate59inter8));
  nand2 gate212(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate213(.a(s_1), .b(gate59inter3), .O(gate59inter10));
  nor2  gate214(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate215(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate216(.a(gate59inter12), .b(gate59inter1), .O(N340));
xor2 gate60( .a(N293), .b(N299), .O(N341) );

  xor2  gate385(.a(N305), .b(N302), .O(gate61inter0));
  nand2 gate386(.a(gate61inter0), .b(s_26), .O(gate61inter1));
  and2  gate387(.a(N305), .b(N302), .O(gate61inter2));
  inv1  gate388(.a(s_26), .O(gate61inter3));
  inv1  gate389(.a(s_27), .O(gate61inter4));
  nand2 gate390(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate391(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate392(.a(N302), .O(gate61inter7));
  inv1  gate393(.a(N305), .O(gate61inter8));
  nand2 gate394(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate395(.a(s_27), .b(gate61inter3), .O(gate61inter10));
  nor2  gate396(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate397(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate398(.a(gate61inter12), .b(gate61inter1), .O(N342));
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate287(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate288(.a(gate65inter0), .b(s_12), .O(gate65inter1));
  and2  gate289(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate290(.a(s_12), .O(gate65inter3));
  inv1  gate291(.a(s_13), .O(gate65inter4));
  nand2 gate292(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate293(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate294(.a(N266), .O(gate65inter7));
  inv1  gate295(.a(N342), .O(gate65inter8));
  nand2 gate296(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate297(.a(s_13), .b(gate65inter3), .O(gate65inter10));
  nor2  gate298(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate299(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate300(.a(gate65inter12), .b(gate65inter1), .O(N346));
xor2 gate66( .a(N267), .b(N343), .O(N347) );

  xor2  gate539(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate540(.a(gate67inter0), .b(s_48), .O(gate67inter1));
  and2  gate541(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate542(.a(s_48), .O(gate67inter3));
  inv1  gate543(.a(s_49), .O(gate67inter4));
  nand2 gate544(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate545(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate546(.a(N268), .O(gate67inter7));
  inv1  gate547(.a(N344), .O(gate67inter8));
  nand2 gate548(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate549(.a(s_49), .b(gate67inter3), .O(gate67inter10));
  nor2  gate550(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate551(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate552(.a(gate67inter12), .b(gate67inter1), .O(N348));
xor2 gate68( .a(N269), .b(N345), .O(N349) );

  xor2  gate399(.a(N338), .b(N270), .O(gate69inter0));
  nand2 gate400(.a(gate69inter0), .b(s_28), .O(gate69inter1));
  and2  gate401(.a(N338), .b(N270), .O(gate69inter2));
  inv1  gate402(.a(s_28), .O(gate69inter3));
  inv1  gate403(.a(s_29), .O(gate69inter4));
  nand2 gate404(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate405(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate406(.a(N270), .O(gate69inter7));
  inv1  gate407(.a(N338), .O(gate69inter8));
  nand2 gate408(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate409(.a(s_29), .b(gate69inter3), .O(gate69inter10));
  nor2  gate410(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate411(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate412(.a(gate69inter12), .b(gate69inter1), .O(N350));

  xor2  gate343(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate344(.a(gate70inter0), .b(s_20), .O(gate70inter1));
  and2  gate345(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate346(.a(s_20), .O(gate70inter3));
  inv1  gate347(.a(s_21), .O(gate70inter4));
  nand2 gate348(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate349(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate350(.a(N271), .O(gate70inter7));
  inv1  gate351(.a(N339), .O(gate70inter8));
  nand2 gate352(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate353(.a(s_21), .b(gate70inter3), .O(gate70inter10));
  nor2  gate354(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate355(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate356(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );

  xor2  gate217(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate218(.a(gate74inter0), .b(s_2), .O(gate74inter1));
  and2  gate219(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate220(.a(s_2), .O(gate74inter3));
  inv1  gate221(.a(s_3), .O(gate74inter4));
  nand2 gate222(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate223(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate224(.a(N315), .O(gate74inter7));
  inv1  gate225(.a(N347), .O(gate74inter8));
  nand2 gate226(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate227(.a(s_3), .b(gate74inter3), .O(gate74inter10));
  nor2  gate228(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate229(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate230(.a(gate74inter12), .b(gate74inter1), .O(N367));
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );

  xor2  gate427(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate428(.a(gate77inter0), .b(s_32), .O(gate77inter1));
  and2  gate429(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate430(.a(s_32), .O(gate77inter3));
  inv1  gate431(.a(s_33), .O(gate77inter4));
  nand2 gate432(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate433(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate434(.a(N318), .O(gate77inter7));
  inv1  gate435(.a(N350), .O(gate77inter8));
  nand2 gate436(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate437(.a(s_33), .b(gate77inter3), .O(gate77inter10));
  nor2  gate438(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate439(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate440(.a(gate77inter12), .b(gate77inter1), .O(N406));

  xor2  gate441(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate442(.a(gate78inter0), .b(s_34), .O(gate78inter1));
  and2  gate443(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate444(.a(s_34), .O(gate78inter3));
  inv1  gate445(.a(s_35), .O(gate78inter4));
  nand2 gate446(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate447(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate448(.a(N319), .O(gate78inter7));
  inv1  gate449(.a(N351), .O(gate78inter8));
  nand2 gate450(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate451(.a(s_35), .b(gate78inter3), .O(gate78inter10));
  nor2  gate452(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate453(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate454(.a(gate78inter12), .b(gate78inter1), .O(N419));
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate581(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate582(.a(gate80inter0), .b(s_54), .O(gate80inter1));
  and2  gate583(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate584(.a(s_54), .O(gate80inter3));
  inv1  gate585(.a(s_55), .O(gate80inter4));
  nand2 gate586(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate587(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate588(.a(N321), .O(gate80inter7));
  inv1  gate589(.a(N353), .O(gate80inter8));
  nand2 gate590(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate591(.a(s_55), .b(gate80inter3), .O(gate80inter10));
  nor2  gate592(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate593(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate594(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );

  xor2  gate315(.a(N695), .b(N13), .O(gate174inter0));
  nand2 gate316(.a(gate174inter0), .b(s_16), .O(gate174inter1));
  and2  gate317(.a(N695), .b(N13), .O(gate174inter2));
  inv1  gate318(.a(s_16), .O(gate174inter3));
  inv1  gate319(.a(s_17), .O(gate174inter4));
  nand2 gate320(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate321(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate322(.a(N13), .O(gate174inter7));
  inv1  gate323(.a(N695), .O(gate174inter8));
  nand2 gate324(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate325(.a(s_17), .b(gate174inter3), .O(gate174inter10));
  nor2  gate326(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate327(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate328(.a(gate174inter12), .b(gate174inter1), .O(N727));
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );

  xor2  gate273(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate274(.a(gate178inter0), .b(s_10), .O(gate178inter1));
  and2  gate275(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate276(.a(s_10), .O(gate178inter3));
  inv1  gate277(.a(s_11), .O(gate178inter4));
  nand2 gate278(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate279(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate280(.a(N29), .O(gate178inter7));
  inv1  gate281(.a(N699), .O(gate178inter8));
  nand2 gate282(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate283(.a(s_11), .b(gate178inter3), .O(gate178inter10));
  nor2  gate284(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate285(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate286(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );

  xor2  gate259(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate260(.a(gate182inter0), .b(s_8), .O(gate182inter1));
  and2  gate261(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate262(.a(s_8), .O(gate182inter3));
  inv1  gate263(.a(s_9), .O(gate182inter4));
  nand2 gate264(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate265(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate266(.a(N45), .O(gate182inter7));
  inv1  gate267(.a(N703), .O(gate182inter8));
  nand2 gate268(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate269(.a(s_9), .b(gate182inter3), .O(gate182inter10));
  nor2  gate270(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate271(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate272(.a(gate182inter12), .b(gate182inter1), .O(N735));

  xor2  gate245(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate246(.a(gate183inter0), .b(s_6), .O(gate183inter1));
  and2  gate247(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate248(.a(s_6), .O(gate183inter3));
  inv1  gate249(.a(s_7), .O(gate183inter4));
  nand2 gate250(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate251(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate252(.a(N49), .O(gate183inter7));
  inv1  gate253(.a(N704), .O(gate183inter8));
  nand2 gate254(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate255(.a(s_7), .b(gate183inter3), .O(gate183inter10));
  nor2  gate256(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate257(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate258(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate455(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate456(.a(gate186inter0), .b(s_36), .O(gate186inter1));
  and2  gate457(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate458(.a(s_36), .O(gate186inter3));
  inv1  gate459(.a(s_37), .O(gate186inter4));
  nand2 gate460(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate461(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate462(.a(N61), .O(gate186inter7));
  inv1  gate463(.a(N707), .O(gate186inter8));
  nand2 gate464(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate465(.a(s_37), .b(gate186inter3), .O(gate186inter10));
  nor2  gate466(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate467(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate468(.a(gate186inter12), .b(gate186inter1), .O(N739));
xor2 gate187( .a(N65), .b(N708), .O(N740) );

  xor2  gate231(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate232(.a(gate188inter0), .b(s_4), .O(gate188inter1));
  and2  gate233(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate234(.a(s_4), .O(gate188inter3));
  inv1  gate235(.a(s_5), .O(gate188inter4));
  nand2 gate236(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate237(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate238(.a(N69), .O(gate188inter7));
  inv1  gate239(.a(N709), .O(gate188inter8));
  nand2 gate240(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate241(.a(s_5), .b(gate188inter3), .O(gate188inter10));
  nor2  gate242(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate243(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate244(.a(gate188inter12), .b(gate188inter1), .O(N741));
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );

  xor2  gate469(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate470(.a(gate195inter0), .b(s_38), .O(gate195inter1));
  and2  gate471(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate472(.a(s_38), .O(gate195inter3));
  inv1  gate473(.a(s_39), .O(gate195inter4));
  nand2 gate474(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate475(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate476(.a(N97), .O(gate195inter7));
  inv1  gate477(.a(N716), .O(gate195inter8));
  nand2 gate478(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate479(.a(s_39), .b(gate195inter3), .O(gate195inter10));
  nor2  gate480(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate481(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate482(.a(gate195inter12), .b(gate195inter1), .O(N748));

  xor2  gate623(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate624(.a(gate196inter0), .b(s_60), .O(gate196inter1));
  and2  gate625(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate626(.a(s_60), .O(gate196inter3));
  inv1  gate627(.a(s_61), .O(gate196inter4));
  nand2 gate628(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate629(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate630(.a(N101), .O(gate196inter7));
  inv1  gate631(.a(N717), .O(gate196inter8));
  nand2 gate632(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate633(.a(s_61), .b(gate196inter3), .O(gate196inter10));
  nor2  gate634(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate635(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate636(.a(gate196inter12), .b(gate196inter1), .O(N749));
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );

  xor2  gate413(.a(N721), .b(N117), .O(gate200inter0));
  nand2 gate414(.a(gate200inter0), .b(s_30), .O(gate200inter1));
  and2  gate415(.a(N721), .b(N117), .O(gate200inter2));
  inv1  gate416(.a(s_30), .O(gate200inter3));
  inv1  gate417(.a(s_31), .O(gate200inter4));
  nand2 gate418(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate419(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate420(.a(N117), .O(gate200inter7));
  inv1  gate421(.a(N721), .O(gate200inter8));
  nand2 gate422(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate423(.a(s_31), .b(gate200inter3), .O(gate200inter10));
  nor2  gate424(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate425(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate426(.a(gate200inter12), .b(gate200inter1), .O(N753));

  xor2  gate525(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate526(.a(gate201inter0), .b(s_46), .O(gate201inter1));
  and2  gate527(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate528(.a(s_46), .O(gate201inter3));
  inv1  gate529(.a(s_47), .O(gate201inter4));
  nand2 gate530(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate531(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate532(.a(N121), .O(gate201inter7));
  inv1  gate533(.a(N722), .O(gate201inter8));
  nand2 gate534(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate535(.a(s_47), .b(gate201inter3), .O(gate201inter10));
  nor2  gate536(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate537(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate538(.a(gate201inter12), .b(gate201inter1), .O(N754));

  xor2  gate609(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate610(.a(gate202inter0), .b(s_58), .O(gate202inter1));
  and2  gate611(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate612(.a(s_58), .O(gate202inter3));
  inv1  gate613(.a(s_59), .O(gate202inter4));
  nand2 gate614(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate615(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate616(.a(N125), .O(gate202inter7));
  inv1  gate617(.a(N723), .O(gate202inter8));
  nand2 gate618(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate619(.a(s_59), .b(gate202inter3), .O(gate202inter10));
  nor2  gate620(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate621(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate622(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule