module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2479(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2480(.a(gate13inter0), .b(s_276), .O(gate13inter1));
  and2  gate2481(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2482(.a(s_276), .O(gate13inter3));
  inv1  gate2483(.a(s_277), .O(gate13inter4));
  nand2 gate2484(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2485(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2486(.a(G9), .O(gate13inter7));
  inv1  gate2487(.a(G10), .O(gate13inter8));
  nand2 gate2488(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2489(.a(s_277), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2490(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2491(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2492(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1611(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1612(.a(gate14inter0), .b(s_152), .O(gate14inter1));
  and2  gate1613(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1614(.a(s_152), .O(gate14inter3));
  inv1  gate1615(.a(s_153), .O(gate14inter4));
  nand2 gate1616(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1617(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1618(.a(G11), .O(gate14inter7));
  inv1  gate1619(.a(G12), .O(gate14inter8));
  nand2 gate1620(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1621(.a(s_153), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1622(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1623(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1624(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate743(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate744(.a(gate16inter0), .b(s_28), .O(gate16inter1));
  and2  gate745(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate746(.a(s_28), .O(gate16inter3));
  inv1  gate747(.a(s_29), .O(gate16inter4));
  nand2 gate748(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate749(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate750(.a(G15), .O(gate16inter7));
  inv1  gate751(.a(G16), .O(gate16inter8));
  nand2 gate752(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate753(.a(s_29), .b(gate16inter3), .O(gate16inter10));
  nor2  gate754(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate755(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate756(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2381(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2382(.a(gate19inter0), .b(s_262), .O(gate19inter1));
  and2  gate2383(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2384(.a(s_262), .O(gate19inter3));
  inv1  gate2385(.a(s_263), .O(gate19inter4));
  nand2 gate2386(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2387(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2388(.a(G21), .O(gate19inter7));
  inv1  gate2389(.a(G22), .O(gate19inter8));
  nand2 gate2390(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2391(.a(s_263), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2392(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2393(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2394(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2115(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2116(.a(gate22inter0), .b(s_224), .O(gate22inter1));
  and2  gate2117(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2118(.a(s_224), .O(gate22inter3));
  inv1  gate2119(.a(s_225), .O(gate22inter4));
  nand2 gate2120(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2121(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2122(.a(G27), .O(gate22inter7));
  inv1  gate2123(.a(G28), .O(gate22inter8));
  nand2 gate2124(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2125(.a(s_225), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2126(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2127(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2128(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2283(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2284(.a(gate24inter0), .b(s_248), .O(gate24inter1));
  and2  gate2285(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2286(.a(s_248), .O(gate24inter3));
  inv1  gate2287(.a(s_249), .O(gate24inter4));
  nand2 gate2288(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2289(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2290(.a(G31), .O(gate24inter7));
  inv1  gate2291(.a(G32), .O(gate24inter8));
  nand2 gate2292(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2293(.a(s_249), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2294(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2295(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2296(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1597(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1598(.a(gate25inter0), .b(s_150), .O(gate25inter1));
  and2  gate1599(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1600(.a(s_150), .O(gate25inter3));
  inv1  gate1601(.a(s_151), .O(gate25inter4));
  nand2 gate1602(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1603(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1604(.a(G1), .O(gate25inter7));
  inv1  gate1605(.a(G5), .O(gate25inter8));
  nand2 gate1606(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1607(.a(s_151), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1608(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1609(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1610(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate575(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate576(.a(gate31inter0), .b(s_4), .O(gate31inter1));
  and2  gate577(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate578(.a(s_4), .O(gate31inter3));
  inv1  gate579(.a(s_5), .O(gate31inter4));
  nand2 gate580(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate581(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate582(.a(G4), .O(gate31inter7));
  inv1  gate583(.a(G8), .O(gate31inter8));
  nand2 gate584(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate585(.a(s_5), .b(gate31inter3), .O(gate31inter10));
  nor2  gate586(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate587(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate588(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1275(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1276(.a(gate34inter0), .b(s_104), .O(gate34inter1));
  and2  gate1277(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1278(.a(s_104), .O(gate34inter3));
  inv1  gate1279(.a(s_105), .O(gate34inter4));
  nand2 gate1280(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1281(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1282(.a(G25), .O(gate34inter7));
  inv1  gate1283(.a(G29), .O(gate34inter8));
  nand2 gate1284(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1285(.a(s_105), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1286(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1287(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1288(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1989(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1990(.a(gate36inter0), .b(s_206), .O(gate36inter1));
  and2  gate1991(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1992(.a(s_206), .O(gate36inter3));
  inv1  gate1993(.a(s_207), .O(gate36inter4));
  nand2 gate1994(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1995(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1996(.a(G26), .O(gate36inter7));
  inv1  gate1997(.a(G30), .O(gate36inter8));
  nand2 gate1998(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1999(.a(s_207), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2000(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2001(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2002(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2297(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2298(.a(gate40inter0), .b(s_250), .O(gate40inter1));
  and2  gate2299(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2300(.a(s_250), .O(gate40inter3));
  inv1  gate2301(.a(s_251), .O(gate40inter4));
  nand2 gate2302(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2303(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2304(.a(G28), .O(gate40inter7));
  inv1  gate2305(.a(G32), .O(gate40inter8));
  nand2 gate2306(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2307(.a(s_251), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2308(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2309(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2310(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate939(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate940(.a(gate41inter0), .b(s_56), .O(gate41inter1));
  and2  gate941(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate942(.a(s_56), .O(gate41inter3));
  inv1  gate943(.a(s_57), .O(gate41inter4));
  nand2 gate944(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate945(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate946(.a(G1), .O(gate41inter7));
  inv1  gate947(.a(G266), .O(gate41inter8));
  nand2 gate948(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate949(.a(s_57), .b(gate41inter3), .O(gate41inter10));
  nor2  gate950(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate951(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate952(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1191(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1192(.a(gate44inter0), .b(s_92), .O(gate44inter1));
  and2  gate1193(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1194(.a(s_92), .O(gate44inter3));
  inv1  gate1195(.a(s_93), .O(gate44inter4));
  nand2 gate1196(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1197(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1198(.a(G4), .O(gate44inter7));
  inv1  gate1199(.a(G269), .O(gate44inter8));
  nand2 gate1200(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1201(.a(s_93), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1202(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1203(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1204(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1443(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1444(.a(gate50inter0), .b(s_128), .O(gate50inter1));
  and2  gate1445(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1446(.a(s_128), .O(gate50inter3));
  inv1  gate1447(.a(s_129), .O(gate50inter4));
  nand2 gate1448(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1449(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1450(.a(G10), .O(gate50inter7));
  inv1  gate1451(.a(G278), .O(gate50inter8));
  nand2 gate1452(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1453(.a(s_129), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1454(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1455(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1456(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2129(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2130(.a(gate51inter0), .b(s_226), .O(gate51inter1));
  and2  gate2131(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2132(.a(s_226), .O(gate51inter3));
  inv1  gate2133(.a(s_227), .O(gate51inter4));
  nand2 gate2134(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2135(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2136(.a(G11), .O(gate51inter7));
  inv1  gate2137(.a(G281), .O(gate51inter8));
  nand2 gate2138(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2139(.a(s_227), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2140(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2141(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2142(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1429(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1430(.a(gate54inter0), .b(s_126), .O(gate54inter1));
  and2  gate1431(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1432(.a(s_126), .O(gate54inter3));
  inv1  gate1433(.a(s_127), .O(gate54inter4));
  nand2 gate1434(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1435(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1436(.a(G14), .O(gate54inter7));
  inv1  gate1437(.a(G284), .O(gate54inter8));
  nand2 gate1438(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1439(.a(s_127), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1440(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1441(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1442(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1065(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1066(.a(gate60inter0), .b(s_74), .O(gate60inter1));
  and2  gate1067(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1068(.a(s_74), .O(gate60inter3));
  inv1  gate1069(.a(s_75), .O(gate60inter4));
  nand2 gate1070(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1071(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1072(.a(G20), .O(gate60inter7));
  inv1  gate1073(.a(G293), .O(gate60inter8));
  nand2 gate1074(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1075(.a(s_75), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1076(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1077(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1078(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1177(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1178(.a(gate65inter0), .b(s_90), .O(gate65inter1));
  and2  gate1179(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1180(.a(s_90), .O(gate65inter3));
  inv1  gate1181(.a(s_91), .O(gate65inter4));
  nand2 gate1182(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1183(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1184(.a(G25), .O(gate65inter7));
  inv1  gate1185(.a(G302), .O(gate65inter8));
  nand2 gate1186(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1187(.a(s_91), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1188(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1189(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1190(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate2241(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2242(.a(gate66inter0), .b(s_242), .O(gate66inter1));
  and2  gate2243(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2244(.a(s_242), .O(gate66inter3));
  inv1  gate2245(.a(s_243), .O(gate66inter4));
  nand2 gate2246(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2247(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2248(.a(G26), .O(gate66inter7));
  inv1  gate2249(.a(G302), .O(gate66inter8));
  nand2 gate2250(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2251(.a(s_243), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2252(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2253(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2254(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2451(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2452(.a(gate69inter0), .b(s_272), .O(gate69inter1));
  and2  gate2453(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2454(.a(s_272), .O(gate69inter3));
  inv1  gate2455(.a(s_273), .O(gate69inter4));
  nand2 gate2456(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2457(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2458(.a(G29), .O(gate69inter7));
  inv1  gate2459(.a(G308), .O(gate69inter8));
  nand2 gate2460(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2461(.a(s_273), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2462(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2463(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2464(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate547(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate548(.a(gate72inter0), .b(s_0), .O(gate72inter1));
  and2  gate549(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate550(.a(s_0), .O(gate72inter3));
  inv1  gate551(.a(s_1), .O(gate72inter4));
  nand2 gate552(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate553(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate554(.a(G32), .O(gate72inter7));
  inv1  gate555(.a(G311), .O(gate72inter8));
  nand2 gate556(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate557(.a(s_1), .b(gate72inter3), .O(gate72inter10));
  nor2  gate558(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate559(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate560(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1219(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1220(.a(gate73inter0), .b(s_96), .O(gate73inter1));
  and2  gate1221(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1222(.a(s_96), .O(gate73inter3));
  inv1  gate1223(.a(s_97), .O(gate73inter4));
  nand2 gate1224(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1225(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1226(.a(G1), .O(gate73inter7));
  inv1  gate1227(.a(G314), .O(gate73inter8));
  nand2 gate1228(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1229(.a(s_97), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1230(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1231(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1232(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1723(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1724(.a(gate75inter0), .b(s_168), .O(gate75inter1));
  and2  gate1725(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1726(.a(s_168), .O(gate75inter3));
  inv1  gate1727(.a(s_169), .O(gate75inter4));
  nand2 gate1728(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1729(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1730(.a(G9), .O(gate75inter7));
  inv1  gate1731(.a(G317), .O(gate75inter8));
  nand2 gate1732(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1733(.a(s_169), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1734(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1735(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1736(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1317(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1318(.a(gate76inter0), .b(s_110), .O(gate76inter1));
  and2  gate1319(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1320(.a(s_110), .O(gate76inter3));
  inv1  gate1321(.a(s_111), .O(gate76inter4));
  nand2 gate1322(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1323(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1324(.a(G13), .O(gate76inter7));
  inv1  gate1325(.a(G317), .O(gate76inter8));
  nand2 gate1326(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1327(.a(s_111), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1328(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1329(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1330(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate687(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate688(.a(gate77inter0), .b(s_20), .O(gate77inter1));
  and2  gate689(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate690(.a(s_20), .O(gate77inter3));
  inv1  gate691(.a(s_21), .O(gate77inter4));
  nand2 gate692(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate693(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate694(.a(G2), .O(gate77inter7));
  inv1  gate695(.a(G320), .O(gate77inter8));
  nand2 gate696(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate697(.a(s_21), .b(gate77inter3), .O(gate77inter10));
  nor2  gate698(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate699(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate700(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1205(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1206(.a(gate78inter0), .b(s_94), .O(gate78inter1));
  and2  gate1207(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1208(.a(s_94), .O(gate78inter3));
  inv1  gate1209(.a(s_95), .O(gate78inter4));
  nand2 gate1210(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1211(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1212(.a(G6), .O(gate78inter7));
  inv1  gate1213(.a(G320), .O(gate78inter8));
  nand2 gate1214(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1215(.a(s_95), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1216(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1217(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1218(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2325(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2326(.a(gate85inter0), .b(s_254), .O(gate85inter1));
  and2  gate2327(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2328(.a(s_254), .O(gate85inter3));
  inv1  gate2329(.a(s_255), .O(gate85inter4));
  nand2 gate2330(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2331(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2332(.a(G4), .O(gate85inter7));
  inv1  gate2333(.a(G332), .O(gate85inter8));
  nand2 gate2334(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2335(.a(s_255), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2336(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2337(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2338(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate841(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate842(.a(gate87inter0), .b(s_42), .O(gate87inter1));
  and2  gate843(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate844(.a(s_42), .O(gate87inter3));
  inv1  gate845(.a(s_43), .O(gate87inter4));
  nand2 gate846(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate847(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate848(.a(G12), .O(gate87inter7));
  inv1  gate849(.a(G335), .O(gate87inter8));
  nand2 gate850(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate851(.a(s_43), .b(gate87inter3), .O(gate87inter10));
  nor2  gate852(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate853(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate854(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2507(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2508(.a(gate94inter0), .b(s_280), .O(gate94inter1));
  and2  gate2509(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2510(.a(s_280), .O(gate94inter3));
  inv1  gate2511(.a(s_281), .O(gate94inter4));
  nand2 gate2512(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2513(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2514(.a(G22), .O(gate94inter7));
  inv1  gate2515(.a(G344), .O(gate94inter8));
  nand2 gate2516(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2517(.a(s_281), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2518(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2519(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2520(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1387(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1388(.a(gate95inter0), .b(s_120), .O(gate95inter1));
  and2  gate1389(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1390(.a(s_120), .O(gate95inter3));
  inv1  gate1391(.a(s_121), .O(gate95inter4));
  nand2 gate1392(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1393(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1394(.a(G26), .O(gate95inter7));
  inv1  gate1395(.a(G347), .O(gate95inter8));
  nand2 gate1396(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1397(.a(s_121), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1398(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1399(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1400(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2367(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2368(.a(gate96inter0), .b(s_260), .O(gate96inter1));
  and2  gate2369(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2370(.a(s_260), .O(gate96inter3));
  inv1  gate2371(.a(s_261), .O(gate96inter4));
  nand2 gate2372(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2373(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2374(.a(G30), .O(gate96inter7));
  inv1  gate2375(.a(G347), .O(gate96inter8));
  nand2 gate2376(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2377(.a(s_261), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2378(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2379(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2380(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate673(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate674(.a(gate98inter0), .b(s_18), .O(gate98inter1));
  and2  gate675(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate676(.a(s_18), .O(gate98inter3));
  inv1  gate677(.a(s_19), .O(gate98inter4));
  nand2 gate678(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate679(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate680(.a(G23), .O(gate98inter7));
  inv1  gate681(.a(G350), .O(gate98inter8));
  nand2 gate682(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate683(.a(s_19), .b(gate98inter3), .O(gate98inter10));
  nor2  gate684(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate685(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate686(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1877(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1878(.a(gate99inter0), .b(s_190), .O(gate99inter1));
  and2  gate1879(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1880(.a(s_190), .O(gate99inter3));
  inv1  gate1881(.a(s_191), .O(gate99inter4));
  nand2 gate1882(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1883(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1884(.a(G27), .O(gate99inter7));
  inv1  gate1885(.a(G353), .O(gate99inter8));
  nand2 gate1886(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1887(.a(s_191), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1888(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1889(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1890(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2395(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2396(.a(gate102inter0), .b(s_264), .O(gate102inter1));
  and2  gate2397(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2398(.a(s_264), .O(gate102inter3));
  inv1  gate2399(.a(s_265), .O(gate102inter4));
  nand2 gate2400(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2401(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2402(.a(G24), .O(gate102inter7));
  inv1  gate2403(.a(G356), .O(gate102inter8));
  nand2 gate2404(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2405(.a(s_265), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2406(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2407(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2408(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1037(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1038(.a(gate105inter0), .b(s_70), .O(gate105inter1));
  and2  gate1039(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1040(.a(s_70), .O(gate105inter3));
  inv1  gate1041(.a(s_71), .O(gate105inter4));
  nand2 gate1042(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1043(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1044(.a(G362), .O(gate105inter7));
  inv1  gate1045(.a(G363), .O(gate105inter8));
  nand2 gate1046(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1047(.a(s_71), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1048(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1049(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1050(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate2213(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2214(.a(gate106inter0), .b(s_238), .O(gate106inter1));
  and2  gate2215(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2216(.a(s_238), .O(gate106inter3));
  inv1  gate2217(.a(s_239), .O(gate106inter4));
  nand2 gate2218(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2219(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2220(.a(G364), .O(gate106inter7));
  inv1  gate2221(.a(G365), .O(gate106inter8));
  nand2 gate2222(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2223(.a(s_239), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2224(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2225(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2226(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1457(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1458(.a(gate108inter0), .b(s_130), .O(gate108inter1));
  and2  gate1459(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1460(.a(s_130), .O(gate108inter3));
  inv1  gate1461(.a(s_131), .O(gate108inter4));
  nand2 gate1462(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1463(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1464(.a(G368), .O(gate108inter7));
  inv1  gate1465(.a(G369), .O(gate108inter8));
  nand2 gate1466(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1467(.a(s_131), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1468(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1469(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1470(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1149(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1150(.a(gate112inter0), .b(s_86), .O(gate112inter1));
  and2  gate1151(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1152(.a(s_86), .O(gate112inter3));
  inv1  gate1153(.a(s_87), .O(gate112inter4));
  nand2 gate1154(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1155(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1156(.a(G376), .O(gate112inter7));
  inv1  gate1157(.a(G377), .O(gate112inter8));
  nand2 gate1158(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1159(.a(s_87), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1160(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1161(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1162(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate729(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate730(.a(gate113inter0), .b(s_26), .O(gate113inter1));
  and2  gate731(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate732(.a(s_26), .O(gate113inter3));
  inv1  gate733(.a(s_27), .O(gate113inter4));
  nand2 gate734(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate735(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate736(.a(G378), .O(gate113inter7));
  inv1  gate737(.a(G379), .O(gate113inter8));
  nand2 gate738(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate739(.a(s_27), .b(gate113inter3), .O(gate113inter10));
  nor2  gate740(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate741(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate742(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1905(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1906(.a(gate116inter0), .b(s_194), .O(gate116inter1));
  and2  gate1907(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1908(.a(s_194), .O(gate116inter3));
  inv1  gate1909(.a(s_195), .O(gate116inter4));
  nand2 gate1910(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1911(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1912(.a(G384), .O(gate116inter7));
  inv1  gate1913(.a(G385), .O(gate116inter8));
  nand2 gate1914(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1915(.a(s_195), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1916(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1917(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1918(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2073(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2074(.a(gate120inter0), .b(s_218), .O(gate120inter1));
  and2  gate2075(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2076(.a(s_218), .O(gate120inter3));
  inv1  gate2077(.a(s_219), .O(gate120inter4));
  nand2 gate2078(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2079(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2080(.a(G392), .O(gate120inter7));
  inv1  gate2081(.a(G393), .O(gate120inter8));
  nand2 gate2082(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2083(.a(s_219), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2084(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2085(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2086(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2227(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2228(.a(gate127inter0), .b(s_240), .O(gate127inter1));
  and2  gate2229(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2230(.a(s_240), .O(gate127inter3));
  inv1  gate2231(.a(s_241), .O(gate127inter4));
  nand2 gate2232(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2233(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2234(.a(G406), .O(gate127inter7));
  inv1  gate2235(.a(G407), .O(gate127inter8));
  nand2 gate2236(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2237(.a(s_241), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2238(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2239(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2240(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1051(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1052(.a(gate128inter0), .b(s_72), .O(gate128inter1));
  and2  gate1053(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1054(.a(s_72), .O(gate128inter3));
  inv1  gate1055(.a(s_73), .O(gate128inter4));
  nand2 gate1056(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1057(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1058(.a(G408), .O(gate128inter7));
  inv1  gate1059(.a(G409), .O(gate128inter8));
  nand2 gate1060(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1061(.a(s_73), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1062(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1063(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1064(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2409(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2410(.a(gate129inter0), .b(s_266), .O(gate129inter1));
  and2  gate2411(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2412(.a(s_266), .O(gate129inter3));
  inv1  gate2413(.a(s_267), .O(gate129inter4));
  nand2 gate2414(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2415(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2416(.a(G410), .O(gate129inter7));
  inv1  gate2417(.a(G411), .O(gate129inter8));
  nand2 gate2418(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2419(.a(s_267), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2420(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2421(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2422(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate1975(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1976(.a(gate130inter0), .b(s_204), .O(gate130inter1));
  and2  gate1977(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1978(.a(s_204), .O(gate130inter3));
  inv1  gate1979(.a(s_205), .O(gate130inter4));
  nand2 gate1980(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1981(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1982(.a(G412), .O(gate130inter7));
  inv1  gate1983(.a(G413), .O(gate130inter8));
  nand2 gate1984(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1985(.a(s_205), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1986(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1987(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1988(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1695(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1696(.a(gate131inter0), .b(s_164), .O(gate131inter1));
  and2  gate1697(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1698(.a(s_164), .O(gate131inter3));
  inv1  gate1699(.a(s_165), .O(gate131inter4));
  nand2 gate1700(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1701(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1702(.a(G414), .O(gate131inter7));
  inv1  gate1703(.a(G415), .O(gate131inter8));
  nand2 gate1704(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1705(.a(s_165), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1706(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1707(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1708(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1513(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1514(.a(gate132inter0), .b(s_138), .O(gate132inter1));
  and2  gate1515(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1516(.a(s_138), .O(gate132inter3));
  inv1  gate1517(.a(s_139), .O(gate132inter4));
  nand2 gate1518(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1519(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1520(.a(G416), .O(gate132inter7));
  inv1  gate1521(.a(G417), .O(gate132inter8));
  nand2 gate1522(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1523(.a(s_139), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1524(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1525(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1526(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1359(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1360(.a(gate134inter0), .b(s_116), .O(gate134inter1));
  and2  gate1361(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1362(.a(s_116), .O(gate134inter3));
  inv1  gate1363(.a(s_117), .O(gate134inter4));
  nand2 gate1364(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1365(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1366(.a(G420), .O(gate134inter7));
  inv1  gate1367(.a(G421), .O(gate134inter8));
  nand2 gate1368(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1369(.a(s_117), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1370(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1371(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1372(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate715(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate716(.a(gate139inter0), .b(s_24), .O(gate139inter1));
  and2  gate717(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate718(.a(s_24), .O(gate139inter3));
  inv1  gate719(.a(s_25), .O(gate139inter4));
  nand2 gate720(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate721(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate722(.a(G438), .O(gate139inter7));
  inv1  gate723(.a(G441), .O(gate139inter8));
  nand2 gate724(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate725(.a(s_25), .b(gate139inter3), .O(gate139inter10));
  nor2  gate726(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate727(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate728(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate2171(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2172(.a(gate141inter0), .b(s_232), .O(gate141inter1));
  and2  gate2173(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2174(.a(s_232), .O(gate141inter3));
  inv1  gate2175(.a(s_233), .O(gate141inter4));
  nand2 gate2176(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2177(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2178(.a(G450), .O(gate141inter7));
  inv1  gate2179(.a(G453), .O(gate141inter8));
  nand2 gate2180(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2181(.a(s_233), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2182(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2183(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2184(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate1289(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1290(.a(gate142inter0), .b(s_106), .O(gate142inter1));
  and2  gate1291(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1292(.a(s_106), .O(gate142inter3));
  inv1  gate1293(.a(s_107), .O(gate142inter4));
  nand2 gate1294(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1295(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1296(.a(G456), .O(gate142inter7));
  inv1  gate1297(.a(G459), .O(gate142inter8));
  nand2 gate1298(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1299(.a(s_107), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1300(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1301(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1302(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1079(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1080(.a(gate147inter0), .b(s_76), .O(gate147inter1));
  and2  gate1081(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1082(.a(s_76), .O(gate147inter3));
  inv1  gate1083(.a(s_77), .O(gate147inter4));
  nand2 gate1084(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1085(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1086(.a(G486), .O(gate147inter7));
  inv1  gate1087(.a(G489), .O(gate147inter8));
  nand2 gate1088(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1089(.a(s_77), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1090(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1091(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1092(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1625(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1626(.a(gate149inter0), .b(s_154), .O(gate149inter1));
  and2  gate1627(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1628(.a(s_154), .O(gate149inter3));
  inv1  gate1629(.a(s_155), .O(gate149inter4));
  nand2 gate1630(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1631(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1632(.a(G498), .O(gate149inter7));
  inv1  gate1633(.a(G501), .O(gate149inter8));
  nand2 gate1634(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1635(.a(s_155), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1636(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1637(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1638(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2003(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2004(.a(gate153inter0), .b(s_208), .O(gate153inter1));
  and2  gate2005(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2006(.a(s_208), .O(gate153inter3));
  inv1  gate2007(.a(s_209), .O(gate153inter4));
  nand2 gate2008(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2009(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2010(.a(G426), .O(gate153inter7));
  inv1  gate2011(.a(G522), .O(gate153inter8));
  nand2 gate2012(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2013(.a(s_209), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2014(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2015(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2016(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1107(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1108(.a(gate157inter0), .b(s_80), .O(gate157inter1));
  and2  gate1109(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1110(.a(s_80), .O(gate157inter3));
  inv1  gate1111(.a(s_81), .O(gate157inter4));
  nand2 gate1112(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1113(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1114(.a(G438), .O(gate157inter7));
  inv1  gate1115(.a(G528), .O(gate157inter8));
  nand2 gate1116(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1117(.a(s_81), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1118(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1119(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1120(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate827(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate828(.a(gate158inter0), .b(s_40), .O(gate158inter1));
  and2  gate829(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate830(.a(s_40), .O(gate158inter3));
  inv1  gate831(.a(s_41), .O(gate158inter4));
  nand2 gate832(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate833(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate834(.a(G441), .O(gate158inter7));
  inv1  gate835(.a(G528), .O(gate158inter8));
  nand2 gate836(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate837(.a(s_41), .b(gate158inter3), .O(gate158inter10));
  nor2  gate838(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate839(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate840(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1583(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1584(.a(gate159inter0), .b(s_148), .O(gate159inter1));
  and2  gate1585(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1586(.a(s_148), .O(gate159inter3));
  inv1  gate1587(.a(s_149), .O(gate159inter4));
  nand2 gate1588(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1589(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1590(.a(G444), .O(gate159inter7));
  inv1  gate1591(.a(G531), .O(gate159inter8));
  nand2 gate1592(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1593(.a(s_149), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1594(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1595(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1596(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2101(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2102(.a(gate161inter0), .b(s_222), .O(gate161inter1));
  and2  gate2103(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2104(.a(s_222), .O(gate161inter3));
  inv1  gate2105(.a(s_223), .O(gate161inter4));
  nand2 gate2106(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2107(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2108(.a(G450), .O(gate161inter7));
  inv1  gate2109(.a(G534), .O(gate161inter8));
  nand2 gate2110(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2111(.a(s_223), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2112(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2113(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2114(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate757(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate758(.a(gate162inter0), .b(s_30), .O(gate162inter1));
  and2  gate759(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate760(.a(s_30), .O(gate162inter3));
  inv1  gate761(.a(s_31), .O(gate162inter4));
  nand2 gate762(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate763(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate764(.a(G453), .O(gate162inter7));
  inv1  gate765(.a(G534), .O(gate162inter8));
  nand2 gate766(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate767(.a(s_31), .b(gate162inter3), .O(gate162inter10));
  nor2  gate768(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate769(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate770(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate701(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate702(.a(gate165inter0), .b(s_22), .O(gate165inter1));
  and2  gate703(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate704(.a(s_22), .O(gate165inter3));
  inv1  gate705(.a(s_23), .O(gate165inter4));
  nand2 gate706(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate707(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate708(.a(G462), .O(gate165inter7));
  inv1  gate709(.a(G540), .O(gate165inter8));
  nand2 gate710(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate711(.a(s_23), .b(gate165inter3), .O(gate165inter10));
  nor2  gate712(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate713(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate714(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2311(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2312(.a(gate171inter0), .b(s_252), .O(gate171inter1));
  and2  gate2313(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2314(.a(s_252), .O(gate171inter3));
  inv1  gate2315(.a(s_253), .O(gate171inter4));
  nand2 gate2316(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2317(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2318(.a(G480), .O(gate171inter7));
  inv1  gate2319(.a(G549), .O(gate171inter8));
  nand2 gate2320(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2321(.a(s_253), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2322(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2323(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2324(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2059(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2060(.a(gate172inter0), .b(s_216), .O(gate172inter1));
  and2  gate2061(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2062(.a(s_216), .O(gate172inter3));
  inv1  gate2063(.a(s_217), .O(gate172inter4));
  nand2 gate2064(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2065(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2066(.a(G483), .O(gate172inter7));
  inv1  gate2067(.a(G549), .O(gate172inter8));
  nand2 gate2068(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2069(.a(s_217), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2070(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2071(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2072(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1639(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1640(.a(gate175inter0), .b(s_156), .O(gate175inter1));
  and2  gate1641(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1642(.a(s_156), .O(gate175inter3));
  inv1  gate1643(.a(s_157), .O(gate175inter4));
  nand2 gate1644(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1645(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1646(.a(G492), .O(gate175inter7));
  inv1  gate1647(.a(G555), .O(gate175inter8));
  nand2 gate1648(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1649(.a(s_157), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1650(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1651(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1652(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1835(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1836(.a(gate176inter0), .b(s_184), .O(gate176inter1));
  and2  gate1837(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1838(.a(s_184), .O(gate176inter3));
  inv1  gate1839(.a(s_185), .O(gate176inter4));
  nand2 gate1840(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1841(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1842(.a(G495), .O(gate176inter7));
  inv1  gate1843(.a(G555), .O(gate176inter8));
  nand2 gate1844(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1845(.a(s_185), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1846(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1847(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1848(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1373(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1374(.a(gate179inter0), .b(s_118), .O(gate179inter1));
  and2  gate1375(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1376(.a(s_118), .O(gate179inter3));
  inv1  gate1377(.a(s_119), .O(gate179inter4));
  nand2 gate1378(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1379(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1380(.a(G504), .O(gate179inter7));
  inv1  gate1381(.a(G561), .O(gate179inter8));
  nand2 gate1382(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1383(.a(s_119), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1384(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1385(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1386(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate953(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate954(.a(gate187inter0), .b(s_58), .O(gate187inter1));
  and2  gate955(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate956(.a(s_58), .O(gate187inter3));
  inv1  gate957(.a(s_59), .O(gate187inter4));
  nand2 gate958(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate959(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate960(.a(G574), .O(gate187inter7));
  inv1  gate961(.a(G575), .O(gate187inter8));
  nand2 gate962(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate963(.a(s_59), .b(gate187inter3), .O(gate187inter10));
  nor2  gate964(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate965(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate966(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate967(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate968(.a(gate193inter0), .b(s_60), .O(gate193inter1));
  and2  gate969(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate970(.a(s_60), .O(gate193inter3));
  inv1  gate971(.a(s_61), .O(gate193inter4));
  nand2 gate972(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate973(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate974(.a(G586), .O(gate193inter7));
  inv1  gate975(.a(G587), .O(gate193inter8));
  nand2 gate976(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate977(.a(s_61), .b(gate193inter3), .O(gate193inter10));
  nor2  gate978(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate979(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate980(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate603(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate604(.a(gate195inter0), .b(s_8), .O(gate195inter1));
  and2  gate605(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate606(.a(s_8), .O(gate195inter3));
  inv1  gate607(.a(s_9), .O(gate195inter4));
  nand2 gate608(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate609(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate610(.a(G590), .O(gate195inter7));
  inv1  gate611(.a(G591), .O(gate195inter8));
  nand2 gate612(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate613(.a(s_9), .b(gate195inter3), .O(gate195inter10));
  nor2  gate614(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate615(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate616(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2339(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2340(.a(gate196inter0), .b(s_256), .O(gate196inter1));
  and2  gate2341(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2342(.a(s_256), .O(gate196inter3));
  inv1  gate2343(.a(s_257), .O(gate196inter4));
  nand2 gate2344(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2345(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2346(.a(G592), .O(gate196inter7));
  inv1  gate2347(.a(G593), .O(gate196inter8));
  nand2 gate2348(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2349(.a(s_257), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2350(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2351(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2352(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2199(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2200(.a(gate202inter0), .b(s_236), .O(gate202inter1));
  and2  gate2201(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2202(.a(s_236), .O(gate202inter3));
  inv1  gate2203(.a(s_237), .O(gate202inter4));
  nand2 gate2204(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2205(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2206(.a(G612), .O(gate202inter7));
  inv1  gate2207(.a(G617), .O(gate202inter8));
  nand2 gate2208(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2209(.a(s_237), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2210(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2211(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2212(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1793(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1794(.a(gate208inter0), .b(s_178), .O(gate208inter1));
  and2  gate1795(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1796(.a(s_178), .O(gate208inter3));
  inv1  gate1797(.a(s_179), .O(gate208inter4));
  nand2 gate1798(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1799(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1800(.a(G627), .O(gate208inter7));
  inv1  gate1801(.a(G637), .O(gate208inter8));
  nand2 gate1802(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1803(.a(s_179), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1804(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1805(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1806(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1961(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1962(.a(gate210inter0), .b(s_202), .O(gate210inter1));
  and2  gate1963(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1964(.a(s_202), .O(gate210inter3));
  inv1  gate1965(.a(s_203), .O(gate210inter4));
  nand2 gate1966(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1967(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1968(.a(G607), .O(gate210inter7));
  inv1  gate1969(.a(G666), .O(gate210inter8));
  nand2 gate1970(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1971(.a(s_203), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1972(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1973(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1974(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2185(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2186(.a(gate222inter0), .b(s_234), .O(gate222inter1));
  and2  gate2187(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2188(.a(s_234), .O(gate222inter3));
  inv1  gate2189(.a(s_235), .O(gate222inter4));
  nand2 gate2190(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2191(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2192(.a(G632), .O(gate222inter7));
  inv1  gate2193(.a(G684), .O(gate222inter8));
  nand2 gate2194(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2195(.a(s_235), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2196(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2197(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2198(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate659(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate660(.a(gate224inter0), .b(s_16), .O(gate224inter1));
  and2  gate661(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate662(.a(s_16), .O(gate224inter3));
  inv1  gate663(.a(s_17), .O(gate224inter4));
  nand2 gate664(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate665(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate666(.a(G637), .O(gate224inter7));
  inv1  gate667(.a(G687), .O(gate224inter8));
  nand2 gate668(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate669(.a(s_17), .b(gate224inter3), .O(gate224inter10));
  nor2  gate670(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate671(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate672(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate2087(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2088(.a(gate225inter0), .b(s_220), .O(gate225inter1));
  and2  gate2089(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2090(.a(s_220), .O(gate225inter3));
  inv1  gate2091(.a(s_221), .O(gate225inter4));
  nand2 gate2092(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2093(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2094(.a(G690), .O(gate225inter7));
  inv1  gate2095(.a(G691), .O(gate225inter8));
  nand2 gate2096(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2097(.a(s_221), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2098(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2099(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2100(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate911(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate912(.a(gate226inter0), .b(s_52), .O(gate226inter1));
  and2  gate913(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate914(.a(s_52), .O(gate226inter3));
  inv1  gate915(.a(s_53), .O(gate226inter4));
  nand2 gate916(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate917(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate918(.a(G692), .O(gate226inter7));
  inv1  gate919(.a(G693), .O(gate226inter8));
  nand2 gate920(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate921(.a(s_53), .b(gate226inter3), .O(gate226inter10));
  nor2  gate922(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate923(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate924(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate869(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate870(.a(gate229inter0), .b(s_46), .O(gate229inter1));
  and2  gate871(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate872(.a(s_46), .O(gate229inter3));
  inv1  gate873(.a(s_47), .O(gate229inter4));
  nand2 gate874(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate875(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate876(.a(G698), .O(gate229inter7));
  inv1  gate877(.a(G699), .O(gate229inter8));
  nand2 gate878(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate879(.a(s_47), .b(gate229inter3), .O(gate229inter10));
  nor2  gate880(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate881(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate882(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1401(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1402(.a(gate233inter0), .b(s_122), .O(gate233inter1));
  and2  gate1403(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1404(.a(s_122), .O(gate233inter3));
  inv1  gate1405(.a(s_123), .O(gate233inter4));
  nand2 gate1406(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1407(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1408(.a(G242), .O(gate233inter7));
  inv1  gate1409(.a(G718), .O(gate233inter8));
  nand2 gate1410(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1411(.a(s_123), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1412(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1413(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1414(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate981(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate982(.a(gate235inter0), .b(s_62), .O(gate235inter1));
  and2  gate983(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate984(.a(s_62), .O(gate235inter3));
  inv1  gate985(.a(s_63), .O(gate235inter4));
  nand2 gate986(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate987(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate988(.a(G248), .O(gate235inter7));
  inv1  gate989(.a(G724), .O(gate235inter8));
  nand2 gate990(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate991(.a(s_63), .b(gate235inter3), .O(gate235inter10));
  nor2  gate992(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate993(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate994(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate561(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate562(.a(gate242inter0), .b(s_2), .O(gate242inter1));
  and2  gate563(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate564(.a(s_2), .O(gate242inter3));
  inv1  gate565(.a(s_3), .O(gate242inter4));
  nand2 gate566(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate567(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate568(.a(G718), .O(gate242inter7));
  inv1  gate569(.a(G730), .O(gate242inter8));
  nand2 gate570(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate571(.a(s_3), .b(gate242inter3), .O(gate242inter10));
  nor2  gate572(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate573(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate574(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1933(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1934(.a(gate243inter0), .b(s_198), .O(gate243inter1));
  and2  gate1935(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1936(.a(s_198), .O(gate243inter3));
  inv1  gate1937(.a(s_199), .O(gate243inter4));
  nand2 gate1938(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1939(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1940(.a(G245), .O(gate243inter7));
  inv1  gate1941(.a(G733), .O(gate243inter8));
  nand2 gate1942(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1943(.a(s_199), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1944(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1945(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1946(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2143(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2144(.a(gate245inter0), .b(s_228), .O(gate245inter1));
  and2  gate2145(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2146(.a(s_228), .O(gate245inter3));
  inv1  gate2147(.a(s_229), .O(gate245inter4));
  nand2 gate2148(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2149(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2150(.a(G248), .O(gate245inter7));
  inv1  gate2151(.a(G736), .O(gate245inter8));
  nand2 gate2152(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2153(.a(s_229), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2154(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2155(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2156(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2353(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2354(.a(gate246inter0), .b(s_258), .O(gate246inter1));
  and2  gate2355(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2356(.a(s_258), .O(gate246inter3));
  inv1  gate2357(.a(s_259), .O(gate246inter4));
  nand2 gate2358(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2359(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2360(.a(G724), .O(gate246inter7));
  inv1  gate2361(.a(G736), .O(gate246inter8));
  nand2 gate2362(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2363(.a(s_259), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2364(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2365(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2366(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2465(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2466(.a(gate248inter0), .b(s_274), .O(gate248inter1));
  and2  gate2467(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2468(.a(s_274), .O(gate248inter3));
  inv1  gate2469(.a(s_275), .O(gate248inter4));
  nand2 gate2470(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2471(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2472(.a(G727), .O(gate248inter7));
  inv1  gate2473(.a(G739), .O(gate248inter8));
  nand2 gate2474(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2475(.a(s_275), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2476(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2477(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2478(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1163(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1164(.a(gate249inter0), .b(s_88), .O(gate249inter1));
  and2  gate1165(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1166(.a(s_88), .O(gate249inter3));
  inv1  gate1167(.a(s_89), .O(gate249inter4));
  nand2 gate1168(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1169(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1170(.a(G254), .O(gate249inter7));
  inv1  gate1171(.a(G742), .O(gate249inter8));
  nand2 gate1172(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1173(.a(s_89), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1174(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1175(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1176(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate589(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate590(.a(gate252inter0), .b(s_6), .O(gate252inter1));
  and2  gate591(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate592(.a(s_6), .O(gate252inter3));
  inv1  gate593(.a(s_7), .O(gate252inter4));
  nand2 gate594(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate595(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate596(.a(G709), .O(gate252inter7));
  inv1  gate597(.a(G745), .O(gate252inter8));
  nand2 gate598(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate599(.a(s_7), .b(gate252inter3), .O(gate252inter10));
  nor2  gate600(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate601(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate602(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate785(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate786(.a(gate253inter0), .b(s_34), .O(gate253inter1));
  and2  gate787(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate788(.a(s_34), .O(gate253inter3));
  inv1  gate789(.a(s_35), .O(gate253inter4));
  nand2 gate790(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate791(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate792(.a(G260), .O(gate253inter7));
  inv1  gate793(.a(G748), .O(gate253inter8));
  nand2 gate794(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate795(.a(s_35), .b(gate253inter3), .O(gate253inter10));
  nor2  gate796(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate797(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate798(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate645(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate646(.a(gate256inter0), .b(s_14), .O(gate256inter1));
  and2  gate647(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate648(.a(s_14), .O(gate256inter3));
  inv1  gate649(.a(s_15), .O(gate256inter4));
  nand2 gate650(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate651(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate652(.a(G715), .O(gate256inter7));
  inv1  gate653(.a(G751), .O(gate256inter8));
  nand2 gate654(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate655(.a(s_15), .b(gate256inter3), .O(gate256inter10));
  nor2  gate656(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate657(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate658(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1135(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1136(.a(gate257inter0), .b(s_84), .O(gate257inter1));
  and2  gate1137(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1138(.a(s_84), .O(gate257inter3));
  inv1  gate1139(.a(s_85), .O(gate257inter4));
  nand2 gate1140(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1141(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1142(.a(G754), .O(gate257inter7));
  inv1  gate1143(.a(G755), .O(gate257inter8));
  nand2 gate1144(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1145(.a(s_85), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1146(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1147(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1148(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate771(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate772(.a(gate262inter0), .b(s_32), .O(gate262inter1));
  and2  gate773(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate774(.a(s_32), .O(gate262inter3));
  inv1  gate775(.a(s_33), .O(gate262inter4));
  nand2 gate776(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate777(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate778(.a(G764), .O(gate262inter7));
  inv1  gate779(.a(G765), .O(gate262inter8));
  nand2 gate780(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate781(.a(s_33), .b(gate262inter3), .O(gate262inter10));
  nor2  gate782(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate783(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate784(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate813(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate814(.a(gate265inter0), .b(s_38), .O(gate265inter1));
  and2  gate815(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate816(.a(s_38), .O(gate265inter3));
  inv1  gate817(.a(s_39), .O(gate265inter4));
  nand2 gate818(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate819(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate820(.a(G642), .O(gate265inter7));
  inv1  gate821(.a(G770), .O(gate265inter8));
  nand2 gate822(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate823(.a(s_39), .b(gate265inter3), .O(gate265inter10));
  nor2  gate824(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate825(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate826(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate617(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate618(.a(gate269inter0), .b(s_10), .O(gate269inter1));
  and2  gate619(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate620(.a(s_10), .O(gate269inter3));
  inv1  gate621(.a(s_11), .O(gate269inter4));
  nand2 gate622(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate623(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate624(.a(G654), .O(gate269inter7));
  inv1  gate625(.a(G782), .O(gate269inter8));
  nand2 gate626(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate627(.a(s_11), .b(gate269inter3), .O(gate269inter10));
  nor2  gate628(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate629(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate630(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1233(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1234(.a(gate272inter0), .b(s_98), .O(gate272inter1));
  and2  gate1235(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1236(.a(s_98), .O(gate272inter3));
  inv1  gate1237(.a(s_99), .O(gate272inter4));
  nand2 gate1238(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1239(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1240(.a(G663), .O(gate272inter7));
  inv1  gate1241(.a(G791), .O(gate272inter8));
  nand2 gate1242(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1243(.a(s_99), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1244(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1245(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1246(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1765(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1766(.a(gate275inter0), .b(s_174), .O(gate275inter1));
  and2  gate1767(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1768(.a(s_174), .O(gate275inter3));
  inv1  gate1769(.a(s_175), .O(gate275inter4));
  nand2 gate1770(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1771(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1772(.a(G645), .O(gate275inter7));
  inv1  gate1773(.a(G797), .O(gate275inter8));
  nand2 gate1774(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1775(.a(s_175), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1776(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1777(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1778(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate995(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate996(.a(gate276inter0), .b(s_64), .O(gate276inter1));
  and2  gate997(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate998(.a(s_64), .O(gate276inter3));
  inv1  gate999(.a(s_65), .O(gate276inter4));
  nand2 gate1000(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1001(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1002(.a(G773), .O(gate276inter7));
  inv1  gate1003(.a(G797), .O(gate276inter8));
  nand2 gate1004(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1005(.a(s_65), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1006(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1007(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1008(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1541(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1542(.a(gate278inter0), .b(s_142), .O(gate278inter1));
  and2  gate1543(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1544(.a(s_142), .O(gate278inter3));
  inv1  gate1545(.a(s_143), .O(gate278inter4));
  nand2 gate1546(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1547(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1548(.a(G776), .O(gate278inter7));
  inv1  gate1549(.a(G800), .O(gate278inter8));
  nand2 gate1550(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1551(.a(s_143), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1552(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1553(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1554(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1891(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1892(.a(gate280inter0), .b(s_192), .O(gate280inter1));
  and2  gate1893(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1894(.a(s_192), .O(gate280inter3));
  inv1  gate1895(.a(s_193), .O(gate280inter4));
  nand2 gate1896(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1897(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1898(.a(G779), .O(gate280inter7));
  inv1  gate1899(.a(G803), .O(gate280inter8));
  nand2 gate1900(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1901(.a(s_193), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1902(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1903(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1904(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1471(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1472(.a(gate285inter0), .b(s_132), .O(gate285inter1));
  and2  gate1473(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1474(.a(s_132), .O(gate285inter3));
  inv1  gate1475(.a(s_133), .O(gate285inter4));
  nand2 gate1476(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1477(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1478(.a(G660), .O(gate285inter7));
  inv1  gate1479(.a(G812), .O(gate285inter8));
  nand2 gate1480(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1481(.a(s_133), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1482(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1483(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1484(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1121(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1122(.a(gate286inter0), .b(s_82), .O(gate286inter1));
  and2  gate1123(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1124(.a(s_82), .O(gate286inter3));
  inv1  gate1125(.a(s_83), .O(gate286inter4));
  nand2 gate1126(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1127(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1128(.a(G788), .O(gate286inter7));
  inv1  gate1129(.a(G812), .O(gate286inter8));
  nand2 gate1130(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1131(.a(s_83), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1132(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1133(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1134(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1947(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1948(.a(gate288inter0), .b(s_200), .O(gate288inter1));
  and2  gate1949(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1950(.a(s_200), .O(gate288inter3));
  inv1  gate1951(.a(s_201), .O(gate288inter4));
  nand2 gate1952(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1953(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1954(.a(G791), .O(gate288inter7));
  inv1  gate1955(.a(G815), .O(gate288inter8));
  nand2 gate1956(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1957(.a(s_201), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1958(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1959(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1960(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1667(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1668(.a(gate293inter0), .b(s_160), .O(gate293inter1));
  and2  gate1669(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1670(.a(s_160), .O(gate293inter3));
  inv1  gate1671(.a(s_161), .O(gate293inter4));
  nand2 gate1672(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1673(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1674(.a(G828), .O(gate293inter7));
  inv1  gate1675(.a(G829), .O(gate293inter8));
  nand2 gate1676(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1677(.a(s_161), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1678(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1679(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1680(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate799(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate800(.a(gate294inter0), .b(s_36), .O(gate294inter1));
  and2  gate801(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate802(.a(s_36), .O(gate294inter3));
  inv1  gate803(.a(s_37), .O(gate294inter4));
  nand2 gate804(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate805(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate806(.a(G832), .O(gate294inter7));
  inv1  gate807(.a(G833), .O(gate294inter8));
  nand2 gate808(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate809(.a(s_37), .b(gate294inter3), .O(gate294inter10));
  nor2  gate810(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate811(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate812(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1919(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1920(.a(gate296inter0), .b(s_196), .O(gate296inter1));
  and2  gate1921(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1922(.a(s_196), .O(gate296inter3));
  inv1  gate1923(.a(s_197), .O(gate296inter4));
  nand2 gate1924(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1925(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1926(.a(G826), .O(gate296inter7));
  inv1  gate1927(.a(G827), .O(gate296inter8));
  nand2 gate1928(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1929(.a(s_197), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1930(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1931(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1932(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1779(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1780(.a(gate391inter0), .b(s_176), .O(gate391inter1));
  and2  gate1781(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1782(.a(s_176), .O(gate391inter3));
  inv1  gate1783(.a(s_177), .O(gate391inter4));
  nand2 gate1784(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1785(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1786(.a(G5), .O(gate391inter7));
  inv1  gate1787(.a(G1048), .O(gate391inter8));
  nand2 gate1788(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1789(.a(s_177), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1790(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1791(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1792(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1303(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1304(.a(gate395inter0), .b(s_108), .O(gate395inter1));
  and2  gate1305(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1306(.a(s_108), .O(gate395inter3));
  inv1  gate1307(.a(s_109), .O(gate395inter4));
  nand2 gate1308(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1309(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1310(.a(G9), .O(gate395inter7));
  inv1  gate1311(.a(G1060), .O(gate395inter8));
  nand2 gate1312(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1313(.a(s_109), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1314(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1315(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1316(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1261(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1262(.a(gate402inter0), .b(s_102), .O(gate402inter1));
  and2  gate1263(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1264(.a(s_102), .O(gate402inter3));
  inv1  gate1265(.a(s_103), .O(gate402inter4));
  nand2 gate1266(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1267(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1268(.a(G16), .O(gate402inter7));
  inv1  gate1269(.a(G1081), .O(gate402inter8));
  nand2 gate1270(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1271(.a(s_103), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1272(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1273(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1274(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1737(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1738(.a(gate404inter0), .b(s_170), .O(gate404inter1));
  and2  gate1739(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1740(.a(s_170), .O(gate404inter3));
  inv1  gate1741(.a(s_171), .O(gate404inter4));
  nand2 gate1742(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1743(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1744(.a(G18), .O(gate404inter7));
  inv1  gate1745(.a(G1087), .O(gate404inter8));
  nand2 gate1746(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1747(.a(s_171), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1748(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1749(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1750(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2157(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2158(.a(gate406inter0), .b(s_230), .O(gate406inter1));
  and2  gate2159(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2160(.a(s_230), .O(gate406inter3));
  inv1  gate2161(.a(s_231), .O(gate406inter4));
  nand2 gate2162(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2163(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2164(.a(G20), .O(gate406inter7));
  inv1  gate2165(.a(G1093), .O(gate406inter8));
  nand2 gate2166(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2167(.a(s_231), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2168(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2169(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2170(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1331(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1332(.a(gate409inter0), .b(s_112), .O(gate409inter1));
  and2  gate1333(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1334(.a(s_112), .O(gate409inter3));
  inv1  gate1335(.a(s_113), .O(gate409inter4));
  nand2 gate1336(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1337(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1338(.a(G23), .O(gate409inter7));
  inv1  gate1339(.a(G1102), .O(gate409inter8));
  nand2 gate1340(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1341(.a(s_113), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1342(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1343(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1344(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1681(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1682(.a(gate424inter0), .b(s_162), .O(gate424inter1));
  and2  gate1683(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1684(.a(s_162), .O(gate424inter3));
  inv1  gate1685(.a(s_163), .O(gate424inter4));
  nand2 gate1686(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1687(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1688(.a(G1042), .O(gate424inter7));
  inv1  gate1689(.a(G1138), .O(gate424inter8));
  nand2 gate1690(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1691(.a(s_163), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1692(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1693(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1694(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1499(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1500(.a(gate426inter0), .b(s_136), .O(gate426inter1));
  and2  gate1501(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1502(.a(s_136), .O(gate426inter3));
  inv1  gate1503(.a(s_137), .O(gate426inter4));
  nand2 gate1504(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1505(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1506(.a(G1045), .O(gate426inter7));
  inv1  gate1507(.a(G1141), .O(gate426inter8));
  nand2 gate1508(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1509(.a(s_137), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1510(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1511(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1512(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2423(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2424(.a(gate428inter0), .b(s_268), .O(gate428inter1));
  and2  gate2425(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2426(.a(s_268), .O(gate428inter3));
  inv1  gate2427(.a(s_269), .O(gate428inter4));
  nand2 gate2428(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2429(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2430(.a(G1048), .O(gate428inter7));
  inv1  gate2431(.a(G1144), .O(gate428inter8));
  nand2 gate2432(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2433(.a(s_269), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2434(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2435(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2436(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1569(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1570(.a(gate432inter0), .b(s_146), .O(gate432inter1));
  and2  gate1571(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1572(.a(s_146), .O(gate432inter3));
  inv1  gate1573(.a(s_147), .O(gate432inter4));
  nand2 gate1574(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1575(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1576(.a(G1054), .O(gate432inter7));
  inv1  gate1577(.a(G1150), .O(gate432inter8));
  nand2 gate1578(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1579(.a(s_147), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1580(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1581(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1582(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2437(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2438(.a(gate442inter0), .b(s_270), .O(gate442inter1));
  and2  gate2439(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2440(.a(s_270), .O(gate442inter3));
  inv1  gate2441(.a(s_271), .O(gate442inter4));
  nand2 gate2442(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2443(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2444(.a(G1069), .O(gate442inter7));
  inv1  gate2445(.a(G1165), .O(gate442inter8));
  nand2 gate2446(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2447(.a(s_271), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2448(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2449(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2450(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1527(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1528(.a(gate448inter0), .b(s_140), .O(gate448inter1));
  and2  gate1529(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1530(.a(s_140), .O(gate448inter3));
  inv1  gate1531(.a(s_141), .O(gate448inter4));
  nand2 gate1532(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1533(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1534(.a(G1078), .O(gate448inter7));
  inv1  gate1535(.a(G1174), .O(gate448inter8));
  nand2 gate1536(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1537(.a(s_141), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1538(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1539(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1540(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1023(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1024(.a(gate449inter0), .b(s_68), .O(gate449inter1));
  and2  gate1025(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1026(.a(s_68), .O(gate449inter3));
  inv1  gate1027(.a(s_69), .O(gate449inter4));
  nand2 gate1028(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1029(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1030(.a(G16), .O(gate449inter7));
  inv1  gate1031(.a(G1177), .O(gate449inter8));
  nand2 gate1032(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1033(.a(s_69), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1034(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1035(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1036(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1345(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1346(.a(gate457inter0), .b(s_114), .O(gate457inter1));
  and2  gate1347(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1348(.a(s_114), .O(gate457inter3));
  inv1  gate1349(.a(s_115), .O(gate457inter4));
  nand2 gate1350(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1351(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1352(.a(G20), .O(gate457inter7));
  inv1  gate1353(.a(G1189), .O(gate457inter8));
  nand2 gate1354(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1355(.a(s_115), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1356(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1357(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1358(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate925(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate926(.a(gate459inter0), .b(s_54), .O(gate459inter1));
  and2  gate927(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate928(.a(s_54), .O(gate459inter3));
  inv1  gate929(.a(s_55), .O(gate459inter4));
  nand2 gate930(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate931(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate932(.a(G21), .O(gate459inter7));
  inv1  gate933(.a(G1192), .O(gate459inter8));
  nand2 gate934(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate935(.a(s_55), .b(gate459inter3), .O(gate459inter10));
  nor2  gate936(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate937(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate938(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate855(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate856(.a(gate460inter0), .b(s_44), .O(gate460inter1));
  and2  gate857(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate858(.a(s_44), .O(gate460inter3));
  inv1  gate859(.a(s_45), .O(gate460inter4));
  nand2 gate860(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate861(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate862(.a(G1096), .O(gate460inter7));
  inv1  gate863(.a(G1192), .O(gate460inter8));
  nand2 gate864(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate865(.a(s_45), .b(gate460inter3), .O(gate460inter10));
  nor2  gate866(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate867(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate868(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2045(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2046(.a(gate461inter0), .b(s_214), .O(gate461inter1));
  and2  gate2047(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2048(.a(s_214), .O(gate461inter3));
  inv1  gate2049(.a(s_215), .O(gate461inter4));
  nand2 gate2050(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2051(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2052(.a(G22), .O(gate461inter7));
  inv1  gate2053(.a(G1195), .O(gate461inter8));
  nand2 gate2054(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2055(.a(s_215), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2056(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2057(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2058(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2493(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2494(.a(gate464inter0), .b(s_278), .O(gate464inter1));
  and2  gate2495(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2496(.a(s_278), .O(gate464inter3));
  inv1  gate2497(.a(s_279), .O(gate464inter4));
  nand2 gate2498(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2499(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2500(.a(G1102), .O(gate464inter7));
  inv1  gate2501(.a(G1198), .O(gate464inter8));
  nand2 gate2502(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2503(.a(s_279), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2504(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2505(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2506(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2255(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2256(.a(gate466inter0), .b(s_244), .O(gate466inter1));
  and2  gate2257(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2258(.a(s_244), .O(gate466inter3));
  inv1  gate2259(.a(s_245), .O(gate466inter4));
  nand2 gate2260(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2261(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2262(.a(G1105), .O(gate466inter7));
  inv1  gate2263(.a(G1201), .O(gate466inter8));
  nand2 gate2264(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2265(.a(s_245), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2266(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2267(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2268(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1247(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1248(.a(gate468inter0), .b(s_100), .O(gate468inter1));
  and2  gate1249(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1250(.a(s_100), .O(gate468inter3));
  inv1  gate1251(.a(s_101), .O(gate468inter4));
  nand2 gate1252(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1253(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1254(.a(G1108), .O(gate468inter7));
  inv1  gate1255(.a(G1204), .O(gate468inter8));
  nand2 gate1256(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1257(.a(s_101), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1258(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1259(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1260(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate897(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate898(.a(gate469inter0), .b(s_50), .O(gate469inter1));
  and2  gate899(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate900(.a(s_50), .O(gate469inter3));
  inv1  gate901(.a(s_51), .O(gate469inter4));
  nand2 gate902(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate903(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate904(.a(G26), .O(gate469inter7));
  inv1  gate905(.a(G1207), .O(gate469inter8));
  nand2 gate906(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate907(.a(s_51), .b(gate469inter3), .O(gate469inter10));
  nor2  gate908(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate909(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate910(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate1415(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1416(.a(gate470inter0), .b(s_124), .O(gate470inter1));
  and2  gate1417(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1418(.a(s_124), .O(gate470inter3));
  inv1  gate1419(.a(s_125), .O(gate470inter4));
  nand2 gate1420(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1421(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1422(.a(G1111), .O(gate470inter7));
  inv1  gate1423(.a(G1207), .O(gate470inter8));
  nand2 gate1424(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1425(.a(s_125), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1426(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1427(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1428(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1485(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1486(.a(gate471inter0), .b(s_134), .O(gate471inter1));
  and2  gate1487(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1488(.a(s_134), .O(gate471inter3));
  inv1  gate1489(.a(s_135), .O(gate471inter4));
  nand2 gate1490(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1491(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1492(.a(G27), .O(gate471inter7));
  inv1  gate1493(.a(G1210), .O(gate471inter8));
  nand2 gate1494(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1495(.a(s_135), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1496(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1497(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1498(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1555(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1556(.a(gate473inter0), .b(s_144), .O(gate473inter1));
  and2  gate1557(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1558(.a(s_144), .O(gate473inter3));
  inv1  gate1559(.a(s_145), .O(gate473inter4));
  nand2 gate1560(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1561(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1562(.a(G28), .O(gate473inter7));
  inv1  gate1563(.a(G1213), .O(gate473inter8));
  nand2 gate1564(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1565(.a(s_145), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1566(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1567(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1568(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate1751(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1752(.a(gate474inter0), .b(s_172), .O(gate474inter1));
  and2  gate1753(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1754(.a(s_172), .O(gate474inter3));
  inv1  gate1755(.a(s_173), .O(gate474inter4));
  nand2 gate1756(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1757(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1758(.a(G1117), .O(gate474inter7));
  inv1  gate1759(.a(G1213), .O(gate474inter8));
  nand2 gate1760(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1761(.a(s_173), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1762(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1763(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1764(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1807(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1808(.a(gate476inter0), .b(s_180), .O(gate476inter1));
  and2  gate1809(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1810(.a(s_180), .O(gate476inter3));
  inv1  gate1811(.a(s_181), .O(gate476inter4));
  nand2 gate1812(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1813(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1814(.a(G1120), .O(gate476inter7));
  inv1  gate1815(.a(G1216), .O(gate476inter8));
  nand2 gate1816(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1817(.a(s_181), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1818(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1819(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1820(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1093(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1094(.a(gate477inter0), .b(s_78), .O(gate477inter1));
  and2  gate1095(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1096(.a(s_78), .O(gate477inter3));
  inv1  gate1097(.a(s_79), .O(gate477inter4));
  nand2 gate1098(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1099(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1100(.a(G30), .O(gate477inter7));
  inv1  gate1101(.a(G1219), .O(gate477inter8));
  nand2 gate1102(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1103(.a(s_79), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1104(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1105(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1106(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1863(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1864(.a(gate482inter0), .b(s_188), .O(gate482inter1));
  and2  gate1865(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1866(.a(s_188), .O(gate482inter3));
  inv1  gate1867(.a(s_189), .O(gate482inter4));
  nand2 gate1868(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1869(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1870(.a(G1129), .O(gate482inter7));
  inv1  gate1871(.a(G1225), .O(gate482inter8));
  nand2 gate1872(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1873(.a(s_189), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1874(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1875(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1876(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1009(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1010(.a(gate486inter0), .b(s_66), .O(gate486inter1));
  and2  gate1011(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1012(.a(s_66), .O(gate486inter3));
  inv1  gate1013(.a(s_67), .O(gate486inter4));
  nand2 gate1014(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1015(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1016(.a(G1234), .O(gate486inter7));
  inv1  gate1017(.a(G1235), .O(gate486inter8));
  nand2 gate1018(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1019(.a(s_67), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1020(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1021(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1022(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1709(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1710(.a(gate488inter0), .b(s_166), .O(gate488inter1));
  and2  gate1711(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1712(.a(s_166), .O(gate488inter3));
  inv1  gate1713(.a(s_167), .O(gate488inter4));
  nand2 gate1714(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1715(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1716(.a(G1238), .O(gate488inter7));
  inv1  gate1717(.a(G1239), .O(gate488inter8));
  nand2 gate1718(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1719(.a(s_167), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1720(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1721(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1722(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2017(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2018(.a(gate490inter0), .b(s_210), .O(gate490inter1));
  and2  gate2019(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2020(.a(s_210), .O(gate490inter3));
  inv1  gate2021(.a(s_211), .O(gate490inter4));
  nand2 gate2022(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2023(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2024(.a(G1242), .O(gate490inter7));
  inv1  gate2025(.a(G1243), .O(gate490inter8));
  nand2 gate2026(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2027(.a(s_211), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2028(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2029(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2030(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1849(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1850(.a(gate492inter0), .b(s_186), .O(gate492inter1));
  and2  gate1851(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1852(.a(s_186), .O(gate492inter3));
  inv1  gate1853(.a(s_187), .O(gate492inter4));
  nand2 gate1854(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1855(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1856(.a(G1246), .O(gate492inter7));
  inv1  gate1857(.a(G1247), .O(gate492inter8));
  nand2 gate1858(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1859(.a(s_187), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1860(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1861(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1862(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1821(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1822(.a(gate493inter0), .b(s_182), .O(gate493inter1));
  and2  gate1823(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1824(.a(s_182), .O(gate493inter3));
  inv1  gate1825(.a(s_183), .O(gate493inter4));
  nand2 gate1826(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1827(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1828(.a(G1248), .O(gate493inter7));
  inv1  gate1829(.a(G1249), .O(gate493inter8));
  nand2 gate1830(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1831(.a(s_183), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1832(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1833(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1834(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate631(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate632(.a(gate494inter0), .b(s_12), .O(gate494inter1));
  and2  gate633(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate634(.a(s_12), .O(gate494inter3));
  inv1  gate635(.a(s_13), .O(gate494inter4));
  nand2 gate636(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate637(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate638(.a(G1250), .O(gate494inter7));
  inv1  gate639(.a(G1251), .O(gate494inter8));
  nand2 gate640(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate641(.a(s_13), .b(gate494inter3), .O(gate494inter10));
  nor2  gate642(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate643(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate644(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate883(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate884(.a(gate496inter0), .b(s_48), .O(gate496inter1));
  and2  gate885(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate886(.a(s_48), .O(gate496inter3));
  inv1  gate887(.a(s_49), .O(gate496inter4));
  nand2 gate888(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate889(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate890(.a(G1254), .O(gate496inter7));
  inv1  gate891(.a(G1255), .O(gate496inter8));
  nand2 gate892(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate893(.a(s_49), .b(gate496inter3), .O(gate496inter10));
  nor2  gate894(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate895(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate896(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1653(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1654(.a(gate497inter0), .b(s_158), .O(gate497inter1));
  and2  gate1655(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1656(.a(s_158), .O(gate497inter3));
  inv1  gate1657(.a(s_159), .O(gate497inter4));
  nand2 gate1658(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1659(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1660(.a(G1256), .O(gate497inter7));
  inv1  gate1661(.a(G1257), .O(gate497inter8));
  nand2 gate1662(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1663(.a(s_159), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1664(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1665(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1666(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2031(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2032(.a(gate502inter0), .b(s_212), .O(gate502inter1));
  and2  gate2033(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2034(.a(s_212), .O(gate502inter3));
  inv1  gate2035(.a(s_213), .O(gate502inter4));
  nand2 gate2036(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2037(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2038(.a(G1266), .O(gate502inter7));
  inv1  gate2039(.a(G1267), .O(gate502inter8));
  nand2 gate2040(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2041(.a(s_213), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2042(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2043(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2044(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2269(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2270(.a(gate514inter0), .b(s_246), .O(gate514inter1));
  and2  gate2271(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2272(.a(s_246), .O(gate514inter3));
  inv1  gate2273(.a(s_247), .O(gate514inter4));
  nand2 gate2274(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2275(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2276(.a(G1290), .O(gate514inter7));
  inv1  gate2277(.a(G1291), .O(gate514inter8));
  nand2 gate2278(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2279(.a(s_247), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2280(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2281(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2282(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule