module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381, s_382, s_383, s_384, s_385, s_386, s_387, s_388, s_389, s_390, s_391, s_392, s_393, s_394, s_395, s_396, s_397, s_398, s_399, s_400, s_401;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate995(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate996(.a(gate9inter0), .b(s_64), .O(gate9inter1));
  and2  gate997(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate998(.a(s_64), .O(gate9inter3));
  inv1  gate999(.a(s_65), .O(gate9inter4));
  nand2 gate1000(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1001(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1002(.a(G1), .O(gate9inter7));
  inv1  gate1003(.a(G2), .O(gate9inter8));
  nand2 gate1004(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1005(.a(s_65), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1006(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1007(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1008(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1373(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1374(.a(gate11inter0), .b(s_118), .O(gate11inter1));
  and2  gate1375(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1376(.a(s_118), .O(gate11inter3));
  inv1  gate1377(.a(s_119), .O(gate11inter4));
  nand2 gate1378(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1379(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1380(.a(G5), .O(gate11inter7));
  inv1  gate1381(.a(G6), .O(gate11inter8));
  nand2 gate1382(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1383(.a(s_119), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1384(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1385(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1386(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2185(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2186(.a(gate12inter0), .b(s_234), .O(gate12inter1));
  and2  gate2187(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2188(.a(s_234), .O(gate12inter3));
  inv1  gate2189(.a(s_235), .O(gate12inter4));
  nand2 gate2190(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2191(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2192(.a(G7), .O(gate12inter7));
  inv1  gate2193(.a(G8), .O(gate12inter8));
  nand2 gate2194(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2195(.a(s_235), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2196(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2197(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2198(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate897(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate898(.a(gate14inter0), .b(s_50), .O(gate14inter1));
  and2  gate899(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate900(.a(s_50), .O(gate14inter3));
  inv1  gate901(.a(s_51), .O(gate14inter4));
  nand2 gate902(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate903(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate904(.a(G11), .O(gate14inter7));
  inv1  gate905(.a(G12), .O(gate14inter8));
  nand2 gate906(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate907(.a(s_51), .b(gate14inter3), .O(gate14inter10));
  nor2  gate908(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate909(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate910(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1625(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1626(.a(gate16inter0), .b(s_154), .O(gate16inter1));
  and2  gate1627(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1628(.a(s_154), .O(gate16inter3));
  inv1  gate1629(.a(s_155), .O(gate16inter4));
  nand2 gate1630(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1631(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1632(.a(G15), .O(gate16inter7));
  inv1  gate1633(.a(G16), .O(gate16inter8));
  nand2 gate1634(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1635(.a(s_155), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1636(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1637(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1638(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2017(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2018(.a(gate17inter0), .b(s_210), .O(gate17inter1));
  and2  gate2019(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2020(.a(s_210), .O(gate17inter3));
  inv1  gate2021(.a(s_211), .O(gate17inter4));
  nand2 gate2022(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2023(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2024(.a(G17), .O(gate17inter7));
  inv1  gate2025(.a(G18), .O(gate17inter8));
  nand2 gate2026(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2027(.a(s_211), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2028(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2029(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2030(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1289(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1290(.a(gate18inter0), .b(s_106), .O(gate18inter1));
  and2  gate1291(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1292(.a(s_106), .O(gate18inter3));
  inv1  gate1293(.a(s_107), .O(gate18inter4));
  nand2 gate1294(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1295(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1296(.a(G19), .O(gate18inter7));
  inv1  gate1297(.a(G20), .O(gate18inter8));
  nand2 gate1298(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1299(.a(s_107), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1300(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1301(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1302(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2941(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2942(.a(gate19inter0), .b(s_342), .O(gate19inter1));
  and2  gate2943(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2944(.a(s_342), .O(gate19inter3));
  inv1  gate2945(.a(s_343), .O(gate19inter4));
  nand2 gate2946(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2947(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2948(.a(G21), .O(gate19inter7));
  inv1  gate2949(.a(G22), .O(gate19inter8));
  nand2 gate2950(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2951(.a(s_343), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2952(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2953(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2954(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate911(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate912(.a(gate20inter0), .b(s_52), .O(gate20inter1));
  and2  gate913(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate914(.a(s_52), .O(gate20inter3));
  inv1  gate915(.a(s_53), .O(gate20inter4));
  nand2 gate916(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate917(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate918(.a(G23), .O(gate20inter7));
  inv1  gate919(.a(G24), .O(gate20inter8));
  nand2 gate920(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate921(.a(s_53), .b(gate20inter3), .O(gate20inter10));
  nor2  gate922(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate923(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate924(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1275(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1276(.a(gate23inter0), .b(s_104), .O(gate23inter1));
  and2  gate1277(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1278(.a(s_104), .O(gate23inter3));
  inv1  gate1279(.a(s_105), .O(gate23inter4));
  nand2 gate1280(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1281(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1282(.a(G29), .O(gate23inter7));
  inv1  gate1283(.a(G30), .O(gate23inter8));
  nand2 gate1284(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1285(.a(s_105), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1286(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1287(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1288(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2661(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2662(.a(gate25inter0), .b(s_302), .O(gate25inter1));
  and2  gate2663(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2664(.a(s_302), .O(gate25inter3));
  inv1  gate2665(.a(s_303), .O(gate25inter4));
  nand2 gate2666(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2667(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2668(.a(G1), .O(gate25inter7));
  inv1  gate2669(.a(G5), .O(gate25inter8));
  nand2 gate2670(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2671(.a(s_303), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2672(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2673(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2674(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate3179(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate3180(.a(gate26inter0), .b(s_376), .O(gate26inter1));
  and2  gate3181(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate3182(.a(s_376), .O(gate26inter3));
  inv1  gate3183(.a(s_377), .O(gate26inter4));
  nand2 gate3184(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate3185(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate3186(.a(G9), .O(gate26inter7));
  inv1  gate3187(.a(G13), .O(gate26inter8));
  nand2 gate3188(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate3189(.a(s_377), .b(gate26inter3), .O(gate26inter10));
  nor2  gate3190(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate3191(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate3192(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate799(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate800(.a(gate29inter0), .b(s_36), .O(gate29inter1));
  and2  gate801(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate802(.a(s_36), .O(gate29inter3));
  inv1  gate803(.a(s_37), .O(gate29inter4));
  nand2 gate804(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate805(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate806(.a(G3), .O(gate29inter7));
  inv1  gate807(.a(G7), .O(gate29inter8));
  nand2 gate808(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate809(.a(s_37), .b(gate29inter3), .O(gate29inter10));
  nor2  gate810(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate811(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate812(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2339(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2340(.a(gate30inter0), .b(s_256), .O(gate30inter1));
  and2  gate2341(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2342(.a(s_256), .O(gate30inter3));
  inv1  gate2343(.a(s_257), .O(gate30inter4));
  nand2 gate2344(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2345(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2346(.a(G11), .O(gate30inter7));
  inv1  gate2347(.a(G15), .O(gate30inter8));
  nand2 gate2348(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2349(.a(s_257), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2350(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2351(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2352(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate827(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate828(.a(gate33inter0), .b(s_40), .O(gate33inter1));
  and2  gate829(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate830(.a(s_40), .O(gate33inter3));
  inv1  gate831(.a(s_41), .O(gate33inter4));
  nand2 gate832(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate833(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate834(.a(G17), .O(gate33inter7));
  inv1  gate835(.a(G21), .O(gate33inter8));
  nand2 gate836(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate837(.a(s_41), .b(gate33inter3), .O(gate33inter10));
  nor2  gate838(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate839(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate840(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1331(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1332(.a(gate34inter0), .b(s_112), .O(gate34inter1));
  and2  gate1333(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1334(.a(s_112), .O(gate34inter3));
  inv1  gate1335(.a(s_113), .O(gate34inter4));
  nand2 gate1336(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1337(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1338(.a(G25), .O(gate34inter7));
  inv1  gate1339(.a(G29), .O(gate34inter8));
  nand2 gate1340(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1341(.a(s_113), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1342(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1343(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1344(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1765(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1766(.a(gate35inter0), .b(s_174), .O(gate35inter1));
  and2  gate1767(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1768(.a(s_174), .O(gate35inter3));
  inv1  gate1769(.a(s_175), .O(gate35inter4));
  nand2 gate1770(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1771(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1772(.a(G18), .O(gate35inter7));
  inv1  gate1773(.a(G22), .O(gate35inter8));
  nand2 gate1774(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1775(.a(s_175), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1776(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1777(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1778(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2367(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2368(.a(gate36inter0), .b(s_260), .O(gate36inter1));
  and2  gate2369(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2370(.a(s_260), .O(gate36inter3));
  inv1  gate2371(.a(s_261), .O(gate36inter4));
  nand2 gate2372(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2373(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2374(.a(G26), .O(gate36inter7));
  inv1  gate2375(.a(G30), .O(gate36inter8));
  nand2 gate2376(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2377(.a(s_261), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2378(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2379(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2380(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1135(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1136(.a(gate38inter0), .b(s_84), .O(gate38inter1));
  and2  gate1137(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1138(.a(s_84), .O(gate38inter3));
  inv1  gate1139(.a(s_85), .O(gate38inter4));
  nand2 gate1140(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1141(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1142(.a(G27), .O(gate38inter7));
  inv1  gate1143(.a(G31), .O(gate38inter8));
  nand2 gate1144(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1145(.a(s_85), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1146(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1147(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1148(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1443(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1444(.a(gate40inter0), .b(s_128), .O(gate40inter1));
  and2  gate1445(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1446(.a(s_128), .O(gate40inter3));
  inv1  gate1447(.a(s_129), .O(gate40inter4));
  nand2 gate1448(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1449(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1450(.a(G28), .O(gate40inter7));
  inv1  gate1451(.a(G32), .O(gate40inter8));
  nand2 gate1452(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1453(.a(s_129), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1454(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1455(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1456(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1709(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1710(.a(gate41inter0), .b(s_166), .O(gate41inter1));
  and2  gate1711(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1712(.a(s_166), .O(gate41inter3));
  inv1  gate1713(.a(s_167), .O(gate41inter4));
  nand2 gate1714(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1715(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1716(.a(G1), .O(gate41inter7));
  inv1  gate1717(.a(G266), .O(gate41inter8));
  nand2 gate1718(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1719(.a(s_167), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1720(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1721(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1722(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate981(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate982(.a(gate42inter0), .b(s_62), .O(gate42inter1));
  and2  gate983(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate984(.a(s_62), .O(gate42inter3));
  inv1  gate985(.a(s_63), .O(gate42inter4));
  nand2 gate986(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate987(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate988(.a(G2), .O(gate42inter7));
  inv1  gate989(.a(G266), .O(gate42inter8));
  nand2 gate990(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate991(.a(s_63), .b(gate42inter3), .O(gate42inter10));
  nor2  gate992(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate993(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate994(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1051(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1052(.a(gate43inter0), .b(s_72), .O(gate43inter1));
  and2  gate1053(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1054(.a(s_72), .O(gate43inter3));
  inv1  gate1055(.a(s_73), .O(gate43inter4));
  nand2 gate1056(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1057(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1058(.a(G3), .O(gate43inter7));
  inv1  gate1059(.a(G269), .O(gate43inter8));
  nand2 gate1060(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1061(.a(s_73), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1062(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1063(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1064(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate3053(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate3054(.a(gate44inter0), .b(s_358), .O(gate44inter1));
  and2  gate3055(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate3056(.a(s_358), .O(gate44inter3));
  inv1  gate3057(.a(s_359), .O(gate44inter4));
  nand2 gate3058(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate3059(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate3060(.a(G4), .O(gate44inter7));
  inv1  gate3061(.a(G269), .O(gate44inter8));
  nand2 gate3062(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate3063(.a(s_359), .b(gate44inter3), .O(gate44inter10));
  nor2  gate3064(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate3065(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate3066(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2689(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2690(.a(gate45inter0), .b(s_306), .O(gate45inter1));
  and2  gate2691(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2692(.a(s_306), .O(gate45inter3));
  inv1  gate2693(.a(s_307), .O(gate45inter4));
  nand2 gate2694(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2695(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2696(.a(G5), .O(gate45inter7));
  inv1  gate2697(.a(G272), .O(gate45inter8));
  nand2 gate2698(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2699(.a(s_307), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2700(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2701(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2702(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1541(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1542(.a(gate46inter0), .b(s_142), .O(gate46inter1));
  and2  gate1543(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1544(.a(s_142), .O(gate46inter3));
  inv1  gate1545(.a(s_143), .O(gate46inter4));
  nand2 gate1546(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1547(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1548(.a(G6), .O(gate46inter7));
  inv1  gate1549(.a(G272), .O(gate46inter8));
  nand2 gate1550(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1551(.a(s_143), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1552(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1553(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1554(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate925(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate926(.a(gate47inter0), .b(s_54), .O(gate47inter1));
  and2  gate927(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate928(.a(s_54), .O(gate47inter3));
  inv1  gate929(.a(s_55), .O(gate47inter4));
  nand2 gate930(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate931(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate932(.a(G7), .O(gate47inter7));
  inv1  gate933(.a(G275), .O(gate47inter8));
  nand2 gate934(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate935(.a(s_55), .b(gate47inter3), .O(gate47inter10));
  nor2  gate936(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate937(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate938(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate953(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate954(.a(gate49inter0), .b(s_58), .O(gate49inter1));
  and2  gate955(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate956(.a(s_58), .O(gate49inter3));
  inv1  gate957(.a(s_59), .O(gate49inter4));
  nand2 gate958(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate959(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate960(.a(G9), .O(gate49inter7));
  inv1  gate961(.a(G278), .O(gate49inter8));
  nand2 gate962(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate963(.a(s_59), .b(gate49inter3), .O(gate49inter10));
  nor2  gate964(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate965(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate966(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1317(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1318(.a(gate50inter0), .b(s_110), .O(gate50inter1));
  and2  gate1319(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1320(.a(s_110), .O(gate50inter3));
  inv1  gate1321(.a(s_111), .O(gate50inter4));
  nand2 gate1322(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1323(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1324(.a(G10), .O(gate50inter7));
  inv1  gate1325(.a(G278), .O(gate50inter8));
  nand2 gate1326(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1327(.a(s_111), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1328(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1329(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1330(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate785(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate786(.a(gate52inter0), .b(s_34), .O(gate52inter1));
  and2  gate787(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate788(.a(s_34), .O(gate52inter3));
  inv1  gate789(.a(s_35), .O(gate52inter4));
  nand2 gate790(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate791(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate792(.a(G12), .O(gate52inter7));
  inv1  gate793(.a(G281), .O(gate52inter8));
  nand2 gate794(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate795(.a(s_35), .b(gate52inter3), .O(gate52inter10));
  nor2  gate796(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate797(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate798(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate575(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate576(.a(gate54inter0), .b(s_4), .O(gate54inter1));
  and2  gate577(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate578(.a(s_4), .O(gate54inter3));
  inv1  gate579(.a(s_5), .O(gate54inter4));
  nand2 gate580(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate581(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate582(.a(G14), .O(gate54inter7));
  inv1  gate583(.a(G284), .O(gate54inter8));
  nand2 gate584(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate585(.a(s_5), .b(gate54inter3), .O(gate54inter10));
  nor2  gate586(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate587(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate588(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate3263(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate3264(.a(gate62inter0), .b(s_388), .O(gate62inter1));
  and2  gate3265(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate3266(.a(s_388), .O(gate62inter3));
  inv1  gate3267(.a(s_389), .O(gate62inter4));
  nand2 gate3268(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate3269(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate3270(.a(G22), .O(gate62inter7));
  inv1  gate3271(.a(G296), .O(gate62inter8));
  nand2 gate3272(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate3273(.a(s_389), .b(gate62inter3), .O(gate62inter10));
  nor2  gate3274(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate3275(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate3276(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate2157(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2158(.a(gate65inter0), .b(s_230), .O(gate65inter1));
  and2  gate2159(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2160(.a(s_230), .O(gate65inter3));
  inv1  gate2161(.a(s_231), .O(gate65inter4));
  nand2 gate2162(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2163(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2164(.a(G25), .O(gate65inter7));
  inv1  gate2165(.a(G302), .O(gate65inter8));
  nand2 gate2166(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2167(.a(s_231), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2168(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2169(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2170(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1023(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1024(.a(gate66inter0), .b(s_68), .O(gate66inter1));
  and2  gate1025(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1026(.a(s_68), .O(gate66inter3));
  inv1  gate1027(.a(s_69), .O(gate66inter4));
  nand2 gate1028(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1029(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1030(.a(G26), .O(gate66inter7));
  inv1  gate1031(.a(G302), .O(gate66inter8));
  nand2 gate1032(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1033(.a(s_69), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1034(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1035(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1036(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate673(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate674(.a(gate67inter0), .b(s_18), .O(gate67inter1));
  and2  gate675(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate676(.a(s_18), .O(gate67inter3));
  inv1  gate677(.a(s_19), .O(gate67inter4));
  nand2 gate678(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate679(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate680(.a(G27), .O(gate67inter7));
  inv1  gate681(.a(G305), .O(gate67inter8));
  nand2 gate682(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate683(.a(s_19), .b(gate67inter3), .O(gate67inter10));
  nor2  gate684(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate685(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate686(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate2003(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2004(.a(gate68inter0), .b(s_208), .O(gate68inter1));
  and2  gate2005(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2006(.a(s_208), .O(gate68inter3));
  inv1  gate2007(.a(s_209), .O(gate68inter4));
  nand2 gate2008(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2009(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2010(.a(G28), .O(gate68inter7));
  inv1  gate2011(.a(G305), .O(gate68inter8));
  nand2 gate2012(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2013(.a(s_209), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2014(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2015(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2016(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate2507(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2508(.a(gate69inter0), .b(s_280), .O(gate69inter1));
  and2  gate2509(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2510(.a(s_280), .O(gate69inter3));
  inv1  gate2511(.a(s_281), .O(gate69inter4));
  nand2 gate2512(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2513(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2514(.a(G29), .O(gate69inter7));
  inv1  gate2515(.a(G308), .O(gate69inter8));
  nand2 gate2516(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2517(.a(s_281), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2518(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2519(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2520(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate3123(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate3124(.a(gate72inter0), .b(s_368), .O(gate72inter1));
  and2  gate3125(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate3126(.a(s_368), .O(gate72inter3));
  inv1  gate3127(.a(s_369), .O(gate72inter4));
  nand2 gate3128(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate3129(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate3130(.a(G32), .O(gate72inter7));
  inv1  gate3131(.a(G311), .O(gate72inter8));
  nand2 gate3132(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate3133(.a(s_369), .b(gate72inter3), .O(gate72inter10));
  nor2  gate3134(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate3135(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate3136(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1345(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1346(.a(gate74inter0), .b(s_114), .O(gate74inter1));
  and2  gate1347(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1348(.a(s_114), .O(gate74inter3));
  inv1  gate1349(.a(s_115), .O(gate74inter4));
  nand2 gate1350(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1351(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1352(.a(G5), .O(gate74inter7));
  inv1  gate1353(.a(G314), .O(gate74inter8));
  nand2 gate1354(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1355(.a(s_115), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1356(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1357(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1358(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate2605(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2606(.a(gate75inter0), .b(s_294), .O(gate75inter1));
  and2  gate2607(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2608(.a(s_294), .O(gate75inter3));
  inv1  gate2609(.a(s_295), .O(gate75inter4));
  nand2 gate2610(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2611(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2612(.a(G9), .O(gate75inter7));
  inv1  gate2613(.a(G317), .O(gate75inter8));
  nand2 gate2614(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2615(.a(s_295), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2616(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2617(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2618(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1583(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1584(.a(gate78inter0), .b(s_148), .O(gate78inter1));
  and2  gate1585(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1586(.a(s_148), .O(gate78inter3));
  inv1  gate1587(.a(s_149), .O(gate78inter4));
  nand2 gate1588(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1589(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1590(.a(G6), .O(gate78inter7));
  inv1  gate1591(.a(G320), .O(gate78inter8));
  nand2 gate1592(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1593(.a(s_149), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1594(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1595(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1596(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2423(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2424(.a(gate82inter0), .b(s_268), .O(gate82inter1));
  and2  gate2425(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2426(.a(s_268), .O(gate82inter3));
  inv1  gate2427(.a(s_269), .O(gate82inter4));
  nand2 gate2428(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2429(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2430(.a(G7), .O(gate82inter7));
  inv1  gate2431(.a(G326), .O(gate82inter8));
  nand2 gate2432(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2433(.a(s_269), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2434(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2435(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2436(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1919(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1920(.a(gate83inter0), .b(s_196), .O(gate83inter1));
  and2  gate1921(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1922(.a(s_196), .O(gate83inter3));
  inv1  gate1923(.a(s_197), .O(gate83inter4));
  nand2 gate1924(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1925(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1926(.a(G11), .O(gate83inter7));
  inv1  gate1927(.a(G329), .O(gate83inter8));
  nand2 gate1928(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1929(.a(s_197), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1930(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1931(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1932(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2465(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2466(.a(gate86inter0), .b(s_274), .O(gate86inter1));
  and2  gate2467(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2468(.a(s_274), .O(gate86inter3));
  inv1  gate2469(.a(s_275), .O(gate86inter4));
  nand2 gate2470(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2471(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2472(.a(G8), .O(gate86inter7));
  inv1  gate2473(.a(G332), .O(gate86inter8));
  nand2 gate2474(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2475(.a(s_275), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2476(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2477(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2478(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2843(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2844(.a(gate87inter0), .b(s_328), .O(gate87inter1));
  and2  gate2845(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2846(.a(s_328), .O(gate87inter3));
  inv1  gate2847(.a(s_329), .O(gate87inter4));
  nand2 gate2848(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2849(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2850(.a(G12), .O(gate87inter7));
  inv1  gate2851(.a(G335), .O(gate87inter8));
  nand2 gate2852(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2853(.a(s_329), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2854(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2855(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2856(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2045(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2046(.a(gate89inter0), .b(s_214), .O(gate89inter1));
  and2  gate2047(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2048(.a(s_214), .O(gate89inter3));
  inv1  gate2049(.a(s_215), .O(gate89inter4));
  nand2 gate2050(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2051(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2052(.a(G17), .O(gate89inter7));
  inv1  gate2053(.a(G338), .O(gate89inter8));
  nand2 gate2054(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2055(.a(s_215), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2056(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2057(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2058(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1891(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1892(.a(gate92inter0), .b(s_192), .O(gate92inter1));
  and2  gate1893(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1894(.a(s_192), .O(gate92inter3));
  inv1  gate1895(.a(s_193), .O(gate92inter4));
  nand2 gate1896(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1897(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1898(.a(G29), .O(gate92inter7));
  inv1  gate1899(.a(G341), .O(gate92inter8));
  nand2 gate1900(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1901(.a(s_193), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1902(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1903(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1904(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2437(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2438(.a(gate102inter0), .b(s_270), .O(gate102inter1));
  and2  gate2439(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2440(.a(s_270), .O(gate102inter3));
  inv1  gate2441(.a(s_271), .O(gate102inter4));
  nand2 gate2442(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2443(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2444(.a(G24), .O(gate102inter7));
  inv1  gate2445(.a(G356), .O(gate102inter8));
  nand2 gate2446(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2447(.a(s_271), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2448(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2449(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2450(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1457(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1458(.a(gate105inter0), .b(s_130), .O(gate105inter1));
  and2  gate1459(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1460(.a(s_130), .O(gate105inter3));
  inv1  gate1461(.a(s_131), .O(gate105inter4));
  nand2 gate1462(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1463(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1464(.a(G362), .O(gate105inter7));
  inv1  gate1465(.a(G363), .O(gate105inter8));
  nand2 gate1466(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1467(.a(s_131), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1468(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1469(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1470(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate869(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate870(.a(gate106inter0), .b(s_46), .O(gate106inter1));
  and2  gate871(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate872(.a(s_46), .O(gate106inter3));
  inv1  gate873(.a(s_47), .O(gate106inter4));
  nand2 gate874(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate875(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate876(.a(G364), .O(gate106inter7));
  inv1  gate877(.a(G365), .O(gate106inter8));
  nand2 gate878(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate879(.a(s_47), .b(gate106inter3), .O(gate106inter10));
  nor2  gate880(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate881(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate882(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1121(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1122(.a(gate109inter0), .b(s_82), .O(gate109inter1));
  and2  gate1123(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1124(.a(s_82), .O(gate109inter3));
  inv1  gate1125(.a(s_83), .O(gate109inter4));
  nand2 gate1126(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1127(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1128(.a(G370), .O(gate109inter7));
  inv1  gate1129(.a(G371), .O(gate109inter8));
  nand2 gate1130(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1131(.a(s_83), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1132(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1133(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1134(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1401(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1402(.a(gate110inter0), .b(s_122), .O(gate110inter1));
  and2  gate1403(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1404(.a(s_122), .O(gate110inter3));
  inv1  gate1405(.a(s_123), .O(gate110inter4));
  nand2 gate1406(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1407(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1408(.a(G372), .O(gate110inter7));
  inv1  gate1409(.a(G373), .O(gate110inter8));
  nand2 gate1410(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1411(.a(s_123), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1412(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1413(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1414(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2969(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2970(.a(gate111inter0), .b(s_346), .O(gate111inter1));
  and2  gate2971(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2972(.a(s_346), .O(gate111inter3));
  inv1  gate2973(.a(s_347), .O(gate111inter4));
  nand2 gate2974(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2975(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2976(.a(G374), .O(gate111inter7));
  inv1  gate2977(.a(G375), .O(gate111inter8));
  nand2 gate2978(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2979(.a(s_347), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2980(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2981(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2982(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1499(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1500(.a(gate112inter0), .b(s_136), .O(gate112inter1));
  and2  gate1501(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1502(.a(s_136), .O(gate112inter3));
  inv1  gate1503(.a(s_137), .O(gate112inter4));
  nand2 gate1504(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1505(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1506(.a(G376), .O(gate112inter7));
  inv1  gate1507(.a(G377), .O(gate112inter8));
  nand2 gate1508(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1509(.a(s_137), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1510(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1511(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1512(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate2759(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2760(.a(gate113inter0), .b(s_316), .O(gate113inter1));
  and2  gate2761(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2762(.a(s_316), .O(gate113inter3));
  inv1  gate2763(.a(s_317), .O(gate113inter4));
  nand2 gate2764(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2765(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2766(.a(G378), .O(gate113inter7));
  inv1  gate2767(.a(G379), .O(gate113inter8));
  nand2 gate2768(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2769(.a(s_317), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2770(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2771(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2772(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1681(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1682(.a(gate115inter0), .b(s_162), .O(gate115inter1));
  and2  gate1683(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1684(.a(s_162), .O(gate115inter3));
  inv1  gate1685(.a(s_163), .O(gate115inter4));
  nand2 gate1686(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1687(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1688(.a(G382), .O(gate115inter7));
  inv1  gate1689(.a(G383), .O(gate115inter8));
  nand2 gate1690(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1691(.a(s_163), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1692(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1693(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1694(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2815(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2816(.a(gate118inter0), .b(s_324), .O(gate118inter1));
  and2  gate2817(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2818(.a(s_324), .O(gate118inter3));
  inv1  gate2819(.a(s_325), .O(gate118inter4));
  nand2 gate2820(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2821(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2822(.a(G388), .O(gate118inter7));
  inv1  gate2823(.a(G389), .O(gate118inter8));
  nand2 gate2824(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2825(.a(s_325), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2826(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2827(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2828(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2535(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2536(.a(gate122inter0), .b(s_284), .O(gate122inter1));
  and2  gate2537(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2538(.a(s_284), .O(gate122inter3));
  inv1  gate2539(.a(s_285), .O(gate122inter4));
  nand2 gate2540(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2541(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2542(.a(G396), .O(gate122inter7));
  inv1  gate2543(.a(G397), .O(gate122inter8));
  nand2 gate2544(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2545(.a(s_285), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2546(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2547(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2548(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1779(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1780(.a(gate125inter0), .b(s_176), .O(gate125inter1));
  and2  gate1781(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1782(.a(s_176), .O(gate125inter3));
  inv1  gate1783(.a(s_177), .O(gate125inter4));
  nand2 gate1784(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1785(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1786(.a(G402), .O(gate125inter7));
  inv1  gate1787(.a(G403), .O(gate125inter8));
  nand2 gate1788(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1789(.a(s_177), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1790(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1791(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1792(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate631(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate632(.a(gate130inter0), .b(s_12), .O(gate130inter1));
  and2  gate633(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate634(.a(s_12), .O(gate130inter3));
  inv1  gate635(.a(s_13), .O(gate130inter4));
  nand2 gate636(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate637(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate638(.a(G412), .O(gate130inter7));
  inv1  gate639(.a(G413), .O(gate130inter8));
  nand2 gate640(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate641(.a(s_13), .b(gate130inter3), .O(gate130inter10));
  nor2  gate642(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate643(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate644(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1905(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1906(.a(gate132inter0), .b(s_194), .O(gate132inter1));
  and2  gate1907(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1908(.a(s_194), .O(gate132inter3));
  inv1  gate1909(.a(s_195), .O(gate132inter4));
  nand2 gate1910(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1911(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1912(.a(G416), .O(gate132inter7));
  inv1  gate1913(.a(G417), .O(gate132inter8));
  nand2 gate1914(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1915(.a(s_195), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1916(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1917(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1918(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2675(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2676(.a(gate136inter0), .b(s_304), .O(gate136inter1));
  and2  gate2677(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2678(.a(s_304), .O(gate136inter3));
  inv1  gate2679(.a(s_305), .O(gate136inter4));
  nand2 gate2680(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2681(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2682(.a(G424), .O(gate136inter7));
  inv1  gate2683(.a(G425), .O(gate136inter8));
  nand2 gate2684(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2685(.a(s_305), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2686(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2687(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2688(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2227(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2228(.a(gate138inter0), .b(s_240), .O(gate138inter1));
  and2  gate2229(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2230(.a(s_240), .O(gate138inter3));
  inv1  gate2231(.a(s_241), .O(gate138inter4));
  nand2 gate2232(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2233(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2234(.a(G432), .O(gate138inter7));
  inv1  gate2235(.a(G435), .O(gate138inter8));
  nand2 gate2236(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2237(.a(s_241), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2238(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2239(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2240(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2171(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2172(.a(gate139inter0), .b(s_232), .O(gate139inter1));
  and2  gate2173(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2174(.a(s_232), .O(gate139inter3));
  inv1  gate2175(.a(s_233), .O(gate139inter4));
  nand2 gate2176(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2177(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2178(.a(G438), .O(gate139inter7));
  inv1  gate2179(.a(G441), .O(gate139inter8));
  nand2 gate2180(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2181(.a(s_233), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2182(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2183(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2184(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2787(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2788(.a(gate140inter0), .b(s_320), .O(gate140inter1));
  and2  gate2789(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2790(.a(s_320), .O(gate140inter3));
  inv1  gate2791(.a(s_321), .O(gate140inter4));
  nand2 gate2792(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2793(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2794(.a(G444), .O(gate140inter7));
  inv1  gate2795(.a(G447), .O(gate140inter8));
  nand2 gate2796(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2797(.a(s_321), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2798(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2799(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2800(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate2871(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate2872(.a(gate141inter0), .b(s_332), .O(gate141inter1));
  and2  gate2873(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate2874(.a(s_332), .O(gate141inter3));
  inv1  gate2875(.a(s_333), .O(gate141inter4));
  nand2 gate2876(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate2877(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate2878(.a(G450), .O(gate141inter7));
  inv1  gate2879(.a(G453), .O(gate141inter8));
  nand2 gate2880(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate2881(.a(s_333), .b(gate141inter3), .O(gate141inter10));
  nor2  gate2882(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate2883(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate2884(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate2451(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2452(.a(gate142inter0), .b(s_272), .O(gate142inter1));
  and2  gate2453(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2454(.a(s_272), .O(gate142inter3));
  inv1  gate2455(.a(s_273), .O(gate142inter4));
  nand2 gate2456(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2457(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2458(.a(G456), .O(gate142inter7));
  inv1  gate2459(.a(G459), .O(gate142inter8));
  nand2 gate2460(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2461(.a(s_273), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2462(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2463(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2464(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate729(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate730(.a(gate146inter0), .b(s_26), .O(gate146inter1));
  and2  gate731(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate732(.a(s_26), .O(gate146inter3));
  inv1  gate733(.a(s_27), .O(gate146inter4));
  nand2 gate734(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate735(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate736(.a(G480), .O(gate146inter7));
  inv1  gate737(.a(G483), .O(gate146inter8));
  nand2 gate738(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate739(.a(s_27), .b(gate146inter3), .O(gate146inter10));
  nor2  gate740(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate741(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate742(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2857(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2858(.a(gate149inter0), .b(s_330), .O(gate149inter1));
  and2  gate2859(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2860(.a(s_330), .O(gate149inter3));
  inv1  gate2861(.a(s_331), .O(gate149inter4));
  nand2 gate2862(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2863(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2864(.a(G498), .O(gate149inter7));
  inv1  gate2865(.a(G501), .O(gate149inter8));
  nand2 gate2866(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2867(.a(s_331), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2868(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2869(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2870(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate771(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate772(.a(gate150inter0), .b(s_32), .O(gate150inter1));
  and2  gate773(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate774(.a(s_32), .O(gate150inter3));
  inv1  gate775(.a(s_33), .O(gate150inter4));
  nand2 gate776(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate777(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate778(.a(G504), .O(gate150inter7));
  inv1  gate779(.a(G507), .O(gate150inter8));
  nand2 gate780(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate781(.a(s_33), .b(gate150inter3), .O(gate150inter10));
  nor2  gate782(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate783(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate784(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1093(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1094(.a(gate152inter0), .b(s_78), .O(gate152inter1));
  and2  gate1095(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1096(.a(s_78), .O(gate152inter3));
  inv1  gate1097(.a(s_79), .O(gate152inter4));
  nand2 gate1098(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1099(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1100(.a(G516), .O(gate152inter7));
  inv1  gate1101(.a(G519), .O(gate152inter8));
  nand2 gate1102(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1103(.a(s_79), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1104(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1105(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1106(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate2619(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2620(.a(gate153inter0), .b(s_296), .O(gate153inter1));
  and2  gate2621(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2622(.a(s_296), .O(gate153inter3));
  inv1  gate2623(.a(s_297), .O(gate153inter4));
  nand2 gate2624(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2625(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2626(.a(G426), .O(gate153inter7));
  inv1  gate2627(.a(G522), .O(gate153inter8));
  nand2 gate2628(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2629(.a(s_297), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2630(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2631(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2632(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1485(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1486(.a(gate155inter0), .b(s_134), .O(gate155inter1));
  and2  gate1487(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1488(.a(s_134), .O(gate155inter3));
  inv1  gate1489(.a(s_135), .O(gate155inter4));
  nand2 gate1490(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1491(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1492(.a(G432), .O(gate155inter7));
  inv1  gate1493(.a(G525), .O(gate155inter8));
  nand2 gate1494(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1495(.a(s_135), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1496(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1497(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1498(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2073(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2074(.a(gate160inter0), .b(s_218), .O(gate160inter1));
  and2  gate2075(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2076(.a(s_218), .O(gate160inter3));
  inv1  gate2077(.a(s_219), .O(gate160inter4));
  nand2 gate2078(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2079(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2080(.a(G447), .O(gate160inter7));
  inv1  gate2081(.a(G531), .O(gate160inter8));
  nand2 gate2082(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2083(.a(s_219), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2084(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2085(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2086(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2325(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2326(.a(gate164inter0), .b(s_254), .O(gate164inter1));
  and2  gate2327(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2328(.a(s_254), .O(gate164inter3));
  inv1  gate2329(.a(s_255), .O(gate164inter4));
  nand2 gate2330(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2331(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2332(.a(G459), .O(gate164inter7));
  inv1  gate2333(.a(G537), .O(gate164inter8));
  nand2 gate2334(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2335(.a(s_255), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2336(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2337(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2338(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1219(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1220(.a(gate168inter0), .b(s_96), .O(gate168inter1));
  and2  gate1221(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1222(.a(s_96), .O(gate168inter3));
  inv1  gate1223(.a(s_97), .O(gate168inter4));
  nand2 gate1224(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1225(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1226(.a(G471), .O(gate168inter7));
  inv1  gate1227(.a(G543), .O(gate168inter8));
  nand2 gate1228(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1229(.a(s_97), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1230(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1231(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1232(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2563(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2564(.a(gate170inter0), .b(s_288), .O(gate170inter1));
  and2  gate2565(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2566(.a(s_288), .O(gate170inter3));
  inv1  gate2567(.a(s_289), .O(gate170inter4));
  nand2 gate2568(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2569(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2570(.a(G477), .O(gate170inter7));
  inv1  gate2571(.a(G546), .O(gate170inter8));
  nand2 gate2572(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2573(.a(s_289), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2574(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2575(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2576(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate589(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate590(.a(gate171inter0), .b(s_6), .O(gate171inter1));
  and2  gate591(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate592(.a(s_6), .O(gate171inter3));
  inv1  gate593(.a(s_7), .O(gate171inter4));
  nand2 gate594(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate595(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate596(.a(G480), .O(gate171inter7));
  inv1  gate597(.a(G549), .O(gate171inter8));
  nand2 gate598(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate599(.a(s_7), .b(gate171inter3), .O(gate171inter10));
  nor2  gate600(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate601(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate602(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate3221(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate3222(.a(gate172inter0), .b(s_382), .O(gate172inter1));
  and2  gate3223(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate3224(.a(s_382), .O(gate172inter3));
  inv1  gate3225(.a(s_383), .O(gate172inter4));
  nand2 gate3226(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate3227(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate3228(.a(G483), .O(gate172inter7));
  inv1  gate3229(.a(G549), .O(gate172inter8));
  nand2 gate3230(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate3231(.a(s_383), .b(gate172inter3), .O(gate172inter10));
  nor2  gate3232(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate3233(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate3234(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2521(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2522(.a(gate174inter0), .b(s_282), .O(gate174inter1));
  and2  gate2523(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2524(.a(s_282), .O(gate174inter3));
  inv1  gate2525(.a(s_283), .O(gate174inter4));
  nand2 gate2526(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2527(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2528(.a(G489), .O(gate174inter7));
  inv1  gate2529(.a(G552), .O(gate174inter8));
  nand2 gate2530(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2531(.a(s_283), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2532(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2533(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2534(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate3249(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate3250(.a(gate176inter0), .b(s_386), .O(gate176inter1));
  and2  gate3251(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate3252(.a(s_386), .O(gate176inter3));
  inv1  gate3253(.a(s_387), .O(gate176inter4));
  nand2 gate3254(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate3255(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate3256(.a(G495), .O(gate176inter7));
  inv1  gate3257(.a(G555), .O(gate176inter8));
  nand2 gate3258(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate3259(.a(s_387), .b(gate176inter3), .O(gate176inter10));
  nor2  gate3260(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate3261(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate3262(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate1415(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1416(.a(gate177inter0), .b(s_124), .O(gate177inter1));
  and2  gate1417(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1418(.a(s_124), .O(gate177inter3));
  inv1  gate1419(.a(s_125), .O(gate177inter4));
  nand2 gate1420(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1421(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1422(.a(G498), .O(gate177inter7));
  inv1  gate1423(.a(G558), .O(gate177inter8));
  nand2 gate1424(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1425(.a(s_125), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1426(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1427(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1428(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate757(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate758(.a(gate179inter0), .b(s_30), .O(gate179inter1));
  and2  gate759(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate760(.a(s_30), .O(gate179inter3));
  inv1  gate761(.a(s_31), .O(gate179inter4));
  nand2 gate762(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate763(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate764(.a(G504), .O(gate179inter7));
  inv1  gate765(.a(G561), .O(gate179inter8));
  nand2 gate766(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate767(.a(s_31), .b(gate179inter3), .O(gate179inter10));
  nor2  gate768(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate769(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate770(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1653(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1654(.a(gate180inter0), .b(s_158), .O(gate180inter1));
  and2  gate1655(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1656(.a(s_158), .O(gate180inter3));
  inv1  gate1657(.a(s_159), .O(gate180inter4));
  nand2 gate1658(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1659(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1660(.a(G507), .O(gate180inter7));
  inv1  gate1661(.a(G561), .O(gate180inter8));
  nand2 gate1662(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1663(.a(s_159), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1664(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1665(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1666(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate687(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate688(.a(gate181inter0), .b(s_20), .O(gate181inter1));
  and2  gate689(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate690(.a(s_20), .O(gate181inter3));
  inv1  gate691(.a(s_21), .O(gate181inter4));
  nand2 gate692(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate693(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate694(.a(G510), .O(gate181inter7));
  inv1  gate695(.a(G564), .O(gate181inter8));
  nand2 gate696(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate697(.a(s_21), .b(gate181inter3), .O(gate181inter10));
  nor2  gate698(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate699(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate700(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2143(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2144(.a(gate182inter0), .b(s_228), .O(gate182inter1));
  and2  gate2145(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2146(.a(s_228), .O(gate182inter3));
  inv1  gate2147(.a(s_229), .O(gate182inter4));
  nand2 gate2148(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2149(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2150(.a(G513), .O(gate182inter7));
  inv1  gate2151(.a(G564), .O(gate182inter8));
  nand2 gate2152(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2153(.a(s_229), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2154(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2155(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2156(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1261(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1262(.a(gate185inter0), .b(s_102), .O(gate185inter1));
  and2  gate1263(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1264(.a(s_102), .O(gate185inter3));
  inv1  gate1265(.a(s_103), .O(gate185inter4));
  nand2 gate1266(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1267(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1268(.a(G570), .O(gate185inter7));
  inv1  gate1269(.a(G571), .O(gate185inter8));
  nand2 gate1270(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1271(.a(s_103), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1272(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1273(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1274(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1359(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1360(.a(gate191inter0), .b(s_116), .O(gate191inter1));
  and2  gate1361(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1362(.a(s_116), .O(gate191inter3));
  inv1  gate1363(.a(s_117), .O(gate191inter4));
  nand2 gate1364(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1365(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1366(.a(G582), .O(gate191inter7));
  inv1  gate1367(.a(G583), .O(gate191inter8));
  nand2 gate1368(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1369(.a(s_117), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1370(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1371(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1372(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2395(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2396(.a(gate194inter0), .b(s_264), .O(gate194inter1));
  and2  gate2397(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2398(.a(s_264), .O(gate194inter3));
  inv1  gate2399(.a(s_265), .O(gate194inter4));
  nand2 gate2400(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2401(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2402(.a(G588), .O(gate194inter7));
  inv1  gate2403(.a(G589), .O(gate194inter8));
  nand2 gate2404(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2405(.a(s_265), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2406(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2407(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2408(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate3319(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate3320(.a(gate197inter0), .b(s_396), .O(gate197inter1));
  and2  gate3321(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate3322(.a(s_396), .O(gate197inter3));
  inv1  gate3323(.a(s_397), .O(gate197inter4));
  nand2 gate3324(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate3325(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate3326(.a(G594), .O(gate197inter7));
  inv1  gate3327(.a(G595), .O(gate197inter8));
  nand2 gate3328(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate3329(.a(s_397), .b(gate197inter3), .O(gate197inter10));
  nor2  gate3330(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate3331(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate3332(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1107(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1108(.a(gate201inter0), .b(s_80), .O(gate201inter1));
  and2  gate1109(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1110(.a(s_80), .O(gate201inter3));
  inv1  gate1111(.a(s_81), .O(gate201inter4));
  nand2 gate1112(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1113(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1114(.a(G602), .O(gate201inter7));
  inv1  gate1115(.a(G607), .O(gate201inter8));
  nand2 gate1116(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1117(.a(s_81), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1118(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1119(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1120(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1079(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1080(.a(gate202inter0), .b(s_76), .O(gate202inter1));
  and2  gate1081(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1082(.a(s_76), .O(gate202inter3));
  inv1  gate1083(.a(s_77), .O(gate202inter4));
  nand2 gate1084(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1085(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1086(.a(G612), .O(gate202inter7));
  inv1  gate1087(.a(G617), .O(gate202inter8));
  nand2 gate1088(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1089(.a(s_77), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1090(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1091(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1092(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate701(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate702(.a(gate203inter0), .b(s_22), .O(gate203inter1));
  and2  gate703(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate704(.a(s_22), .O(gate203inter3));
  inv1  gate705(.a(s_23), .O(gate203inter4));
  nand2 gate706(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate707(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate708(.a(G602), .O(gate203inter7));
  inv1  gate709(.a(G612), .O(gate203inter8));
  nand2 gate710(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate711(.a(s_23), .b(gate203inter3), .O(gate203inter10));
  nor2  gate712(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate713(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate714(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate2241(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2242(.a(gate204inter0), .b(s_242), .O(gate204inter1));
  and2  gate2243(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2244(.a(s_242), .O(gate204inter3));
  inv1  gate2245(.a(s_243), .O(gate204inter4));
  nand2 gate2246(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2247(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2248(.a(G607), .O(gate204inter7));
  inv1  gate2249(.a(G617), .O(gate204inter8));
  nand2 gate2250(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2251(.a(s_243), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2252(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2253(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2254(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate603(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate604(.a(gate207inter0), .b(s_8), .O(gate207inter1));
  and2  gate605(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate606(.a(s_8), .O(gate207inter3));
  inv1  gate607(.a(s_9), .O(gate207inter4));
  nand2 gate608(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate609(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate610(.a(G622), .O(gate207inter7));
  inv1  gate611(.a(G632), .O(gate207inter8));
  nand2 gate612(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate613(.a(s_9), .b(gate207inter3), .O(gate207inter10));
  nor2  gate614(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate615(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate616(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1205(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1206(.a(gate210inter0), .b(s_94), .O(gate210inter1));
  and2  gate1207(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1208(.a(s_94), .O(gate210inter3));
  inv1  gate1209(.a(s_95), .O(gate210inter4));
  nand2 gate1210(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1211(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1212(.a(G607), .O(gate210inter7));
  inv1  gate1213(.a(G666), .O(gate210inter8));
  nand2 gate1214(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1215(.a(s_95), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1216(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1217(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1218(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1177(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1178(.a(gate211inter0), .b(s_90), .O(gate211inter1));
  and2  gate1179(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1180(.a(s_90), .O(gate211inter3));
  inv1  gate1181(.a(s_91), .O(gate211inter4));
  nand2 gate1182(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1183(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1184(.a(G612), .O(gate211inter7));
  inv1  gate1185(.a(G669), .O(gate211inter8));
  nand2 gate1186(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1187(.a(s_91), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1188(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1189(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1190(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate743(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate744(.a(gate212inter0), .b(s_28), .O(gate212inter1));
  and2  gate745(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate746(.a(s_28), .O(gate212inter3));
  inv1  gate747(.a(s_29), .O(gate212inter4));
  nand2 gate748(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate749(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate750(.a(G617), .O(gate212inter7));
  inv1  gate751(.a(G669), .O(gate212inter8));
  nand2 gate752(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate753(.a(s_29), .b(gate212inter3), .O(gate212inter10));
  nor2  gate754(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate755(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate756(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate813(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate814(.a(gate213inter0), .b(s_38), .O(gate213inter1));
  and2  gate815(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate816(.a(s_38), .O(gate213inter3));
  inv1  gate817(.a(s_39), .O(gate213inter4));
  nand2 gate818(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate819(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate820(.a(G602), .O(gate213inter7));
  inv1  gate821(.a(G672), .O(gate213inter8));
  nand2 gate822(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate823(.a(s_39), .b(gate213inter3), .O(gate213inter10));
  nor2  gate824(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate825(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate826(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2647(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2648(.a(gate214inter0), .b(s_300), .O(gate214inter1));
  and2  gate2649(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2650(.a(s_300), .O(gate214inter3));
  inv1  gate2651(.a(s_301), .O(gate214inter4));
  nand2 gate2652(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2653(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2654(.a(G612), .O(gate214inter7));
  inv1  gate2655(.a(G672), .O(gate214inter8));
  nand2 gate2656(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2657(.a(s_301), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2658(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2659(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2660(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2115(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2116(.a(gate216inter0), .b(s_224), .O(gate216inter1));
  and2  gate2117(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2118(.a(s_224), .O(gate216inter3));
  inv1  gate2119(.a(s_225), .O(gate216inter4));
  nand2 gate2120(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2121(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2122(.a(G617), .O(gate216inter7));
  inv1  gate2123(.a(G675), .O(gate216inter8));
  nand2 gate2124(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2125(.a(s_225), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2126(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2127(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2128(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2983(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2984(.a(gate219inter0), .b(s_348), .O(gate219inter1));
  and2  gate2985(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2986(.a(s_348), .O(gate219inter3));
  inv1  gate2987(.a(s_349), .O(gate219inter4));
  nand2 gate2988(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2989(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2990(.a(G632), .O(gate219inter7));
  inv1  gate2991(.a(G681), .O(gate219inter8));
  nand2 gate2992(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2993(.a(s_349), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2994(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2995(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2996(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2927(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2928(.a(gate220inter0), .b(s_340), .O(gate220inter1));
  and2  gate2929(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2930(.a(s_340), .O(gate220inter3));
  inv1  gate2931(.a(s_341), .O(gate220inter4));
  nand2 gate2932(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2933(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2934(.a(G637), .O(gate220inter7));
  inv1  gate2935(.a(G681), .O(gate220inter8));
  nand2 gate2936(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2937(.a(s_341), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2938(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2939(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2940(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1667(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1668(.a(gate224inter0), .b(s_160), .O(gate224inter1));
  and2  gate1669(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1670(.a(s_160), .O(gate224inter3));
  inv1  gate1671(.a(s_161), .O(gate224inter4));
  nand2 gate1672(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1673(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1674(.a(G637), .O(gate224inter7));
  inv1  gate1675(.a(G687), .O(gate224inter8));
  nand2 gate1676(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1677(.a(s_161), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1678(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1679(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1680(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2997(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2998(.a(gate227inter0), .b(s_350), .O(gate227inter1));
  and2  gate2999(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate3000(.a(s_350), .O(gate227inter3));
  inv1  gate3001(.a(s_351), .O(gate227inter4));
  nand2 gate3002(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate3003(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate3004(.a(G694), .O(gate227inter7));
  inv1  gate3005(.a(G695), .O(gate227inter8));
  nand2 gate3006(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate3007(.a(s_351), .b(gate227inter3), .O(gate227inter10));
  nor2  gate3008(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate3009(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate3010(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1065(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1066(.a(gate233inter0), .b(s_74), .O(gate233inter1));
  and2  gate1067(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1068(.a(s_74), .O(gate233inter3));
  inv1  gate1069(.a(s_75), .O(gate233inter4));
  nand2 gate1070(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1071(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1072(.a(G242), .O(gate233inter7));
  inv1  gate1073(.a(G718), .O(gate233inter8));
  nand2 gate1074(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1075(.a(s_75), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1076(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1077(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1078(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1877(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1878(.a(gate234inter0), .b(s_190), .O(gate234inter1));
  and2  gate1879(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1880(.a(s_190), .O(gate234inter3));
  inv1  gate1881(.a(s_191), .O(gate234inter4));
  nand2 gate1882(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1883(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1884(.a(G245), .O(gate234inter7));
  inv1  gate1885(.a(G721), .O(gate234inter8));
  nand2 gate1886(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1887(.a(s_191), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1888(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1889(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1890(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2479(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2480(.a(gate236inter0), .b(s_276), .O(gate236inter1));
  and2  gate2481(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2482(.a(s_276), .O(gate236inter3));
  inv1  gate2483(.a(s_277), .O(gate236inter4));
  nand2 gate2484(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2485(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2486(.a(G251), .O(gate236inter7));
  inv1  gate2487(.a(G727), .O(gate236inter8));
  nand2 gate2488(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2489(.a(s_277), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2490(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2491(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2492(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate547(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate548(.a(gate238inter0), .b(s_0), .O(gate238inter1));
  and2  gate549(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate550(.a(s_0), .O(gate238inter3));
  inv1  gate551(.a(s_1), .O(gate238inter4));
  nand2 gate552(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate553(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate554(.a(G257), .O(gate238inter7));
  inv1  gate555(.a(G709), .O(gate238inter8));
  nand2 gate556(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate557(.a(s_1), .b(gate238inter3), .O(gate238inter10));
  nor2  gate558(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate559(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate560(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1611(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1612(.a(gate239inter0), .b(s_152), .O(gate239inter1));
  and2  gate1613(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1614(.a(s_152), .O(gate239inter3));
  inv1  gate1615(.a(s_153), .O(gate239inter4));
  nand2 gate1616(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1617(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1618(.a(G260), .O(gate239inter7));
  inv1  gate1619(.a(G712), .O(gate239inter8));
  nand2 gate1620(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1621(.a(s_153), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1622(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1623(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1624(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate3081(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate3082(.a(gate240inter0), .b(s_362), .O(gate240inter1));
  and2  gate3083(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate3084(.a(s_362), .O(gate240inter3));
  inv1  gate3085(.a(s_363), .O(gate240inter4));
  nand2 gate3086(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate3087(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate3088(.a(G263), .O(gate240inter7));
  inv1  gate3089(.a(G715), .O(gate240inter8));
  nand2 gate3090(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate3091(.a(s_363), .b(gate240inter3), .O(gate240inter10));
  nor2  gate3092(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate3093(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate3094(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1191(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1192(.a(gate243inter0), .b(s_92), .O(gate243inter1));
  and2  gate1193(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1194(.a(s_92), .O(gate243inter3));
  inv1  gate1195(.a(s_93), .O(gate243inter4));
  nand2 gate1196(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1197(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1198(.a(G245), .O(gate243inter7));
  inv1  gate1199(.a(G733), .O(gate243inter8));
  nand2 gate1200(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1201(.a(s_93), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1202(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1203(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1204(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate3025(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate3026(.a(gate244inter0), .b(s_354), .O(gate244inter1));
  and2  gate3027(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate3028(.a(s_354), .O(gate244inter3));
  inv1  gate3029(.a(s_355), .O(gate244inter4));
  nand2 gate3030(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate3031(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate3032(.a(G721), .O(gate244inter7));
  inv1  gate3033(.a(G733), .O(gate244inter8));
  nand2 gate3034(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate3035(.a(s_355), .b(gate244inter3), .O(gate244inter10));
  nor2  gate3036(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate3037(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate3038(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate3109(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate3110(.a(gate245inter0), .b(s_366), .O(gate245inter1));
  and2  gate3111(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate3112(.a(s_366), .O(gate245inter3));
  inv1  gate3113(.a(s_367), .O(gate245inter4));
  nand2 gate3114(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate3115(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate3116(.a(G248), .O(gate245inter7));
  inv1  gate3117(.a(G736), .O(gate245inter8));
  nand2 gate3118(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate3119(.a(s_367), .b(gate245inter3), .O(gate245inter10));
  nor2  gate3120(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate3121(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate3122(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2773(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2774(.a(gate246inter0), .b(s_318), .O(gate246inter1));
  and2  gate2775(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2776(.a(s_318), .O(gate246inter3));
  inv1  gate2777(.a(s_319), .O(gate246inter4));
  nand2 gate2778(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2779(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2780(.a(G724), .O(gate246inter7));
  inv1  gate2781(.a(G736), .O(gate246inter8));
  nand2 gate2782(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2783(.a(s_319), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2784(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2785(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2786(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2353(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2354(.a(gate248inter0), .b(s_258), .O(gate248inter1));
  and2  gate2355(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2356(.a(s_258), .O(gate248inter3));
  inv1  gate2357(.a(s_259), .O(gate248inter4));
  nand2 gate2358(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2359(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2360(.a(G727), .O(gate248inter7));
  inv1  gate2361(.a(G739), .O(gate248inter8));
  nand2 gate2362(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2363(.a(s_259), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2364(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2365(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2366(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate3235(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate3236(.a(gate254inter0), .b(s_384), .O(gate254inter1));
  and2  gate3237(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate3238(.a(s_384), .O(gate254inter3));
  inv1  gate3239(.a(s_385), .O(gate254inter4));
  nand2 gate3240(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate3241(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate3242(.a(G712), .O(gate254inter7));
  inv1  gate3243(.a(G748), .O(gate254inter8));
  nand2 gate3244(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate3245(.a(s_385), .b(gate254inter3), .O(gate254inter10));
  nor2  gate3246(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate3247(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate3248(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1751(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1752(.a(gate258inter0), .b(s_172), .O(gate258inter1));
  and2  gate1753(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1754(.a(s_172), .O(gate258inter3));
  inv1  gate1755(.a(s_173), .O(gate258inter4));
  nand2 gate1756(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1757(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1758(.a(G756), .O(gate258inter7));
  inv1  gate1759(.a(G757), .O(gate258inter8));
  nand2 gate1760(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1761(.a(s_173), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1762(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1763(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1764(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate561(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate562(.a(gate259inter0), .b(s_2), .O(gate259inter1));
  and2  gate563(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate564(.a(s_2), .O(gate259inter3));
  inv1  gate565(.a(s_3), .O(gate259inter4));
  nand2 gate566(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate567(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate568(.a(G758), .O(gate259inter7));
  inv1  gate569(.a(G759), .O(gate259inter8));
  nand2 gate570(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate571(.a(s_3), .b(gate259inter3), .O(gate259inter10));
  nor2  gate572(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate573(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate574(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate3011(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate3012(.a(gate261inter0), .b(s_352), .O(gate261inter1));
  and2  gate3013(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate3014(.a(s_352), .O(gate261inter3));
  inv1  gate3015(.a(s_353), .O(gate261inter4));
  nand2 gate3016(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate3017(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate3018(.a(G762), .O(gate261inter7));
  inv1  gate3019(.a(G763), .O(gate261inter8));
  nand2 gate3020(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate3021(.a(s_353), .b(gate261inter3), .O(gate261inter10));
  nor2  gate3022(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate3023(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate3024(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate2087(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2088(.a(gate266inter0), .b(s_220), .O(gate266inter1));
  and2  gate2089(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2090(.a(s_220), .O(gate266inter3));
  inv1  gate2091(.a(s_221), .O(gate266inter4));
  nand2 gate2092(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2093(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2094(.a(G645), .O(gate266inter7));
  inv1  gate2095(.a(G773), .O(gate266inter8));
  nand2 gate2096(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2097(.a(s_221), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2098(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2099(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2100(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1303(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1304(.a(gate267inter0), .b(s_108), .O(gate267inter1));
  and2  gate1305(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1306(.a(s_108), .O(gate267inter3));
  inv1  gate1307(.a(s_109), .O(gate267inter4));
  nand2 gate1308(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1309(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1310(.a(G648), .O(gate267inter7));
  inv1  gate1311(.a(G776), .O(gate267inter8));
  nand2 gate1312(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1313(.a(s_109), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1314(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1315(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1316(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2591(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2592(.a(gate268inter0), .b(s_292), .O(gate268inter1));
  and2  gate2593(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2594(.a(s_292), .O(gate268inter3));
  inv1  gate2595(.a(s_293), .O(gate268inter4));
  nand2 gate2596(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2597(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2598(.a(G651), .O(gate268inter7));
  inv1  gate2599(.a(G779), .O(gate268inter8));
  nand2 gate2600(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2601(.a(s_293), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2602(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2603(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2604(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate3151(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate3152(.a(gate270inter0), .b(s_372), .O(gate270inter1));
  and2  gate3153(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate3154(.a(s_372), .O(gate270inter3));
  inv1  gate3155(.a(s_373), .O(gate270inter4));
  nand2 gate3156(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate3157(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate3158(.a(G657), .O(gate270inter7));
  inv1  gate3159(.a(G785), .O(gate270inter8));
  nand2 gate3160(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate3161(.a(s_373), .b(gate270inter3), .O(gate270inter10));
  nor2  gate3162(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate3163(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate3164(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2885(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2886(.a(gate271inter0), .b(s_334), .O(gate271inter1));
  and2  gate2887(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2888(.a(s_334), .O(gate271inter3));
  inv1  gate2889(.a(s_335), .O(gate271inter4));
  nand2 gate2890(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2891(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2892(.a(G660), .O(gate271inter7));
  inv1  gate2893(.a(G788), .O(gate271inter8));
  nand2 gate2894(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2895(.a(s_335), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2896(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2897(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2898(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2255(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2256(.a(gate273inter0), .b(s_244), .O(gate273inter1));
  and2  gate2257(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2258(.a(s_244), .O(gate273inter3));
  inv1  gate2259(.a(s_245), .O(gate273inter4));
  nand2 gate2260(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2261(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2262(.a(G642), .O(gate273inter7));
  inv1  gate2263(.a(G794), .O(gate273inter8));
  nand2 gate2264(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2265(.a(s_245), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2266(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2267(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2268(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1513(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1514(.a(gate275inter0), .b(s_138), .O(gate275inter1));
  and2  gate1515(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1516(.a(s_138), .O(gate275inter3));
  inv1  gate1517(.a(s_139), .O(gate275inter4));
  nand2 gate1518(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1519(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1520(.a(G645), .O(gate275inter7));
  inv1  gate1521(.a(G797), .O(gate275inter8));
  nand2 gate1522(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1523(.a(s_139), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1524(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1525(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1526(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate2731(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2732(.a(gate276inter0), .b(s_312), .O(gate276inter1));
  and2  gate2733(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2734(.a(s_312), .O(gate276inter3));
  inv1  gate2735(.a(s_313), .O(gate276inter4));
  nand2 gate2736(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2737(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2738(.a(G773), .O(gate276inter7));
  inv1  gate2739(.a(G797), .O(gate276inter8));
  nand2 gate2740(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2741(.a(s_313), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2742(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2743(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2744(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1793(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1794(.a(gate277inter0), .b(s_178), .O(gate277inter1));
  and2  gate1795(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1796(.a(s_178), .O(gate277inter3));
  inv1  gate1797(.a(s_179), .O(gate277inter4));
  nand2 gate1798(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1799(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1800(.a(G648), .O(gate277inter7));
  inv1  gate1801(.a(G800), .O(gate277inter8));
  nand2 gate1802(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1803(.a(s_179), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1804(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1805(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1806(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate967(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate968(.a(gate280inter0), .b(s_60), .O(gate280inter1));
  and2  gate969(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate970(.a(s_60), .O(gate280inter3));
  inv1  gate971(.a(s_61), .O(gate280inter4));
  nand2 gate972(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate973(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate974(.a(G779), .O(gate280inter7));
  inv1  gate975(.a(G803), .O(gate280inter8));
  nand2 gate976(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate977(.a(s_61), .b(gate280inter3), .O(gate280inter10));
  nor2  gate978(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate979(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate980(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1821(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1822(.a(gate283inter0), .b(s_182), .O(gate283inter1));
  and2  gate1823(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1824(.a(s_182), .O(gate283inter3));
  inv1  gate1825(.a(s_183), .O(gate283inter4));
  nand2 gate1826(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1827(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1828(.a(G657), .O(gate283inter7));
  inv1  gate1829(.a(G809), .O(gate283inter8));
  nand2 gate1830(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1831(.a(s_183), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1832(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1833(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1834(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1569(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1570(.a(gate286inter0), .b(s_146), .O(gate286inter1));
  and2  gate1571(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1572(.a(s_146), .O(gate286inter3));
  inv1  gate1573(.a(s_147), .O(gate286inter4));
  nand2 gate1574(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1575(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1576(.a(G788), .O(gate286inter7));
  inv1  gate1577(.a(G812), .O(gate286inter8));
  nand2 gate1578(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1579(.a(s_147), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1580(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1581(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1582(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2059(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2060(.a(gate287inter0), .b(s_216), .O(gate287inter1));
  and2  gate2061(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2062(.a(s_216), .O(gate287inter3));
  inv1  gate2063(.a(s_217), .O(gate287inter4));
  nand2 gate2064(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2065(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2066(.a(G663), .O(gate287inter7));
  inv1  gate2067(.a(G815), .O(gate287inter8));
  nand2 gate2068(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2069(.a(s_217), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2070(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2071(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2072(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate3137(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate3138(.a(gate288inter0), .b(s_370), .O(gate288inter1));
  and2  gate3139(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate3140(.a(s_370), .O(gate288inter3));
  inv1  gate3141(.a(s_371), .O(gate288inter4));
  nand2 gate3142(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate3143(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate3144(.a(G791), .O(gate288inter7));
  inv1  gate3145(.a(G815), .O(gate288inter8));
  nand2 gate3146(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate3147(.a(s_371), .b(gate288inter3), .O(gate288inter10));
  nor2  gate3148(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate3149(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate3150(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate3207(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate3208(.a(gate289inter0), .b(s_380), .O(gate289inter1));
  and2  gate3209(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate3210(.a(s_380), .O(gate289inter3));
  inv1  gate3211(.a(s_381), .O(gate289inter4));
  nand2 gate3212(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate3213(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate3214(.a(G818), .O(gate289inter7));
  inv1  gate3215(.a(G819), .O(gate289inter8));
  nand2 gate3216(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate3217(.a(s_381), .b(gate289inter3), .O(gate289inter10));
  nor2  gate3218(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate3219(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate3220(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2381(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2382(.a(gate291inter0), .b(s_262), .O(gate291inter1));
  and2  gate2383(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2384(.a(s_262), .O(gate291inter3));
  inv1  gate2385(.a(s_263), .O(gate291inter4));
  nand2 gate2386(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2387(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2388(.a(G822), .O(gate291inter7));
  inv1  gate2389(.a(G823), .O(gate291inter8));
  nand2 gate2390(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2391(.a(s_263), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2392(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2393(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2394(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1835(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1836(.a(gate292inter0), .b(s_184), .O(gate292inter1));
  and2  gate1837(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1838(.a(s_184), .O(gate292inter3));
  inv1  gate1839(.a(s_185), .O(gate292inter4));
  nand2 gate1840(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1841(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1842(.a(G824), .O(gate292inter7));
  inv1  gate1843(.a(G825), .O(gate292inter8));
  nand2 gate1844(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1845(.a(s_185), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1846(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1847(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1848(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2031(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2032(.a(gate294inter0), .b(s_212), .O(gate294inter1));
  and2  gate2033(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2034(.a(s_212), .O(gate294inter3));
  inv1  gate2035(.a(s_213), .O(gate294inter4));
  nand2 gate2036(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2037(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2038(.a(G832), .O(gate294inter7));
  inv1  gate2039(.a(G833), .O(gate294inter8));
  nand2 gate2040(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2041(.a(s_213), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2042(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2043(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2044(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1737(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1738(.a(gate296inter0), .b(s_170), .O(gate296inter1));
  and2  gate1739(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1740(.a(s_170), .O(gate296inter3));
  inv1  gate1741(.a(s_171), .O(gate296inter4));
  nand2 gate1742(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1743(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1744(.a(G826), .O(gate296inter7));
  inv1  gate1745(.a(G827), .O(gate296inter8));
  nand2 gate1746(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1747(.a(s_171), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1748(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1749(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1750(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1723(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1724(.a(gate387inter0), .b(s_168), .O(gate387inter1));
  and2  gate1725(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1726(.a(s_168), .O(gate387inter3));
  inv1  gate1727(.a(s_169), .O(gate387inter4));
  nand2 gate1728(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1729(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1730(.a(G1), .O(gate387inter7));
  inv1  gate1731(.a(G1036), .O(gate387inter8));
  nand2 gate1732(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1733(.a(s_169), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1734(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1735(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1736(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2633(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2634(.a(gate391inter0), .b(s_298), .O(gate391inter1));
  and2  gate2635(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2636(.a(s_298), .O(gate391inter3));
  inv1  gate2637(.a(s_299), .O(gate391inter4));
  nand2 gate2638(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2639(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2640(.a(G5), .O(gate391inter7));
  inv1  gate2641(.a(G1048), .O(gate391inter8));
  nand2 gate2642(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2643(.a(s_299), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2644(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2645(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2646(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1247(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1248(.a(gate392inter0), .b(s_100), .O(gate392inter1));
  and2  gate1249(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1250(.a(s_100), .O(gate392inter3));
  inv1  gate1251(.a(s_101), .O(gate392inter4));
  nand2 gate1252(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1253(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1254(.a(G6), .O(gate392inter7));
  inv1  gate1255(.a(G1051), .O(gate392inter8));
  nand2 gate1256(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1257(.a(s_101), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1258(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1259(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1260(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate3067(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate3068(.a(gate393inter0), .b(s_360), .O(gate393inter1));
  and2  gate3069(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate3070(.a(s_360), .O(gate393inter3));
  inv1  gate3071(.a(s_361), .O(gate393inter4));
  nand2 gate3072(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate3073(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate3074(.a(G7), .O(gate393inter7));
  inv1  gate3075(.a(G1054), .O(gate393inter8));
  nand2 gate3076(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate3077(.a(s_361), .b(gate393inter3), .O(gate393inter10));
  nor2  gate3078(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate3079(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate3080(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1037(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1038(.a(gate397inter0), .b(s_70), .O(gate397inter1));
  and2  gate1039(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1040(.a(s_70), .O(gate397inter3));
  inv1  gate1041(.a(s_71), .O(gate397inter4));
  nand2 gate1042(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1043(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1044(.a(G11), .O(gate397inter7));
  inv1  gate1045(.a(G1066), .O(gate397inter8));
  nand2 gate1046(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1047(.a(s_71), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1048(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1049(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1050(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1961(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1962(.a(gate398inter0), .b(s_202), .O(gate398inter1));
  and2  gate1963(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1964(.a(s_202), .O(gate398inter3));
  inv1  gate1965(.a(s_203), .O(gate398inter4));
  nand2 gate1966(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1967(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1968(.a(G12), .O(gate398inter7));
  inv1  gate1969(.a(G1069), .O(gate398inter8));
  nand2 gate1970(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1971(.a(s_203), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1972(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1973(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1974(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate2213(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2214(.a(gate399inter0), .b(s_238), .O(gate399inter1));
  and2  gate2215(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2216(.a(s_238), .O(gate399inter3));
  inv1  gate2217(.a(s_239), .O(gate399inter4));
  nand2 gate2218(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2219(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2220(.a(G13), .O(gate399inter7));
  inv1  gate2221(.a(G1072), .O(gate399inter8));
  nand2 gate2222(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2223(.a(s_239), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2224(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2225(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2226(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2311(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2312(.a(gate400inter0), .b(s_252), .O(gate400inter1));
  and2  gate2313(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2314(.a(s_252), .O(gate400inter3));
  inv1  gate2315(.a(s_253), .O(gate400inter4));
  nand2 gate2316(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2317(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2318(.a(G14), .O(gate400inter7));
  inv1  gate2319(.a(G1075), .O(gate400inter8));
  nand2 gate2320(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2321(.a(s_253), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2322(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2323(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2324(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1933(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1934(.a(gate402inter0), .b(s_198), .O(gate402inter1));
  and2  gate1935(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1936(.a(s_198), .O(gate402inter3));
  inv1  gate1937(.a(s_199), .O(gate402inter4));
  nand2 gate1938(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1939(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1940(.a(G16), .O(gate402inter7));
  inv1  gate1941(.a(G1081), .O(gate402inter8));
  nand2 gate1942(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1943(.a(s_199), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1944(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1945(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1946(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate3039(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate3040(.a(gate404inter0), .b(s_356), .O(gate404inter1));
  and2  gate3041(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate3042(.a(s_356), .O(gate404inter3));
  inv1  gate3043(.a(s_357), .O(gate404inter4));
  nand2 gate3044(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate3045(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate3046(.a(G18), .O(gate404inter7));
  inv1  gate3047(.a(G1087), .O(gate404inter8));
  nand2 gate3048(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate3049(.a(s_357), .b(gate404inter3), .O(gate404inter10));
  nor2  gate3050(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate3051(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate3052(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1863(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1864(.a(gate405inter0), .b(s_188), .O(gate405inter1));
  and2  gate1865(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1866(.a(s_188), .O(gate405inter3));
  inv1  gate1867(.a(s_189), .O(gate405inter4));
  nand2 gate1868(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1869(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1870(.a(G19), .O(gate405inter7));
  inv1  gate1871(.a(G1090), .O(gate405inter8));
  nand2 gate1872(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1873(.a(s_189), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1874(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1875(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1876(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate3277(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate3278(.a(gate406inter0), .b(s_390), .O(gate406inter1));
  and2  gate3279(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate3280(.a(s_390), .O(gate406inter3));
  inv1  gate3281(.a(s_391), .O(gate406inter4));
  nand2 gate3282(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate3283(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate3284(.a(G20), .O(gate406inter7));
  inv1  gate3285(.a(G1093), .O(gate406inter8));
  nand2 gate3286(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate3287(.a(s_391), .b(gate406inter3), .O(gate406inter10));
  nor2  gate3288(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate3289(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate3290(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate883(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate884(.a(gate409inter0), .b(s_48), .O(gate409inter1));
  and2  gate885(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate886(.a(s_48), .O(gate409inter3));
  inv1  gate887(.a(s_49), .O(gate409inter4));
  nand2 gate888(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate889(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate890(.a(G23), .O(gate409inter7));
  inv1  gate891(.a(G1102), .O(gate409inter8));
  nand2 gate892(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate893(.a(s_49), .b(gate409inter3), .O(gate409inter10));
  nor2  gate894(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate895(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate896(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate841(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate842(.a(gate410inter0), .b(s_42), .O(gate410inter1));
  and2  gate843(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate844(.a(s_42), .O(gate410inter3));
  inv1  gate845(.a(s_43), .O(gate410inter4));
  nand2 gate846(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate847(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate848(.a(G24), .O(gate410inter7));
  inv1  gate849(.a(G1105), .O(gate410inter8));
  nand2 gate850(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate851(.a(s_43), .b(gate410inter3), .O(gate410inter10));
  nor2  gate852(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate853(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate854(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate939(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate940(.a(gate412inter0), .b(s_56), .O(gate412inter1));
  and2  gate941(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate942(.a(s_56), .O(gate412inter3));
  inv1  gate943(.a(s_57), .O(gate412inter4));
  nand2 gate944(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate945(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate946(.a(G26), .O(gate412inter7));
  inv1  gate947(.a(G1111), .O(gate412inter8));
  nand2 gate948(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate949(.a(s_57), .b(gate412inter3), .O(gate412inter10));
  nor2  gate950(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate951(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate952(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1233(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1234(.a(gate413inter0), .b(s_98), .O(gate413inter1));
  and2  gate1235(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1236(.a(s_98), .O(gate413inter3));
  inv1  gate1237(.a(s_99), .O(gate413inter4));
  nand2 gate1238(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1239(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1240(.a(G27), .O(gate413inter7));
  inv1  gate1241(.a(G1114), .O(gate413inter8));
  nand2 gate1242(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1243(.a(s_99), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1244(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1245(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1246(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1947(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1948(.a(gate414inter0), .b(s_200), .O(gate414inter1));
  and2  gate1949(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1950(.a(s_200), .O(gate414inter3));
  inv1  gate1951(.a(s_201), .O(gate414inter4));
  nand2 gate1952(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1953(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1954(.a(G28), .O(gate414inter7));
  inv1  gate1955(.a(G1117), .O(gate414inter8));
  nand2 gate1956(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1957(.a(s_201), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1958(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1959(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1960(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1555(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1556(.a(gate417inter0), .b(s_144), .O(gate417inter1));
  and2  gate1557(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1558(.a(s_144), .O(gate417inter3));
  inv1  gate1559(.a(s_145), .O(gate417inter4));
  nand2 gate1560(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1561(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1562(.a(G31), .O(gate417inter7));
  inv1  gate1563(.a(G1126), .O(gate417inter8));
  nand2 gate1564(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1565(.a(s_145), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1566(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1567(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1568(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2283(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2284(.a(gate418inter0), .b(s_248), .O(gate418inter1));
  and2  gate2285(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2286(.a(s_248), .O(gate418inter3));
  inv1  gate2287(.a(s_249), .O(gate418inter4));
  nand2 gate2288(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2289(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2290(.a(G32), .O(gate418inter7));
  inv1  gate2291(.a(G1129), .O(gate418inter8));
  nand2 gate2292(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2293(.a(s_249), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2294(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2295(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2296(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate3291(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate3292(.a(gate419inter0), .b(s_392), .O(gate419inter1));
  and2  gate3293(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate3294(.a(s_392), .O(gate419inter3));
  inv1  gate3295(.a(s_393), .O(gate419inter4));
  nand2 gate3296(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate3297(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate3298(.a(G1), .O(gate419inter7));
  inv1  gate3299(.a(G1132), .O(gate419inter8));
  nand2 gate3300(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate3301(.a(s_393), .b(gate419inter3), .O(gate419inter10));
  nor2  gate3302(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate3303(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate3304(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate617(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate618(.a(gate422inter0), .b(s_10), .O(gate422inter1));
  and2  gate619(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate620(.a(s_10), .O(gate422inter3));
  inv1  gate621(.a(s_11), .O(gate422inter4));
  nand2 gate622(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate623(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate624(.a(G1039), .O(gate422inter7));
  inv1  gate625(.a(G1135), .O(gate422inter8));
  nand2 gate626(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate627(.a(s_11), .b(gate422inter3), .O(gate422inter10));
  nor2  gate628(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate629(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate630(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1695(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1696(.a(gate423inter0), .b(s_164), .O(gate423inter1));
  and2  gate1697(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1698(.a(s_164), .O(gate423inter3));
  inv1  gate1699(.a(s_165), .O(gate423inter4));
  nand2 gate1700(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1701(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1702(.a(G3), .O(gate423inter7));
  inv1  gate1703(.a(G1138), .O(gate423inter8));
  nand2 gate1704(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1705(.a(s_165), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1706(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1707(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1708(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2899(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2900(.a(gate424inter0), .b(s_336), .O(gate424inter1));
  and2  gate2901(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2902(.a(s_336), .O(gate424inter3));
  inv1  gate2903(.a(s_337), .O(gate424inter4));
  nand2 gate2904(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2905(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2906(.a(G1042), .O(gate424inter7));
  inv1  gate2907(.a(G1138), .O(gate424inter8));
  nand2 gate2908(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2909(.a(s_337), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2910(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2911(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2912(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate3305(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate3306(.a(gate428inter0), .b(s_394), .O(gate428inter1));
  and2  gate3307(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate3308(.a(s_394), .O(gate428inter3));
  inv1  gate3309(.a(s_395), .O(gate428inter4));
  nand2 gate3310(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate3311(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate3312(.a(G1048), .O(gate428inter7));
  inv1  gate3313(.a(G1144), .O(gate428inter8));
  nand2 gate3314(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate3315(.a(s_395), .b(gate428inter3), .O(gate428inter10));
  nor2  gate3316(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate3317(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate3318(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2297(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2298(.a(gate431inter0), .b(s_250), .O(gate431inter1));
  and2  gate2299(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2300(.a(s_250), .O(gate431inter3));
  inv1  gate2301(.a(s_251), .O(gate431inter4));
  nand2 gate2302(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2303(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2304(.a(G7), .O(gate431inter7));
  inv1  gate2305(.a(G1150), .O(gate431inter8));
  nand2 gate2306(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2307(.a(s_251), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2308(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2309(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2310(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2493(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2494(.a(gate432inter0), .b(s_278), .O(gate432inter1));
  and2  gate2495(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2496(.a(s_278), .O(gate432inter3));
  inv1  gate2497(.a(s_279), .O(gate432inter4));
  nand2 gate2498(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2499(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2500(.a(G1054), .O(gate432inter7));
  inv1  gate2501(.a(G1150), .O(gate432inter8));
  nand2 gate2502(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2503(.a(s_279), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2504(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2505(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2506(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate3333(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate3334(.a(gate433inter0), .b(s_398), .O(gate433inter1));
  and2  gate3335(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate3336(.a(s_398), .O(gate433inter3));
  inv1  gate3337(.a(s_399), .O(gate433inter4));
  nand2 gate3338(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate3339(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate3340(.a(G8), .O(gate433inter7));
  inv1  gate3341(.a(G1153), .O(gate433inter8));
  nand2 gate3342(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate3343(.a(s_399), .b(gate433inter3), .O(gate433inter10));
  nor2  gate3344(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate3345(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate3346(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1163(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1164(.a(gate434inter0), .b(s_88), .O(gate434inter1));
  and2  gate1165(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1166(.a(s_88), .O(gate434inter3));
  inv1  gate1167(.a(s_89), .O(gate434inter4));
  nand2 gate1168(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1169(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1170(.a(G1057), .O(gate434inter7));
  inv1  gate1171(.a(G1153), .O(gate434inter8));
  nand2 gate1172(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1173(.a(s_89), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1174(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1175(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1176(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate2409(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2410(.a(gate436inter0), .b(s_266), .O(gate436inter1));
  and2  gate2411(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2412(.a(s_266), .O(gate436inter3));
  inv1  gate2413(.a(s_267), .O(gate436inter4));
  nand2 gate2414(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2415(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2416(.a(G1060), .O(gate436inter7));
  inv1  gate2417(.a(G1156), .O(gate436inter8));
  nand2 gate2418(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2419(.a(s_267), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2420(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2421(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2422(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate2801(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2802(.a(gate437inter0), .b(s_322), .O(gate437inter1));
  and2  gate2803(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2804(.a(s_322), .O(gate437inter3));
  inv1  gate2805(.a(s_323), .O(gate437inter4));
  nand2 gate2806(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2807(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2808(.a(G10), .O(gate437inter7));
  inv1  gate2809(.a(G1159), .O(gate437inter8));
  nand2 gate2810(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2811(.a(s_323), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2812(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2813(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2814(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate3347(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate3348(.a(gate439inter0), .b(s_400), .O(gate439inter1));
  and2  gate3349(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate3350(.a(s_400), .O(gate439inter3));
  inv1  gate3351(.a(s_401), .O(gate439inter4));
  nand2 gate3352(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate3353(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate3354(.a(G11), .O(gate439inter7));
  inv1  gate3355(.a(G1162), .O(gate439inter8));
  nand2 gate3356(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate3357(.a(s_401), .b(gate439inter3), .O(gate439inter10));
  nor2  gate3358(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate3359(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate3360(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2577(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2578(.a(gate442inter0), .b(s_290), .O(gate442inter1));
  and2  gate2579(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2580(.a(s_290), .O(gate442inter3));
  inv1  gate2581(.a(s_291), .O(gate442inter4));
  nand2 gate2582(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2583(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2584(.a(G1069), .O(gate442inter7));
  inv1  gate2585(.a(G1165), .O(gate442inter8));
  nand2 gate2586(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2587(.a(s_291), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2588(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2589(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2590(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1639(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1640(.a(gate445inter0), .b(s_156), .O(gate445inter1));
  and2  gate1641(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1642(.a(s_156), .O(gate445inter3));
  inv1  gate1643(.a(s_157), .O(gate445inter4));
  nand2 gate1644(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1645(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1646(.a(G14), .O(gate445inter7));
  inv1  gate1647(.a(G1171), .O(gate445inter8));
  nand2 gate1648(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1649(.a(s_157), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1650(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1651(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1652(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate3193(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate3194(.a(gate446inter0), .b(s_378), .O(gate446inter1));
  and2  gate3195(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate3196(.a(s_378), .O(gate446inter3));
  inv1  gate3197(.a(s_379), .O(gate446inter4));
  nand2 gate3198(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate3199(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate3200(.a(G1075), .O(gate446inter7));
  inv1  gate3201(.a(G1171), .O(gate446inter8));
  nand2 gate3202(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate3203(.a(s_379), .b(gate446inter3), .O(gate446inter10));
  nor2  gate3204(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate3205(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate3206(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1975(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1976(.a(gate447inter0), .b(s_204), .O(gate447inter1));
  and2  gate1977(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1978(.a(s_204), .O(gate447inter3));
  inv1  gate1979(.a(s_205), .O(gate447inter4));
  nand2 gate1980(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1981(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1982(.a(G15), .O(gate447inter7));
  inv1  gate1983(.a(G1174), .O(gate447inter8));
  nand2 gate1984(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1985(.a(s_205), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1986(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1987(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1988(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2913(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2914(.a(gate448inter0), .b(s_338), .O(gate448inter1));
  and2  gate2915(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2916(.a(s_338), .O(gate448inter3));
  inv1  gate2917(.a(s_339), .O(gate448inter4));
  nand2 gate2918(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2919(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2920(.a(G1078), .O(gate448inter7));
  inv1  gate2921(.a(G1174), .O(gate448inter8));
  nand2 gate2922(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2923(.a(s_339), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2924(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2925(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2926(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2717(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2718(.a(gate451inter0), .b(s_310), .O(gate451inter1));
  and2  gate2719(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2720(.a(s_310), .O(gate451inter3));
  inv1  gate2721(.a(s_311), .O(gate451inter4));
  nand2 gate2722(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2723(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2724(.a(G17), .O(gate451inter7));
  inv1  gate2725(.a(G1180), .O(gate451inter8));
  nand2 gate2726(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2727(.a(s_311), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2728(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2729(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2730(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1849(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1850(.a(gate454inter0), .b(s_186), .O(gate454inter1));
  and2  gate1851(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1852(.a(s_186), .O(gate454inter3));
  inv1  gate1853(.a(s_187), .O(gate454inter4));
  nand2 gate1854(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1855(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1856(.a(G1087), .O(gate454inter7));
  inv1  gate1857(.a(G1183), .O(gate454inter8));
  nand2 gate1858(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1859(.a(s_187), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1860(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1861(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1862(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2955(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2956(.a(gate461inter0), .b(s_344), .O(gate461inter1));
  and2  gate2957(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2958(.a(s_344), .O(gate461inter3));
  inv1  gate2959(.a(s_345), .O(gate461inter4));
  nand2 gate2960(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2961(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2962(.a(G22), .O(gate461inter7));
  inv1  gate2963(.a(G1195), .O(gate461inter8));
  nand2 gate2964(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2965(.a(s_345), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2966(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2967(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2968(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate855(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate856(.a(gate462inter0), .b(s_44), .O(gate462inter1));
  and2  gate857(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate858(.a(s_44), .O(gate462inter3));
  inv1  gate859(.a(s_45), .O(gate462inter4));
  nand2 gate860(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate861(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate862(.a(G1099), .O(gate462inter7));
  inv1  gate863(.a(G1195), .O(gate462inter8));
  nand2 gate864(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate865(.a(s_45), .b(gate462inter3), .O(gate462inter10));
  nor2  gate866(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate867(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate868(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2199(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2200(.a(gate465inter0), .b(s_236), .O(gate465inter1));
  and2  gate2201(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2202(.a(s_236), .O(gate465inter3));
  inv1  gate2203(.a(s_237), .O(gate465inter4));
  nand2 gate2204(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2205(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2206(.a(G24), .O(gate465inter7));
  inv1  gate2207(.a(G1201), .O(gate465inter8));
  nand2 gate2208(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2209(.a(s_237), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2210(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2211(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2212(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1149(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1150(.a(gate467inter0), .b(s_86), .O(gate467inter1));
  and2  gate1151(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1152(.a(s_86), .O(gate467inter3));
  inv1  gate1153(.a(s_87), .O(gate467inter4));
  nand2 gate1154(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1155(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1156(.a(G25), .O(gate467inter7));
  inv1  gate1157(.a(G1204), .O(gate467inter8));
  nand2 gate1158(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1159(.a(s_87), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1160(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1161(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1162(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1471(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1472(.a(gate468inter0), .b(s_132), .O(gate468inter1));
  and2  gate1473(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1474(.a(s_132), .O(gate468inter3));
  inv1  gate1475(.a(s_133), .O(gate468inter4));
  nand2 gate1476(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1477(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1478(.a(G1108), .O(gate468inter7));
  inv1  gate1479(.a(G1204), .O(gate468inter8));
  nand2 gate1480(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1481(.a(s_133), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1482(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1483(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1484(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1387(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1388(.a(gate471inter0), .b(s_120), .O(gate471inter1));
  and2  gate1389(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1390(.a(s_120), .O(gate471inter3));
  inv1  gate1391(.a(s_121), .O(gate471inter4));
  nand2 gate1392(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1393(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1394(.a(G27), .O(gate471inter7));
  inv1  gate1395(.a(G1210), .O(gate471inter8));
  nand2 gate1396(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1397(.a(s_121), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1398(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1399(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1400(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2829(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2830(.a(gate475inter0), .b(s_326), .O(gate475inter1));
  and2  gate2831(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2832(.a(s_326), .O(gate475inter3));
  inv1  gate2833(.a(s_327), .O(gate475inter4));
  nand2 gate2834(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2835(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2836(.a(G29), .O(gate475inter7));
  inv1  gate2837(.a(G1216), .O(gate475inter8));
  nand2 gate2838(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2839(.a(s_327), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2840(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2841(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2842(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2745(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2746(.a(gate477inter0), .b(s_314), .O(gate477inter1));
  and2  gate2747(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2748(.a(s_314), .O(gate477inter3));
  inv1  gate2749(.a(s_315), .O(gate477inter4));
  nand2 gate2750(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2751(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2752(.a(G30), .O(gate477inter7));
  inv1  gate2753(.a(G1219), .O(gate477inter8));
  nand2 gate2754(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2755(.a(s_315), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2756(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2757(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2758(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2703(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2704(.a(gate479inter0), .b(s_308), .O(gate479inter1));
  and2  gate2705(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2706(.a(s_308), .O(gate479inter3));
  inv1  gate2707(.a(s_309), .O(gate479inter4));
  nand2 gate2708(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2709(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2710(.a(G31), .O(gate479inter7));
  inv1  gate2711(.a(G1222), .O(gate479inter8));
  nand2 gate2712(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2713(.a(s_309), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2714(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2715(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2716(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1527(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1528(.a(gate480inter0), .b(s_140), .O(gate480inter1));
  and2  gate1529(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1530(.a(s_140), .O(gate480inter3));
  inv1  gate1531(.a(s_141), .O(gate480inter4));
  nand2 gate1532(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1533(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1534(.a(G1126), .O(gate480inter7));
  inv1  gate1535(.a(G1222), .O(gate480inter8));
  nand2 gate1536(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1537(.a(s_141), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1538(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1539(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1540(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2549(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2550(.a(gate483inter0), .b(s_286), .O(gate483inter1));
  and2  gate2551(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2552(.a(s_286), .O(gate483inter3));
  inv1  gate2553(.a(s_287), .O(gate483inter4));
  nand2 gate2554(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2555(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2556(.a(G1228), .O(gate483inter7));
  inv1  gate2557(.a(G1229), .O(gate483inter8));
  nand2 gate2558(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2559(.a(s_287), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2560(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2561(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2562(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate715(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate716(.a(gate484inter0), .b(s_24), .O(gate484inter1));
  and2  gate717(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate718(.a(s_24), .O(gate484inter3));
  inv1  gate719(.a(s_25), .O(gate484inter4));
  nand2 gate720(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate721(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate722(.a(G1230), .O(gate484inter7));
  inv1  gate723(.a(G1231), .O(gate484inter8));
  nand2 gate724(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate725(.a(s_25), .b(gate484inter3), .O(gate484inter10));
  nor2  gate726(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate727(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate728(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate659(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate660(.a(gate486inter0), .b(s_16), .O(gate486inter1));
  and2  gate661(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate662(.a(s_16), .O(gate486inter3));
  inv1  gate663(.a(s_17), .O(gate486inter4));
  nand2 gate664(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate665(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate666(.a(G1234), .O(gate486inter7));
  inv1  gate667(.a(G1235), .O(gate486inter8));
  nand2 gate668(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate669(.a(s_17), .b(gate486inter3), .O(gate486inter10));
  nor2  gate670(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate671(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate672(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1597(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1598(.a(gate489inter0), .b(s_150), .O(gate489inter1));
  and2  gate1599(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1600(.a(s_150), .O(gate489inter3));
  inv1  gate1601(.a(s_151), .O(gate489inter4));
  nand2 gate1602(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1603(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1604(.a(G1240), .O(gate489inter7));
  inv1  gate1605(.a(G1241), .O(gate489inter8));
  nand2 gate1606(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1607(.a(s_151), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1608(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1609(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1610(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1429(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1430(.a(gate491inter0), .b(s_126), .O(gate491inter1));
  and2  gate1431(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1432(.a(s_126), .O(gate491inter3));
  inv1  gate1433(.a(s_127), .O(gate491inter4));
  nand2 gate1434(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1435(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1436(.a(G1244), .O(gate491inter7));
  inv1  gate1437(.a(G1245), .O(gate491inter8));
  nand2 gate1438(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1439(.a(s_127), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1440(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1441(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1442(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1807(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1808(.a(gate492inter0), .b(s_180), .O(gate492inter1));
  and2  gate1809(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1810(.a(s_180), .O(gate492inter3));
  inv1  gate1811(.a(s_181), .O(gate492inter4));
  nand2 gate1812(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1813(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1814(.a(G1246), .O(gate492inter7));
  inv1  gate1815(.a(G1247), .O(gate492inter8));
  nand2 gate1816(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1817(.a(s_181), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1818(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1819(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1820(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate3095(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate3096(.a(gate493inter0), .b(s_364), .O(gate493inter1));
  and2  gate3097(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate3098(.a(s_364), .O(gate493inter3));
  inv1  gate3099(.a(s_365), .O(gate493inter4));
  nand2 gate3100(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate3101(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate3102(.a(G1248), .O(gate493inter7));
  inv1  gate3103(.a(G1249), .O(gate493inter8));
  nand2 gate3104(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate3105(.a(s_365), .b(gate493inter3), .O(gate493inter10));
  nor2  gate3106(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate3107(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate3108(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1009(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1010(.a(gate494inter0), .b(s_66), .O(gate494inter1));
  and2  gate1011(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1012(.a(s_66), .O(gate494inter3));
  inv1  gate1013(.a(s_67), .O(gate494inter4));
  nand2 gate1014(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1015(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1016(.a(G1250), .O(gate494inter7));
  inv1  gate1017(.a(G1251), .O(gate494inter8));
  nand2 gate1018(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1019(.a(s_67), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1020(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1021(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1022(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1989(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1990(.a(gate496inter0), .b(s_206), .O(gate496inter1));
  and2  gate1991(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1992(.a(s_206), .O(gate496inter3));
  inv1  gate1993(.a(s_207), .O(gate496inter4));
  nand2 gate1994(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1995(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1996(.a(G1254), .O(gate496inter7));
  inv1  gate1997(.a(G1255), .O(gate496inter8));
  nand2 gate1998(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1999(.a(s_207), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2000(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2001(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2002(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate3165(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate3166(.a(gate497inter0), .b(s_374), .O(gate497inter1));
  and2  gate3167(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate3168(.a(s_374), .O(gate497inter3));
  inv1  gate3169(.a(s_375), .O(gate497inter4));
  nand2 gate3170(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate3171(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate3172(.a(G1256), .O(gate497inter7));
  inv1  gate3173(.a(G1257), .O(gate497inter8));
  nand2 gate3174(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate3175(.a(s_375), .b(gate497inter3), .O(gate497inter10));
  nor2  gate3176(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate3177(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate3178(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2269(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2270(.a(gate500inter0), .b(s_246), .O(gate500inter1));
  and2  gate2271(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2272(.a(s_246), .O(gate500inter3));
  inv1  gate2273(.a(s_247), .O(gate500inter4));
  nand2 gate2274(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2275(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2276(.a(G1262), .O(gate500inter7));
  inv1  gate2277(.a(G1263), .O(gate500inter8));
  nand2 gate2278(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2279(.a(s_247), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2280(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2281(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2282(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate645(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate646(.a(gate501inter0), .b(s_14), .O(gate501inter1));
  and2  gate647(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate648(.a(s_14), .O(gate501inter3));
  inv1  gate649(.a(s_15), .O(gate501inter4));
  nand2 gate650(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate651(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate652(.a(G1264), .O(gate501inter7));
  inv1  gate653(.a(G1265), .O(gate501inter8));
  nand2 gate654(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate655(.a(s_15), .b(gate501inter3), .O(gate501inter10));
  nor2  gate656(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate657(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate658(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2101(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2102(.a(gate506inter0), .b(s_222), .O(gate506inter1));
  and2  gate2103(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2104(.a(s_222), .O(gate506inter3));
  inv1  gate2105(.a(s_223), .O(gate506inter4));
  nand2 gate2106(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2107(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2108(.a(G1274), .O(gate506inter7));
  inv1  gate2109(.a(G1275), .O(gate506inter8));
  nand2 gate2110(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2111(.a(s_223), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2112(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2113(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2114(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2129(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2130(.a(gate513inter0), .b(s_226), .O(gate513inter1));
  and2  gate2131(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2132(.a(s_226), .O(gate513inter3));
  inv1  gate2133(.a(s_227), .O(gate513inter4));
  nand2 gate2134(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2135(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2136(.a(G1288), .O(gate513inter7));
  inv1  gate2137(.a(G1289), .O(gate513inter8));
  nand2 gate2138(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2139(.a(s_227), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2140(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2141(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2142(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule