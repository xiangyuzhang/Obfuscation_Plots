module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate757(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate758(.a(gate12inter0), .b(s_30), .O(gate12inter1));
  and2  gate759(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate760(.a(s_30), .O(gate12inter3));
  inv1  gate761(.a(s_31), .O(gate12inter4));
  nand2 gate762(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate763(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate764(.a(G7), .O(gate12inter7));
  inv1  gate765(.a(G8), .O(gate12inter8));
  nand2 gate766(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate767(.a(s_31), .b(gate12inter3), .O(gate12inter10));
  nor2  gate768(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate769(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate770(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1233(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1234(.a(gate16inter0), .b(s_98), .O(gate16inter1));
  and2  gate1235(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1236(.a(s_98), .O(gate16inter3));
  inv1  gate1237(.a(s_99), .O(gate16inter4));
  nand2 gate1238(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1239(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1240(.a(G15), .O(gate16inter7));
  inv1  gate1241(.a(G16), .O(gate16inter8));
  nand2 gate1242(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1243(.a(s_99), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1244(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1245(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1246(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1261(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1262(.a(gate36inter0), .b(s_102), .O(gate36inter1));
  and2  gate1263(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1264(.a(s_102), .O(gate36inter3));
  inv1  gate1265(.a(s_103), .O(gate36inter4));
  nand2 gate1266(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1267(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1268(.a(G26), .O(gate36inter7));
  inv1  gate1269(.a(G30), .O(gate36inter8));
  nand2 gate1270(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1271(.a(s_103), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1272(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1273(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1274(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate771(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate772(.a(gate44inter0), .b(s_32), .O(gate44inter1));
  and2  gate773(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate774(.a(s_32), .O(gate44inter3));
  inv1  gate775(.a(s_33), .O(gate44inter4));
  nand2 gate776(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate777(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate778(.a(G4), .O(gate44inter7));
  inv1  gate779(.a(G269), .O(gate44inter8));
  nand2 gate780(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate781(.a(s_33), .b(gate44inter3), .O(gate44inter10));
  nor2  gate782(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate783(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate784(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate617(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate618(.a(gate45inter0), .b(s_10), .O(gate45inter1));
  and2  gate619(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate620(.a(s_10), .O(gate45inter3));
  inv1  gate621(.a(s_11), .O(gate45inter4));
  nand2 gate622(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate623(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate624(.a(G5), .O(gate45inter7));
  inv1  gate625(.a(G272), .O(gate45inter8));
  nand2 gate626(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate627(.a(s_11), .b(gate45inter3), .O(gate45inter10));
  nor2  gate628(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate629(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate630(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1387(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1388(.a(gate52inter0), .b(s_120), .O(gate52inter1));
  and2  gate1389(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1390(.a(s_120), .O(gate52inter3));
  inv1  gate1391(.a(s_121), .O(gate52inter4));
  nand2 gate1392(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1393(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1394(.a(G12), .O(gate52inter7));
  inv1  gate1395(.a(G281), .O(gate52inter8));
  nand2 gate1396(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1397(.a(s_121), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1398(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1399(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1400(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1303(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1304(.a(gate53inter0), .b(s_108), .O(gate53inter1));
  and2  gate1305(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1306(.a(s_108), .O(gate53inter3));
  inv1  gate1307(.a(s_109), .O(gate53inter4));
  nand2 gate1308(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1309(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1310(.a(G13), .O(gate53inter7));
  inv1  gate1311(.a(G284), .O(gate53inter8));
  nand2 gate1312(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1313(.a(s_109), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1314(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1315(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1316(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1135(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1136(.a(gate58inter0), .b(s_84), .O(gate58inter1));
  and2  gate1137(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1138(.a(s_84), .O(gate58inter3));
  inv1  gate1139(.a(s_85), .O(gate58inter4));
  nand2 gate1140(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1141(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1142(.a(G18), .O(gate58inter7));
  inv1  gate1143(.a(G290), .O(gate58inter8));
  nand2 gate1144(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1145(.a(s_85), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1146(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1147(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1148(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1163(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1164(.a(gate81inter0), .b(s_88), .O(gate81inter1));
  and2  gate1165(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1166(.a(s_88), .O(gate81inter3));
  inv1  gate1167(.a(s_89), .O(gate81inter4));
  nand2 gate1168(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1169(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1170(.a(G3), .O(gate81inter7));
  inv1  gate1171(.a(G326), .O(gate81inter8));
  nand2 gate1172(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1173(.a(s_89), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1174(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1175(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1176(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1331(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1332(.a(gate85inter0), .b(s_112), .O(gate85inter1));
  and2  gate1333(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1334(.a(s_112), .O(gate85inter3));
  inv1  gate1335(.a(s_113), .O(gate85inter4));
  nand2 gate1336(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1337(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1338(.a(G4), .O(gate85inter7));
  inv1  gate1339(.a(G332), .O(gate85inter8));
  nand2 gate1340(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1341(.a(s_113), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1342(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1343(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1344(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1359(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1360(.a(gate109inter0), .b(s_116), .O(gate109inter1));
  and2  gate1361(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1362(.a(s_116), .O(gate109inter3));
  inv1  gate1363(.a(s_117), .O(gate109inter4));
  nand2 gate1364(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1365(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1366(.a(G370), .O(gate109inter7));
  inv1  gate1367(.a(G371), .O(gate109inter8));
  nand2 gate1368(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1369(.a(s_117), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1370(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1371(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1372(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1093(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1094(.a(gate111inter0), .b(s_78), .O(gate111inter1));
  and2  gate1095(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1096(.a(s_78), .O(gate111inter3));
  inv1  gate1097(.a(s_79), .O(gate111inter4));
  nand2 gate1098(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1099(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1100(.a(G374), .O(gate111inter7));
  inv1  gate1101(.a(G375), .O(gate111inter8));
  nand2 gate1102(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1103(.a(s_79), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1104(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1105(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1106(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1107(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1108(.a(gate125inter0), .b(s_80), .O(gate125inter1));
  and2  gate1109(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1110(.a(s_80), .O(gate125inter3));
  inv1  gate1111(.a(s_81), .O(gate125inter4));
  nand2 gate1112(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1113(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1114(.a(G402), .O(gate125inter7));
  inv1  gate1115(.a(G403), .O(gate125inter8));
  nand2 gate1116(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1117(.a(s_81), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1118(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1119(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1120(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate785(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate786(.a(gate128inter0), .b(s_34), .O(gate128inter1));
  and2  gate787(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate788(.a(s_34), .O(gate128inter3));
  inv1  gate789(.a(s_35), .O(gate128inter4));
  nand2 gate790(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate791(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate792(.a(G408), .O(gate128inter7));
  inv1  gate793(.a(G409), .O(gate128inter8));
  nand2 gate794(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate795(.a(s_35), .b(gate128inter3), .O(gate128inter10));
  nor2  gate796(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate797(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate798(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate715(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate716(.a(gate133inter0), .b(s_24), .O(gate133inter1));
  and2  gate717(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate718(.a(s_24), .O(gate133inter3));
  inv1  gate719(.a(s_25), .O(gate133inter4));
  nand2 gate720(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate721(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate722(.a(G418), .O(gate133inter7));
  inv1  gate723(.a(G419), .O(gate133inter8));
  nand2 gate724(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate725(.a(s_25), .b(gate133inter3), .O(gate133inter10));
  nor2  gate726(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate727(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate728(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate995(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate996(.a(gate136inter0), .b(s_64), .O(gate136inter1));
  and2  gate997(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate998(.a(s_64), .O(gate136inter3));
  inv1  gate999(.a(s_65), .O(gate136inter4));
  nand2 gate1000(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1001(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1002(.a(G424), .O(gate136inter7));
  inv1  gate1003(.a(G425), .O(gate136inter8));
  nand2 gate1004(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1005(.a(s_65), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1006(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1007(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1008(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate589(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate590(.a(gate141inter0), .b(s_6), .O(gate141inter1));
  and2  gate591(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate592(.a(s_6), .O(gate141inter3));
  inv1  gate593(.a(s_7), .O(gate141inter4));
  nand2 gate594(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate595(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate596(.a(G450), .O(gate141inter7));
  inv1  gate597(.a(G453), .O(gate141inter8));
  nand2 gate598(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate599(.a(s_7), .b(gate141inter3), .O(gate141inter10));
  nor2  gate600(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate601(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate602(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate813(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate814(.a(gate155inter0), .b(s_38), .O(gate155inter1));
  and2  gate815(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate816(.a(s_38), .O(gate155inter3));
  inv1  gate817(.a(s_39), .O(gate155inter4));
  nand2 gate818(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate819(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate820(.a(G432), .O(gate155inter7));
  inv1  gate821(.a(G525), .O(gate155inter8));
  nand2 gate822(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate823(.a(s_39), .b(gate155inter3), .O(gate155inter10));
  nor2  gate824(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate825(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate826(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1247(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1248(.a(gate158inter0), .b(s_100), .O(gate158inter1));
  and2  gate1249(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1250(.a(s_100), .O(gate158inter3));
  inv1  gate1251(.a(s_101), .O(gate158inter4));
  nand2 gate1252(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1253(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1254(.a(G441), .O(gate158inter7));
  inv1  gate1255(.a(G528), .O(gate158inter8));
  nand2 gate1256(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1257(.a(s_101), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1258(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1259(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1260(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate743(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate744(.a(gate159inter0), .b(s_28), .O(gate159inter1));
  and2  gate745(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate746(.a(s_28), .O(gate159inter3));
  inv1  gate747(.a(s_29), .O(gate159inter4));
  nand2 gate748(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate749(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate750(.a(G444), .O(gate159inter7));
  inv1  gate751(.a(G531), .O(gate159inter8));
  nand2 gate752(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate753(.a(s_29), .b(gate159inter3), .O(gate159inter10));
  nor2  gate754(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate755(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate756(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1345(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1346(.a(gate167inter0), .b(s_114), .O(gate167inter1));
  and2  gate1347(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1348(.a(s_114), .O(gate167inter3));
  inv1  gate1349(.a(s_115), .O(gate167inter4));
  nand2 gate1350(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1351(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1352(.a(G468), .O(gate167inter7));
  inv1  gate1353(.a(G543), .O(gate167inter8));
  nand2 gate1354(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1355(.a(s_115), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1356(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1357(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1358(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1065(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1066(.a(gate174inter0), .b(s_74), .O(gate174inter1));
  and2  gate1067(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1068(.a(s_74), .O(gate174inter3));
  inv1  gate1069(.a(s_75), .O(gate174inter4));
  nand2 gate1070(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1071(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1072(.a(G489), .O(gate174inter7));
  inv1  gate1073(.a(G552), .O(gate174inter8));
  nand2 gate1074(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1075(.a(s_75), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1076(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1077(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1078(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1219(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1220(.a(gate177inter0), .b(s_96), .O(gate177inter1));
  and2  gate1221(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1222(.a(s_96), .O(gate177inter3));
  inv1  gate1223(.a(s_97), .O(gate177inter4));
  nand2 gate1224(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1225(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1226(.a(G498), .O(gate177inter7));
  inv1  gate1227(.a(G558), .O(gate177inter8));
  nand2 gate1228(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1229(.a(s_97), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1230(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1231(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1232(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate855(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate856(.a(gate195inter0), .b(s_44), .O(gate195inter1));
  and2  gate857(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate858(.a(s_44), .O(gate195inter3));
  inv1  gate859(.a(s_45), .O(gate195inter4));
  nand2 gate860(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate861(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate862(.a(G590), .O(gate195inter7));
  inv1  gate863(.a(G591), .O(gate195inter8));
  nand2 gate864(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate865(.a(s_45), .b(gate195inter3), .O(gate195inter10));
  nor2  gate866(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate867(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate868(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate659(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate660(.a(gate196inter0), .b(s_16), .O(gate196inter1));
  and2  gate661(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate662(.a(s_16), .O(gate196inter3));
  inv1  gate663(.a(s_17), .O(gate196inter4));
  nand2 gate664(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate665(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate666(.a(G592), .O(gate196inter7));
  inv1  gate667(.a(G593), .O(gate196inter8));
  nand2 gate668(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate669(.a(s_17), .b(gate196inter3), .O(gate196inter10));
  nor2  gate670(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate671(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate672(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate547(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate548(.a(gate198inter0), .b(s_0), .O(gate198inter1));
  and2  gate549(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate550(.a(s_0), .O(gate198inter3));
  inv1  gate551(.a(s_1), .O(gate198inter4));
  nand2 gate552(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate553(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate554(.a(G596), .O(gate198inter7));
  inv1  gate555(.a(G597), .O(gate198inter8));
  nand2 gate556(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate557(.a(s_1), .b(gate198inter3), .O(gate198inter10));
  nor2  gate558(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate559(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate560(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1037(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1038(.a(gate206inter0), .b(s_70), .O(gate206inter1));
  and2  gate1039(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1040(.a(s_70), .O(gate206inter3));
  inv1  gate1041(.a(s_71), .O(gate206inter4));
  nand2 gate1042(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1043(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1044(.a(G632), .O(gate206inter7));
  inv1  gate1045(.a(G637), .O(gate206inter8));
  nand2 gate1046(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1047(.a(s_71), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1048(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1049(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1050(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1205(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1206(.a(gate219inter0), .b(s_94), .O(gate219inter1));
  and2  gate1207(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1208(.a(s_94), .O(gate219inter3));
  inv1  gate1209(.a(s_95), .O(gate219inter4));
  nand2 gate1210(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1211(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1212(.a(G632), .O(gate219inter7));
  inv1  gate1213(.a(G681), .O(gate219inter8));
  nand2 gate1214(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1215(.a(s_95), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1216(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1217(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1218(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate799(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate800(.a(gate224inter0), .b(s_36), .O(gate224inter1));
  and2  gate801(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate802(.a(s_36), .O(gate224inter3));
  inv1  gate803(.a(s_37), .O(gate224inter4));
  nand2 gate804(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate805(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate806(.a(G637), .O(gate224inter7));
  inv1  gate807(.a(G687), .O(gate224inter8));
  nand2 gate808(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate809(.a(s_37), .b(gate224inter3), .O(gate224inter10));
  nor2  gate810(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate811(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate812(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate883(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate884(.a(gate225inter0), .b(s_48), .O(gate225inter1));
  and2  gate885(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate886(.a(s_48), .O(gate225inter3));
  inv1  gate887(.a(s_49), .O(gate225inter4));
  nand2 gate888(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate889(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate890(.a(G690), .O(gate225inter7));
  inv1  gate891(.a(G691), .O(gate225inter8));
  nand2 gate892(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate893(.a(s_49), .b(gate225inter3), .O(gate225inter10));
  nor2  gate894(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate895(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate896(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate925(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate926(.a(gate227inter0), .b(s_54), .O(gate227inter1));
  and2  gate927(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate928(.a(s_54), .O(gate227inter3));
  inv1  gate929(.a(s_55), .O(gate227inter4));
  nand2 gate930(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate931(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate932(.a(G694), .O(gate227inter7));
  inv1  gate933(.a(G695), .O(gate227inter8));
  nand2 gate934(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate935(.a(s_55), .b(gate227inter3), .O(gate227inter10));
  nor2  gate936(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate937(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate938(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1275(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1276(.a(gate228inter0), .b(s_104), .O(gate228inter1));
  and2  gate1277(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1278(.a(s_104), .O(gate228inter3));
  inv1  gate1279(.a(s_105), .O(gate228inter4));
  nand2 gate1280(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1281(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1282(.a(G696), .O(gate228inter7));
  inv1  gate1283(.a(G697), .O(gate228inter8));
  nand2 gate1284(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1285(.a(s_105), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1286(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1287(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1288(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1191(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1192(.a(gate240inter0), .b(s_92), .O(gate240inter1));
  and2  gate1193(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1194(.a(s_92), .O(gate240inter3));
  inv1  gate1195(.a(s_93), .O(gate240inter4));
  nand2 gate1196(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1197(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1198(.a(G263), .O(gate240inter7));
  inv1  gate1199(.a(G715), .O(gate240inter8));
  nand2 gate1200(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1201(.a(s_93), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1202(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1203(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1204(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1079(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1080(.a(gate248inter0), .b(s_76), .O(gate248inter1));
  and2  gate1081(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1082(.a(s_76), .O(gate248inter3));
  inv1  gate1083(.a(s_77), .O(gate248inter4));
  nand2 gate1084(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1085(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1086(.a(G727), .O(gate248inter7));
  inv1  gate1087(.a(G739), .O(gate248inter8));
  nand2 gate1088(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1089(.a(s_77), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1090(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1091(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1092(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1051(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1052(.a(gate256inter0), .b(s_72), .O(gate256inter1));
  and2  gate1053(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1054(.a(s_72), .O(gate256inter3));
  inv1  gate1055(.a(s_73), .O(gate256inter4));
  nand2 gate1056(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1057(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1058(.a(G715), .O(gate256inter7));
  inv1  gate1059(.a(G751), .O(gate256inter8));
  nand2 gate1060(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1061(.a(s_73), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1062(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1063(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1064(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1009(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1010(.a(gate263inter0), .b(s_66), .O(gate263inter1));
  and2  gate1011(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1012(.a(s_66), .O(gate263inter3));
  inv1  gate1013(.a(s_67), .O(gate263inter4));
  nand2 gate1014(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1015(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1016(.a(G766), .O(gate263inter7));
  inv1  gate1017(.a(G767), .O(gate263inter8));
  nand2 gate1018(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1019(.a(s_67), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1020(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1021(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1022(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate841(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate842(.a(gate264inter0), .b(s_42), .O(gate264inter1));
  and2  gate843(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate844(.a(s_42), .O(gate264inter3));
  inv1  gate845(.a(s_43), .O(gate264inter4));
  nand2 gate846(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate847(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate848(.a(G768), .O(gate264inter7));
  inv1  gate849(.a(G769), .O(gate264inter8));
  nand2 gate850(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate851(.a(s_43), .b(gate264inter3), .O(gate264inter10));
  nor2  gate852(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate853(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate854(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate911(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate912(.a(gate266inter0), .b(s_52), .O(gate266inter1));
  and2  gate913(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate914(.a(s_52), .O(gate266inter3));
  inv1  gate915(.a(s_53), .O(gate266inter4));
  nand2 gate916(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate917(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate918(.a(G645), .O(gate266inter7));
  inv1  gate919(.a(G773), .O(gate266inter8));
  nand2 gate920(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate921(.a(s_53), .b(gate266inter3), .O(gate266inter10));
  nor2  gate922(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate923(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate924(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate827(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate828(.a(gate270inter0), .b(s_40), .O(gate270inter1));
  and2  gate829(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate830(.a(s_40), .O(gate270inter3));
  inv1  gate831(.a(s_41), .O(gate270inter4));
  nand2 gate832(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate833(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate834(.a(G657), .O(gate270inter7));
  inv1  gate835(.a(G785), .O(gate270inter8));
  nand2 gate836(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate837(.a(s_41), .b(gate270inter3), .O(gate270inter10));
  nor2  gate838(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate839(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate840(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate729(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate730(.a(gate276inter0), .b(s_26), .O(gate276inter1));
  and2  gate731(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate732(.a(s_26), .O(gate276inter3));
  inv1  gate733(.a(s_27), .O(gate276inter4));
  nand2 gate734(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate735(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate736(.a(G773), .O(gate276inter7));
  inv1  gate737(.a(G797), .O(gate276inter8));
  nand2 gate738(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate739(.a(s_27), .b(gate276inter3), .O(gate276inter10));
  nor2  gate740(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate741(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate742(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate687(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate688(.a(gate290inter0), .b(s_20), .O(gate290inter1));
  and2  gate689(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate690(.a(s_20), .O(gate290inter3));
  inv1  gate691(.a(s_21), .O(gate290inter4));
  nand2 gate692(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate693(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate694(.a(G820), .O(gate290inter7));
  inv1  gate695(.a(G821), .O(gate290inter8));
  nand2 gate696(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate697(.a(s_21), .b(gate290inter3), .O(gate290inter10));
  nor2  gate698(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate699(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate700(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate561(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate562(.a(gate293inter0), .b(s_2), .O(gate293inter1));
  and2  gate563(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate564(.a(s_2), .O(gate293inter3));
  inv1  gate565(.a(s_3), .O(gate293inter4));
  nand2 gate566(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate567(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate568(.a(G828), .O(gate293inter7));
  inv1  gate569(.a(G829), .O(gate293inter8));
  nand2 gate570(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate571(.a(s_3), .b(gate293inter3), .O(gate293inter10));
  nor2  gate572(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate573(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate574(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate897(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate898(.a(gate295inter0), .b(s_50), .O(gate295inter1));
  and2  gate899(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate900(.a(s_50), .O(gate295inter3));
  inv1  gate901(.a(s_51), .O(gate295inter4));
  nand2 gate902(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate903(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate904(.a(G830), .O(gate295inter7));
  inv1  gate905(.a(G831), .O(gate295inter8));
  nand2 gate906(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate907(.a(s_51), .b(gate295inter3), .O(gate295inter10));
  nor2  gate908(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate909(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate910(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1177(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1178(.a(gate387inter0), .b(s_90), .O(gate387inter1));
  and2  gate1179(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1180(.a(s_90), .O(gate387inter3));
  inv1  gate1181(.a(s_91), .O(gate387inter4));
  nand2 gate1182(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1183(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1184(.a(G1), .O(gate387inter7));
  inv1  gate1185(.a(G1036), .O(gate387inter8));
  nand2 gate1186(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1187(.a(s_91), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1188(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1189(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1190(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate953(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate954(.a(gate397inter0), .b(s_58), .O(gate397inter1));
  and2  gate955(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate956(.a(s_58), .O(gate397inter3));
  inv1  gate957(.a(s_59), .O(gate397inter4));
  nand2 gate958(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate959(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate960(.a(G11), .O(gate397inter7));
  inv1  gate961(.a(G1066), .O(gate397inter8));
  nand2 gate962(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate963(.a(s_59), .b(gate397inter3), .O(gate397inter10));
  nor2  gate964(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate965(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate966(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1149(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1150(.a(gate408inter0), .b(s_86), .O(gate408inter1));
  and2  gate1151(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1152(.a(s_86), .O(gate408inter3));
  inv1  gate1153(.a(s_87), .O(gate408inter4));
  nand2 gate1154(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1155(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1156(.a(G22), .O(gate408inter7));
  inv1  gate1157(.a(G1099), .O(gate408inter8));
  nand2 gate1158(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1159(.a(s_87), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1160(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1161(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1162(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1373(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1374(.a(gate419inter0), .b(s_118), .O(gate419inter1));
  and2  gate1375(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1376(.a(s_118), .O(gate419inter3));
  inv1  gate1377(.a(s_119), .O(gate419inter4));
  nand2 gate1378(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1379(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1380(.a(G1), .O(gate419inter7));
  inv1  gate1381(.a(G1132), .O(gate419inter8));
  nand2 gate1382(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1383(.a(s_119), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1384(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1385(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1386(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1317(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1318(.a(gate421inter0), .b(s_110), .O(gate421inter1));
  and2  gate1319(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1320(.a(s_110), .O(gate421inter3));
  inv1  gate1321(.a(s_111), .O(gate421inter4));
  nand2 gate1322(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1323(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1324(.a(G2), .O(gate421inter7));
  inv1  gate1325(.a(G1135), .O(gate421inter8));
  nand2 gate1326(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1327(.a(s_111), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1328(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1329(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1330(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate631(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate632(.a(gate428inter0), .b(s_12), .O(gate428inter1));
  and2  gate633(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate634(.a(s_12), .O(gate428inter3));
  inv1  gate635(.a(s_13), .O(gate428inter4));
  nand2 gate636(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate637(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate638(.a(G1048), .O(gate428inter7));
  inv1  gate639(.a(G1144), .O(gate428inter8));
  nand2 gate640(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate641(.a(s_13), .b(gate428inter3), .O(gate428inter10));
  nor2  gate642(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate643(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate644(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate869(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate870(.a(gate430inter0), .b(s_46), .O(gate430inter1));
  and2  gate871(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate872(.a(s_46), .O(gate430inter3));
  inv1  gate873(.a(s_47), .O(gate430inter4));
  nand2 gate874(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate875(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate876(.a(G1051), .O(gate430inter7));
  inv1  gate877(.a(G1147), .O(gate430inter8));
  nand2 gate878(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate879(.a(s_47), .b(gate430inter3), .O(gate430inter10));
  nor2  gate880(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate881(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate882(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1289(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1290(.a(gate441inter0), .b(s_106), .O(gate441inter1));
  and2  gate1291(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1292(.a(s_106), .O(gate441inter3));
  inv1  gate1293(.a(s_107), .O(gate441inter4));
  nand2 gate1294(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1295(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1296(.a(G12), .O(gate441inter7));
  inv1  gate1297(.a(G1165), .O(gate441inter8));
  nand2 gate1298(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1299(.a(s_107), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1300(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1301(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1302(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate967(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate968(.a(gate445inter0), .b(s_60), .O(gate445inter1));
  and2  gate969(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate970(.a(s_60), .O(gate445inter3));
  inv1  gate971(.a(s_61), .O(gate445inter4));
  nand2 gate972(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate973(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate974(.a(G14), .O(gate445inter7));
  inv1  gate975(.a(G1171), .O(gate445inter8));
  nand2 gate976(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate977(.a(s_61), .b(gate445inter3), .O(gate445inter10));
  nor2  gate978(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate979(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate980(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate673(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate674(.a(gate446inter0), .b(s_18), .O(gate446inter1));
  and2  gate675(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate676(.a(s_18), .O(gate446inter3));
  inv1  gate677(.a(s_19), .O(gate446inter4));
  nand2 gate678(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate679(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate680(.a(G1075), .O(gate446inter7));
  inv1  gate681(.a(G1171), .O(gate446inter8));
  nand2 gate682(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate683(.a(s_19), .b(gate446inter3), .O(gate446inter10));
  nor2  gate684(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate685(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate686(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate701(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate702(.a(gate458inter0), .b(s_22), .O(gate458inter1));
  and2  gate703(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate704(.a(s_22), .O(gate458inter3));
  inv1  gate705(.a(s_23), .O(gate458inter4));
  nand2 gate706(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate707(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate708(.a(G1093), .O(gate458inter7));
  inv1  gate709(.a(G1189), .O(gate458inter8));
  nand2 gate710(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate711(.a(s_23), .b(gate458inter3), .O(gate458inter10));
  nor2  gate712(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate713(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate714(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate645(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate646(.a(gate459inter0), .b(s_14), .O(gate459inter1));
  and2  gate647(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate648(.a(s_14), .O(gate459inter3));
  inv1  gate649(.a(s_15), .O(gate459inter4));
  nand2 gate650(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate651(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate652(.a(G21), .O(gate459inter7));
  inv1  gate653(.a(G1192), .O(gate459inter8));
  nand2 gate654(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate655(.a(s_15), .b(gate459inter3), .O(gate459inter10));
  nor2  gate656(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate657(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate658(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate939(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate940(.a(gate465inter0), .b(s_56), .O(gate465inter1));
  and2  gate941(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate942(.a(s_56), .O(gate465inter3));
  inv1  gate943(.a(s_57), .O(gate465inter4));
  nand2 gate944(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate945(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate946(.a(G24), .O(gate465inter7));
  inv1  gate947(.a(G1201), .O(gate465inter8));
  nand2 gate948(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate949(.a(s_57), .b(gate465inter3), .O(gate465inter10));
  nor2  gate950(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate951(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate952(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate603(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate604(.a(gate471inter0), .b(s_8), .O(gate471inter1));
  and2  gate605(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate606(.a(s_8), .O(gate471inter3));
  inv1  gate607(.a(s_9), .O(gate471inter4));
  nand2 gate608(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate609(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate610(.a(G27), .O(gate471inter7));
  inv1  gate611(.a(G1210), .O(gate471inter8));
  nand2 gate612(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate613(.a(s_9), .b(gate471inter3), .O(gate471inter10));
  nor2  gate614(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate615(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate616(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate575(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate576(.a(gate483inter0), .b(s_4), .O(gate483inter1));
  and2  gate577(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate578(.a(s_4), .O(gate483inter3));
  inv1  gate579(.a(s_5), .O(gate483inter4));
  nand2 gate580(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate581(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate582(.a(G1228), .O(gate483inter7));
  inv1  gate583(.a(G1229), .O(gate483inter8));
  nand2 gate584(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate585(.a(s_5), .b(gate483inter3), .O(gate483inter10));
  nor2  gate586(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate587(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate588(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1023(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1024(.a(gate504inter0), .b(s_68), .O(gate504inter1));
  and2  gate1025(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1026(.a(s_68), .O(gate504inter3));
  inv1  gate1027(.a(s_69), .O(gate504inter4));
  nand2 gate1028(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1029(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1030(.a(G1270), .O(gate504inter7));
  inv1  gate1031(.a(G1271), .O(gate504inter8));
  nand2 gate1032(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1033(.a(s_69), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1034(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1035(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1036(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1121(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1122(.a(gate510inter0), .b(s_82), .O(gate510inter1));
  and2  gate1123(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1124(.a(s_82), .O(gate510inter3));
  inv1  gate1125(.a(s_83), .O(gate510inter4));
  nand2 gate1126(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1127(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1128(.a(G1282), .O(gate510inter7));
  inv1  gate1129(.a(G1283), .O(gate510inter8));
  nand2 gate1130(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1131(.a(s_83), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1132(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1133(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1134(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate981(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate982(.a(gate513inter0), .b(s_62), .O(gate513inter1));
  and2  gate983(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate984(.a(s_62), .O(gate513inter3));
  inv1  gate985(.a(s_63), .O(gate513inter4));
  nand2 gate986(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate987(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate988(.a(G1288), .O(gate513inter7));
  inv1  gate989(.a(G1289), .O(gate513inter8));
  nand2 gate990(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate991(.a(s_63), .b(gate513inter3), .O(gate513inter10));
  nor2  gate992(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate993(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate994(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule