module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1639(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1640(.a(gate11inter0), .b(s_156), .O(gate11inter1));
  and2  gate1641(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1642(.a(s_156), .O(gate11inter3));
  inv1  gate1643(.a(s_157), .O(gate11inter4));
  nand2 gate1644(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1645(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1646(.a(G5), .O(gate11inter7));
  inv1  gate1647(.a(G6), .O(gate11inter8));
  nand2 gate1648(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1649(.a(s_157), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1650(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1651(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1652(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate645(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate646(.a(gate12inter0), .b(s_14), .O(gate12inter1));
  and2  gate647(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate648(.a(s_14), .O(gate12inter3));
  inv1  gate649(.a(s_15), .O(gate12inter4));
  nand2 gate650(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate651(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate652(.a(G7), .O(gate12inter7));
  inv1  gate653(.a(G8), .O(gate12inter8));
  nand2 gate654(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate655(.a(s_15), .b(gate12inter3), .O(gate12inter10));
  nor2  gate656(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate657(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate658(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2171(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2172(.a(gate13inter0), .b(s_232), .O(gate13inter1));
  and2  gate2173(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2174(.a(s_232), .O(gate13inter3));
  inv1  gate2175(.a(s_233), .O(gate13inter4));
  nand2 gate2176(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2177(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2178(.a(G9), .O(gate13inter7));
  inv1  gate2179(.a(G10), .O(gate13inter8));
  nand2 gate2180(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2181(.a(s_233), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2182(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2183(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2184(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1499(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1500(.a(gate14inter0), .b(s_136), .O(gate14inter1));
  and2  gate1501(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1502(.a(s_136), .O(gate14inter3));
  inv1  gate1503(.a(s_137), .O(gate14inter4));
  nand2 gate1504(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1505(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1506(.a(G11), .O(gate14inter7));
  inv1  gate1507(.a(G12), .O(gate14inter8));
  nand2 gate1508(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1509(.a(s_137), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1510(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1511(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1512(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate2017(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2018(.a(gate15inter0), .b(s_210), .O(gate15inter1));
  and2  gate2019(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2020(.a(s_210), .O(gate15inter3));
  inv1  gate2021(.a(s_211), .O(gate15inter4));
  nand2 gate2022(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2023(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2024(.a(G13), .O(gate15inter7));
  inv1  gate2025(.a(G14), .O(gate15inter8));
  nand2 gate2026(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2027(.a(s_211), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2028(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2029(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2030(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate2269(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2270(.a(gate17inter0), .b(s_246), .O(gate17inter1));
  and2  gate2271(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2272(.a(s_246), .O(gate17inter3));
  inv1  gate2273(.a(s_247), .O(gate17inter4));
  nand2 gate2274(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2275(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2276(.a(G17), .O(gate17inter7));
  inv1  gate2277(.a(G18), .O(gate17inter8));
  nand2 gate2278(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2279(.a(s_247), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2280(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2281(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2282(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate925(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate926(.a(gate19inter0), .b(s_54), .O(gate19inter1));
  and2  gate927(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate928(.a(s_54), .O(gate19inter3));
  inv1  gate929(.a(s_55), .O(gate19inter4));
  nand2 gate930(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate931(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate932(.a(G21), .O(gate19inter7));
  inv1  gate933(.a(G22), .O(gate19inter8));
  nand2 gate934(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate935(.a(s_55), .b(gate19inter3), .O(gate19inter10));
  nor2  gate936(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate937(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate938(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1205(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1206(.a(gate20inter0), .b(s_94), .O(gate20inter1));
  and2  gate1207(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1208(.a(s_94), .O(gate20inter3));
  inv1  gate1209(.a(s_95), .O(gate20inter4));
  nand2 gate1210(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1211(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1212(.a(G23), .O(gate20inter7));
  inv1  gate1213(.a(G24), .O(gate20inter8));
  nand2 gate1214(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1215(.a(s_95), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1216(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1217(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1218(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1387(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1388(.a(gate24inter0), .b(s_120), .O(gate24inter1));
  and2  gate1389(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1390(.a(s_120), .O(gate24inter3));
  inv1  gate1391(.a(s_121), .O(gate24inter4));
  nand2 gate1392(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1393(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1394(.a(G31), .O(gate24inter7));
  inv1  gate1395(.a(G32), .O(gate24inter8));
  nand2 gate1396(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1397(.a(s_121), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1398(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1399(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1400(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate785(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate786(.a(gate26inter0), .b(s_34), .O(gate26inter1));
  and2  gate787(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate788(.a(s_34), .O(gate26inter3));
  inv1  gate789(.a(s_35), .O(gate26inter4));
  nand2 gate790(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate791(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate792(.a(G9), .O(gate26inter7));
  inv1  gate793(.a(G13), .O(gate26inter8));
  nand2 gate794(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate795(.a(s_35), .b(gate26inter3), .O(gate26inter10));
  nor2  gate796(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate797(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate798(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1765(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1766(.a(gate28inter0), .b(s_174), .O(gate28inter1));
  and2  gate1767(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1768(.a(s_174), .O(gate28inter3));
  inv1  gate1769(.a(s_175), .O(gate28inter4));
  nand2 gate1770(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1771(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1772(.a(G10), .O(gate28inter7));
  inv1  gate1773(.a(G14), .O(gate28inter8));
  nand2 gate1774(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1775(.a(s_175), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1776(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1777(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1778(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2773(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2774(.a(gate29inter0), .b(s_318), .O(gate29inter1));
  and2  gate2775(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2776(.a(s_318), .O(gate29inter3));
  inv1  gate2777(.a(s_319), .O(gate29inter4));
  nand2 gate2778(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2779(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2780(.a(G3), .O(gate29inter7));
  inv1  gate2781(.a(G7), .O(gate29inter8));
  nand2 gate2782(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2783(.a(s_319), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2784(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2785(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2786(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate883(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate884(.a(gate30inter0), .b(s_48), .O(gate30inter1));
  and2  gate885(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate886(.a(s_48), .O(gate30inter3));
  inv1  gate887(.a(s_49), .O(gate30inter4));
  nand2 gate888(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate889(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate890(.a(G11), .O(gate30inter7));
  inv1  gate891(.a(G15), .O(gate30inter8));
  nand2 gate892(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate893(.a(s_49), .b(gate30inter3), .O(gate30inter10));
  nor2  gate894(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate895(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate896(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1527(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1528(.a(gate36inter0), .b(s_140), .O(gate36inter1));
  and2  gate1529(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1530(.a(s_140), .O(gate36inter3));
  inv1  gate1531(.a(s_141), .O(gate36inter4));
  nand2 gate1532(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1533(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1534(.a(G26), .O(gate36inter7));
  inv1  gate1535(.a(G30), .O(gate36inter8));
  nand2 gate1536(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1537(.a(s_141), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1538(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1539(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1540(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1471(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1472(.a(gate37inter0), .b(s_132), .O(gate37inter1));
  and2  gate1473(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1474(.a(s_132), .O(gate37inter3));
  inv1  gate1475(.a(s_133), .O(gate37inter4));
  nand2 gate1476(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1477(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1478(.a(G19), .O(gate37inter7));
  inv1  gate1479(.a(G23), .O(gate37inter8));
  nand2 gate1480(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1481(.a(s_133), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1482(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1483(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1484(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2437(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2438(.a(gate38inter0), .b(s_270), .O(gate38inter1));
  and2  gate2439(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2440(.a(s_270), .O(gate38inter3));
  inv1  gate2441(.a(s_271), .O(gate38inter4));
  nand2 gate2442(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2443(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2444(.a(G27), .O(gate38inter7));
  inv1  gate2445(.a(G31), .O(gate38inter8));
  nand2 gate2446(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2447(.a(s_271), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2448(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2449(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2450(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1149(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1150(.a(gate40inter0), .b(s_86), .O(gate40inter1));
  and2  gate1151(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1152(.a(s_86), .O(gate40inter3));
  inv1  gate1153(.a(s_87), .O(gate40inter4));
  nand2 gate1154(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1155(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1156(.a(G28), .O(gate40inter7));
  inv1  gate1157(.a(G32), .O(gate40inter8));
  nand2 gate1158(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1159(.a(s_87), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1160(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1161(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1162(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate673(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate674(.a(gate43inter0), .b(s_18), .O(gate43inter1));
  and2  gate675(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate676(.a(s_18), .O(gate43inter3));
  inv1  gate677(.a(s_19), .O(gate43inter4));
  nand2 gate678(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate679(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate680(.a(G3), .O(gate43inter7));
  inv1  gate681(.a(G269), .O(gate43inter8));
  nand2 gate682(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate683(.a(s_19), .b(gate43inter3), .O(gate43inter10));
  nor2  gate684(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate685(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate686(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1891(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1892(.a(gate44inter0), .b(s_192), .O(gate44inter1));
  and2  gate1893(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1894(.a(s_192), .O(gate44inter3));
  inv1  gate1895(.a(s_193), .O(gate44inter4));
  nand2 gate1896(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1897(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1898(.a(G4), .O(gate44inter7));
  inv1  gate1899(.a(G269), .O(gate44inter8));
  nand2 gate1900(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1901(.a(s_193), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1902(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1903(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1904(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1849(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1850(.a(gate47inter0), .b(s_186), .O(gate47inter1));
  and2  gate1851(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1852(.a(s_186), .O(gate47inter3));
  inv1  gate1853(.a(s_187), .O(gate47inter4));
  nand2 gate1854(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1855(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1856(.a(G7), .O(gate47inter7));
  inv1  gate1857(.a(G275), .O(gate47inter8));
  nand2 gate1858(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1859(.a(s_187), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1860(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1861(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1862(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2591(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2592(.a(gate48inter0), .b(s_292), .O(gate48inter1));
  and2  gate2593(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2594(.a(s_292), .O(gate48inter3));
  inv1  gate2595(.a(s_293), .O(gate48inter4));
  nand2 gate2596(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2597(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2598(.a(G8), .O(gate48inter7));
  inv1  gate2599(.a(G275), .O(gate48inter8));
  nand2 gate2600(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2601(.a(s_293), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2602(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2603(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2604(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2493(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2494(.a(gate50inter0), .b(s_278), .O(gate50inter1));
  and2  gate2495(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2496(.a(s_278), .O(gate50inter3));
  inv1  gate2497(.a(s_279), .O(gate50inter4));
  nand2 gate2498(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2499(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2500(.a(G10), .O(gate50inter7));
  inv1  gate2501(.a(G278), .O(gate50inter8));
  nand2 gate2502(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2503(.a(s_279), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2504(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2505(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2506(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1541(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1542(.a(gate51inter0), .b(s_142), .O(gate51inter1));
  and2  gate1543(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1544(.a(s_142), .O(gate51inter3));
  inv1  gate1545(.a(s_143), .O(gate51inter4));
  nand2 gate1546(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1547(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1548(.a(G11), .O(gate51inter7));
  inv1  gate1549(.a(G281), .O(gate51inter8));
  nand2 gate1550(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1551(.a(s_143), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1552(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1553(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1554(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2297(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2298(.a(gate55inter0), .b(s_250), .O(gate55inter1));
  and2  gate2299(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2300(.a(s_250), .O(gate55inter3));
  inv1  gate2301(.a(s_251), .O(gate55inter4));
  nand2 gate2302(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2303(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2304(.a(G15), .O(gate55inter7));
  inv1  gate2305(.a(G287), .O(gate55inter8));
  nand2 gate2306(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2307(.a(s_251), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2308(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2309(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2310(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1961(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1962(.a(gate69inter0), .b(s_202), .O(gate69inter1));
  and2  gate1963(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1964(.a(s_202), .O(gate69inter3));
  inv1  gate1965(.a(s_203), .O(gate69inter4));
  nand2 gate1966(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1967(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1968(.a(G29), .O(gate69inter7));
  inv1  gate1969(.a(G308), .O(gate69inter8));
  nand2 gate1970(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1971(.a(s_203), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1972(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1973(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1974(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2633(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2634(.a(gate74inter0), .b(s_298), .O(gate74inter1));
  and2  gate2635(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2636(.a(s_298), .O(gate74inter3));
  inv1  gate2637(.a(s_299), .O(gate74inter4));
  nand2 gate2638(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2639(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2640(.a(G5), .O(gate74inter7));
  inv1  gate2641(.a(G314), .O(gate74inter8));
  nand2 gate2642(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2643(.a(s_299), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2644(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2645(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2646(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate2507(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2508(.a(gate75inter0), .b(s_280), .O(gate75inter1));
  and2  gate2509(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2510(.a(s_280), .O(gate75inter3));
  inv1  gate2511(.a(s_281), .O(gate75inter4));
  nand2 gate2512(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2513(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2514(.a(G9), .O(gate75inter7));
  inv1  gate2515(.a(G317), .O(gate75inter8));
  nand2 gate2516(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2517(.a(s_281), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2518(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2519(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2520(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2535(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2536(.a(gate79inter0), .b(s_284), .O(gate79inter1));
  and2  gate2537(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2538(.a(s_284), .O(gate79inter3));
  inv1  gate2539(.a(s_285), .O(gate79inter4));
  nand2 gate2540(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2541(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2542(.a(G10), .O(gate79inter7));
  inv1  gate2543(.a(G323), .O(gate79inter8));
  nand2 gate2544(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2545(.a(s_285), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2546(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2547(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2548(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1905(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1906(.a(gate81inter0), .b(s_194), .O(gate81inter1));
  and2  gate1907(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1908(.a(s_194), .O(gate81inter3));
  inv1  gate1909(.a(s_195), .O(gate81inter4));
  nand2 gate1910(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1911(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1912(.a(G3), .O(gate81inter7));
  inv1  gate1913(.a(G326), .O(gate81inter8));
  nand2 gate1914(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1915(.a(s_195), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1916(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1917(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1918(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate2101(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2102(.a(gate82inter0), .b(s_222), .O(gate82inter1));
  and2  gate2103(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2104(.a(s_222), .O(gate82inter3));
  inv1  gate2105(.a(s_223), .O(gate82inter4));
  nand2 gate2106(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2107(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2108(.a(G7), .O(gate82inter7));
  inv1  gate2109(.a(G326), .O(gate82inter8));
  nand2 gate2110(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2111(.a(s_223), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2112(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2113(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2114(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate911(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate912(.a(gate92inter0), .b(s_52), .O(gate92inter1));
  and2  gate913(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate914(.a(s_52), .O(gate92inter3));
  inv1  gate915(.a(s_53), .O(gate92inter4));
  nand2 gate916(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate917(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate918(.a(G29), .O(gate92inter7));
  inv1  gate919(.a(G341), .O(gate92inter8));
  nand2 gate920(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate921(.a(s_53), .b(gate92inter3), .O(gate92inter10));
  nor2  gate922(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate923(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate924(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2787(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2788(.a(gate96inter0), .b(s_320), .O(gate96inter1));
  and2  gate2789(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2790(.a(s_320), .O(gate96inter3));
  inv1  gate2791(.a(s_321), .O(gate96inter4));
  nand2 gate2792(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2793(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2794(.a(G30), .O(gate96inter7));
  inv1  gate2795(.a(G347), .O(gate96inter8));
  nand2 gate2796(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2797(.a(s_321), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2798(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2799(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2800(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2745(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2746(.a(gate97inter0), .b(s_314), .O(gate97inter1));
  and2  gate2747(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2748(.a(s_314), .O(gate97inter3));
  inv1  gate2749(.a(s_315), .O(gate97inter4));
  nand2 gate2750(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2751(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2752(.a(G19), .O(gate97inter7));
  inv1  gate2753(.a(G350), .O(gate97inter8));
  nand2 gate2754(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2755(.a(s_315), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2756(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2757(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2758(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2647(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2648(.a(gate102inter0), .b(s_300), .O(gate102inter1));
  and2  gate2649(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2650(.a(s_300), .O(gate102inter3));
  inv1  gate2651(.a(s_301), .O(gate102inter4));
  nand2 gate2652(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2653(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2654(.a(G24), .O(gate102inter7));
  inv1  gate2655(.a(G356), .O(gate102inter8));
  nand2 gate2656(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2657(.a(s_301), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2658(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2659(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2660(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2115(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2116(.a(gate106inter0), .b(s_224), .O(gate106inter1));
  and2  gate2117(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2118(.a(s_224), .O(gate106inter3));
  inv1  gate2119(.a(s_225), .O(gate106inter4));
  nand2 gate2120(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2121(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2122(.a(G364), .O(gate106inter7));
  inv1  gate2123(.a(G365), .O(gate106inter8));
  nand2 gate2124(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2125(.a(s_225), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2126(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2127(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2128(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2353(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2354(.a(gate107inter0), .b(s_258), .O(gate107inter1));
  and2  gate2355(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2356(.a(s_258), .O(gate107inter3));
  inv1  gate2357(.a(s_259), .O(gate107inter4));
  nand2 gate2358(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2359(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2360(.a(G366), .O(gate107inter7));
  inv1  gate2361(.a(G367), .O(gate107inter8));
  nand2 gate2362(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2363(.a(s_259), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2364(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2365(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2366(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1247(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1248(.a(gate108inter0), .b(s_100), .O(gate108inter1));
  and2  gate1249(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1250(.a(s_100), .O(gate108inter3));
  inv1  gate1251(.a(s_101), .O(gate108inter4));
  nand2 gate1252(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1253(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1254(.a(G368), .O(gate108inter7));
  inv1  gate1255(.a(G369), .O(gate108inter8));
  nand2 gate1256(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1257(.a(s_101), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1258(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1259(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1260(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1625(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1626(.a(gate110inter0), .b(s_154), .O(gate110inter1));
  and2  gate1627(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1628(.a(s_154), .O(gate110inter3));
  inv1  gate1629(.a(s_155), .O(gate110inter4));
  nand2 gate1630(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1631(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1632(.a(G372), .O(gate110inter7));
  inv1  gate1633(.a(G373), .O(gate110inter8));
  nand2 gate1634(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1635(.a(s_155), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1636(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1637(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1638(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate2409(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2410(.a(gate113inter0), .b(s_266), .O(gate113inter1));
  and2  gate2411(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2412(.a(s_266), .O(gate113inter3));
  inv1  gate2413(.a(s_267), .O(gate113inter4));
  nand2 gate2414(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2415(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2416(.a(G378), .O(gate113inter7));
  inv1  gate2417(.a(G379), .O(gate113inter8));
  nand2 gate2418(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2419(.a(s_267), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2420(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2421(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2422(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate1779(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1780(.a(gate114inter0), .b(s_176), .O(gate114inter1));
  and2  gate1781(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1782(.a(s_176), .O(gate114inter3));
  inv1  gate1783(.a(s_177), .O(gate114inter4));
  nand2 gate1784(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1785(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1786(.a(G380), .O(gate114inter7));
  inv1  gate1787(.a(G381), .O(gate114inter8));
  nand2 gate1788(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1789(.a(s_177), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1790(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1791(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1792(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1695(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1696(.a(gate115inter0), .b(s_164), .O(gate115inter1));
  and2  gate1697(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1698(.a(s_164), .O(gate115inter3));
  inv1  gate1699(.a(s_165), .O(gate115inter4));
  nand2 gate1700(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1701(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1702(.a(G382), .O(gate115inter7));
  inv1  gate1703(.a(G383), .O(gate115inter8));
  nand2 gate1704(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1705(.a(s_165), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1706(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1707(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1708(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1093(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1094(.a(gate118inter0), .b(s_78), .O(gate118inter1));
  and2  gate1095(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1096(.a(s_78), .O(gate118inter3));
  inv1  gate1097(.a(s_79), .O(gate118inter4));
  nand2 gate1098(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1099(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1100(.a(G388), .O(gate118inter7));
  inv1  gate1101(.a(G389), .O(gate118inter8));
  nand2 gate1102(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1103(.a(s_79), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1104(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1105(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1106(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate729(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate730(.a(gate121inter0), .b(s_26), .O(gate121inter1));
  and2  gate731(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate732(.a(s_26), .O(gate121inter3));
  inv1  gate733(.a(s_27), .O(gate121inter4));
  nand2 gate734(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate735(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate736(.a(G394), .O(gate121inter7));
  inv1  gate737(.a(G395), .O(gate121inter8));
  nand2 gate738(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate739(.a(s_27), .b(gate121inter3), .O(gate121inter10));
  nor2  gate740(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate741(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate742(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2157(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2158(.a(gate122inter0), .b(s_230), .O(gate122inter1));
  and2  gate2159(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2160(.a(s_230), .O(gate122inter3));
  inv1  gate2161(.a(s_231), .O(gate122inter4));
  nand2 gate2162(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2163(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2164(.a(G396), .O(gate122inter7));
  inv1  gate2165(.a(G397), .O(gate122inter8));
  nand2 gate2166(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2167(.a(s_231), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2168(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2169(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2170(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate2451(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2452(.a(gate123inter0), .b(s_272), .O(gate123inter1));
  and2  gate2453(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2454(.a(s_272), .O(gate123inter3));
  inv1  gate2455(.a(s_273), .O(gate123inter4));
  nand2 gate2456(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2457(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2458(.a(G398), .O(gate123inter7));
  inv1  gate2459(.a(G399), .O(gate123inter8));
  nand2 gate2460(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2461(.a(s_273), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2462(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2463(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2464(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate715(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate716(.a(gate125inter0), .b(s_24), .O(gate125inter1));
  and2  gate717(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate718(.a(s_24), .O(gate125inter3));
  inv1  gate719(.a(s_25), .O(gate125inter4));
  nand2 gate720(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate721(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate722(.a(G402), .O(gate125inter7));
  inv1  gate723(.a(G403), .O(gate125inter8));
  nand2 gate724(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate725(.a(s_25), .b(gate125inter3), .O(gate125inter10));
  nor2  gate726(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate727(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate728(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1751(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1752(.a(gate126inter0), .b(s_172), .O(gate126inter1));
  and2  gate1753(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1754(.a(s_172), .O(gate126inter3));
  inv1  gate1755(.a(s_173), .O(gate126inter4));
  nand2 gate1756(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1757(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1758(.a(G404), .O(gate126inter7));
  inv1  gate1759(.a(G405), .O(gate126inter8));
  nand2 gate1760(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1761(.a(s_173), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1762(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1763(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1764(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2255(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2256(.a(gate128inter0), .b(s_244), .O(gate128inter1));
  and2  gate2257(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2258(.a(s_244), .O(gate128inter3));
  inv1  gate2259(.a(s_245), .O(gate128inter4));
  nand2 gate2260(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2261(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2262(.a(G408), .O(gate128inter7));
  inv1  gate2263(.a(G409), .O(gate128inter8));
  nand2 gate2264(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2265(.a(s_245), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2266(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2267(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2268(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2661(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2662(.a(gate129inter0), .b(s_302), .O(gate129inter1));
  and2  gate2663(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2664(.a(s_302), .O(gate129inter3));
  inv1  gate2665(.a(s_303), .O(gate129inter4));
  nand2 gate2666(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2667(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2668(.a(G410), .O(gate129inter7));
  inv1  gate2669(.a(G411), .O(gate129inter8));
  nand2 gate2670(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2671(.a(s_303), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2672(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2673(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2674(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2563(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2564(.a(gate131inter0), .b(s_288), .O(gate131inter1));
  and2  gate2565(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2566(.a(s_288), .O(gate131inter3));
  inv1  gate2567(.a(s_289), .O(gate131inter4));
  nand2 gate2568(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2569(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2570(.a(G414), .O(gate131inter7));
  inv1  gate2571(.a(G415), .O(gate131inter8));
  nand2 gate2572(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2573(.a(s_289), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2574(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2575(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2576(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1457(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1458(.a(gate133inter0), .b(s_130), .O(gate133inter1));
  and2  gate1459(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1460(.a(s_130), .O(gate133inter3));
  inv1  gate1461(.a(s_131), .O(gate133inter4));
  nand2 gate1462(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1463(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1464(.a(G418), .O(gate133inter7));
  inv1  gate1465(.a(G419), .O(gate133inter8));
  nand2 gate1466(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1467(.a(s_131), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1468(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1469(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1470(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2339(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2340(.a(gate137inter0), .b(s_256), .O(gate137inter1));
  and2  gate2341(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2342(.a(s_256), .O(gate137inter3));
  inv1  gate2343(.a(s_257), .O(gate137inter4));
  nand2 gate2344(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2345(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2346(.a(G426), .O(gate137inter7));
  inv1  gate2347(.a(G429), .O(gate137inter8));
  nand2 gate2348(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2349(.a(s_257), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2350(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2351(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2352(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1065(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1066(.a(gate140inter0), .b(s_74), .O(gate140inter1));
  and2  gate1067(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1068(.a(s_74), .O(gate140inter3));
  inv1  gate1069(.a(s_75), .O(gate140inter4));
  nand2 gate1070(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1071(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1072(.a(G444), .O(gate140inter7));
  inv1  gate1073(.a(G447), .O(gate140inter8));
  nand2 gate1074(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1075(.a(s_75), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1076(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1077(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1078(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2381(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2382(.a(gate142inter0), .b(s_262), .O(gate142inter1));
  and2  gate2383(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2384(.a(s_262), .O(gate142inter3));
  inv1  gate2385(.a(s_263), .O(gate142inter4));
  nand2 gate2386(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2387(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2388(.a(G456), .O(gate142inter7));
  inv1  gate2389(.a(G459), .O(gate142inter8));
  nand2 gate2390(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2391(.a(s_263), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2392(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2393(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2394(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate855(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate856(.a(gate144inter0), .b(s_44), .O(gate144inter1));
  and2  gate857(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate858(.a(s_44), .O(gate144inter3));
  inv1  gate859(.a(s_45), .O(gate144inter4));
  nand2 gate860(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate861(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate862(.a(G468), .O(gate144inter7));
  inv1  gate863(.a(G471), .O(gate144inter8));
  nand2 gate864(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate865(.a(s_45), .b(gate144inter3), .O(gate144inter10));
  nor2  gate866(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate867(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate868(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2087(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2088(.a(gate145inter0), .b(s_220), .O(gate145inter1));
  and2  gate2089(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2090(.a(s_220), .O(gate145inter3));
  inv1  gate2091(.a(s_221), .O(gate145inter4));
  nand2 gate2092(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2093(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2094(.a(G474), .O(gate145inter7));
  inv1  gate2095(.a(G477), .O(gate145inter8));
  nand2 gate2096(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2097(.a(s_221), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2098(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2099(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2100(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate743(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate744(.a(gate146inter0), .b(s_28), .O(gate146inter1));
  and2  gate745(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate746(.a(s_28), .O(gate146inter3));
  inv1  gate747(.a(s_29), .O(gate146inter4));
  nand2 gate748(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate749(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate750(.a(G480), .O(gate146inter7));
  inv1  gate751(.a(G483), .O(gate146inter8));
  nand2 gate752(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate753(.a(s_29), .b(gate146inter3), .O(gate146inter10));
  nor2  gate754(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate755(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate756(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1737(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1738(.a(gate147inter0), .b(s_170), .O(gate147inter1));
  and2  gate1739(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1740(.a(s_170), .O(gate147inter3));
  inv1  gate1741(.a(s_171), .O(gate147inter4));
  nand2 gate1742(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1743(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1744(.a(G486), .O(gate147inter7));
  inv1  gate1745(.a(G489), .O(gate147inter8));
  nand2 gate1746(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1747(.a(s_171), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1748(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1749(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1750(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1331(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1332(.a(gate150inter0), .b(s_112), .O(gate150inter1));
  and2  gate1333(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1334(.a(s_112), .O(gate150inter3));
  inv1  gate1335(.a(s_113), .O(gate150inter4));
  nand2 gate1336(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1337(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1338(.a(G504), .O(gate150inter7));
  inv1  gate1339(.a(G507), .O(gate150inter8));
  nand2 gate1340(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1341(.a(s_113), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1342(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1343(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1344(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1303(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1304(.a(gate154inter0), .b(s_108), .O(gate154inter1));
  and2  gate1305(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1306(.a(s_108), .O(gate154inter3));
  inv1  gate1307(.a(s_109), .O(gate154inter4));
  nand2 gate1308(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1309(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1310(.a(G429), .O(gate154inter7));
  inv1  gate1311(.a(G522), .O(gate154inter8));
  nand2 gate1312(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1313(.a(s_109), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1314(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1315(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1316(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate827(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate828(.a(gate155inter0), .b(s_40), .O(gate155inter1));
  and2  gate829(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate830(.a(s_40), .O(gate155inter3));
  inv1  gate831(.a(s_41), .O(gate155inter4));
  nand2 gate832(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate833(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate834(.a(G432), .O(gate155inter7));
  inv1  gate835(.a(G525), .O(gate155inter8));
  nand2 gate836(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate837(.a(s_41), .b(gate155inter3), .O(gate155inter10));
  nor2  gate838(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate839(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate840(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2045(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2046(.a(gate156inter0), .b(s_214), .O(gate156inter1));
  and2  gate2047(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2048(.a(s_214), .O(gate156inter3));
  inv1  gate2049(.a(s_215), .O(gate156inter4));
  nand2 gate2050(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2051(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2052(.a(G435), .O(gate156inter7));
  inv1  gate2053(.a(G525), .O(gate156inter8));
  nand2 gate2054(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2055(.a(s_215), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2056(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2057(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2058(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2423(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2424(.a(gate157inter0), .b(s_268), .O(gate157inter1));
  and2  gate2425(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2426(.a(s_268), .O(gate157inter3));
  inv1  gate2427(.a(s_269), .O(gate157inter4));
  nand2 gate2428(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2429(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2430(.a(G438), .O(gate157inter7));
  inv1  gate2431(.a(G528), .O(gate157inter8));
  nand2 gate2432(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2433(.a(s_269), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2434(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2435(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2436(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate841(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate842(.a(gate158inter0), .b(s_42), .O(gate158inter1));
  and2  gate843(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate844(.a(s_42), .O(gate158inter3));
  inv1  gate845(.a(s_43), .O(gate158inter4));
  nand2 gate846(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate847(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate848(.a(G441), .O(gate158inter7));
  inv1  gate849(.a(G528), .O(gate158inter8));
  nand2 gate850(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate851(.a(s_43), .b(gate158inter3), .O(gate158inter10));
  nor2  gate852(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate853(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate854(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2311(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2312(.a(gate159inter0), .b(s_252), .O(gate159inter1));
  and2  gate2313(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2314(.a(s_252), .O(gate159inter3));
  inv1  gate2315(.a(s_253), .O(gate159inter4));
  nand2 gate2316(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2317(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2318(.a(G444), .O(gate159inter7));
  inv1  gate2319(.a(G531), .O(gate159inter8));
  nand2 gate2320(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2321(.a(s_253), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2322(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2323(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2324(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2815(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2816(.a(gate160inter0), .b(s_324), .O(gate160inter1));
  and2  gate2817(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2818(.a(s_324), .O(gate160inter3));
  inv1  gate2819(.a(s_325), .O(gate160inter4));
  nand2 gate2820(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2821(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2822(.a(G447), .O(gate160inter7));
  inv1  gate2823(.a(G531), .O(gate160inter8));
  nand2 gate2824(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2825(.a(s_325), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2826(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2827(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2828(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1611(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1612(.a(gate162inter0), .b(s_152), .O(gate162inter1));
  and2  gate1613(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1614(.a(s_152), .O(gate162inter3));
  inv1  gate1615(.a(s_153), .O(gate162inter4));
  nand2 gate1616(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1617(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1618(.a(G453), .O(gate162inter7));
  inv1  gate1619(.a(G534), .O(gate162inter8));
  nand2 gate1620(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1621(.a(s_153), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1622(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1623(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1624(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2521(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2522(.a(gate165inter0), .b(s_282), .O(gate165inter1));
  and2  gate2523(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2524(.a(s_282), .O(gate165inter3));
  inv1  gate2525(.a(s_283), .O(gate165inter4));
  nand2 gate2526(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2527(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2528(.a(G462), .O(gate165inter7));
  inv1  gate2529(.a(G540), .O(gate165inter8));
  nand2 gate2530(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2531(.a(s_283), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2532(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2533(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2534(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2395(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2396(.a(gate168inter0), .b(s_264), .O(gate168inter1));
  and2  gate2397(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2398(.a(s_264), .O(gate168inter3));
  inv1  gate2399(.a(s_265), .O(gate168inter4));
  nand2 gate2400(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2401(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2402(.a(G471), .O(gate168inter7));
  inv1  gate2403(.a(G543), .O(gate168inter8));
  nand2 gate2404(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2405(.a(s_265), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2406(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2407(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2408(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2283(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2284(.a(gate169inter0), .b(s_248), .O(gate169inter1));
  and2  gate2285(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2286(.a(s_248), .O(gate169inter3));
  inv1  gate2287(.a(s_249), .O(gate169inter4));
  nand2 gate2288(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2289(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2290(.a(G474), .O(gate169inter7));
  inv1  gate2291(.a(G546), .O(gate169inter8));
  nand2 gate2292(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2293(.a(s_249), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2294(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2295(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2296(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1415(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1416(.a(gate171inter0), .b(s_124), .O(gate171inter1));
  and2  gate1417(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1418(.a(s_124), .O(gate171inter3));
  inv1  gate1419(.a(s_125), .O(gate171inter4));
  nand2 gate1420(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1421(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1422(.a(G480), .O(gate171inter7));
  inv1  gate1423(.a(G549), .O(gate171inter8));
  nand2 gate1424(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1425(.a(s_125), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1426(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1427(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1428(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2605(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2606(.a(gate173inter0), .b(s_294), .O(gate173inter1));
  and2  gate2607(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2608(.a(s_294), .O(gate173inter3));
  inv1  gate2609(.a(s_295), .O(gate173inter4));
  nand2 gate2610(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2611(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2612(.a(G486), .O(gate173inter7));
  inv1  gate2613(.a(G552), .O(gate173inter8));
  nand2 gate2614(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2615(.a(s_295), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2616(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2617(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2618(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate799(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate800(.a(gate174inter0), .b(s_36), .O(gate174inter1));
  and2  gate801(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate802(.a(s_36), .O(gate174inter3));
  inv1  gate803(.a(s_37), .O(gate174inter4));
  nand2 gate804(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate805(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate806(.a(G489), .O(gate174inter7));
  inv1  gate807(.a(G552), .O(gate174inter8));
  nand2 gate808(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate809(.a(s_37), .b(gate174inter3), .O(gate174inter10));
  nor2  gate810(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate811(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate812(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate757(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate758(.a(gate177inter0), .b(s_30), .O(gate177inter1));
  and2  gate759(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate760(.a(s_30), .O(gate177inter3));
  inv1  gate761(.a(s_31), .O(gate177inter4));
  nand2 gate762(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate763(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate764(.a(G498), .O(gate177inter7));
  inv1  gate765(.a(G558), .O(gate177inter8));
  nand2 gate766(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate767(.a(s_31), .b(gate177inter3), .O(gate177inter10));
  nor2  gate768(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate769(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate770(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1401(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1402(.a(gate179inter0), .b(s_122), .O(gate179inter1));
  and2  gate1403(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1404(.a(s_122), .O(gate179inter3));
  inv1  gate1405(.a(s_123), .O(gate179inter4));
  nand2 gate1406(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1407(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1408(.a(G504), .O(gate179inter7));
  inv1  gate1409(.a(G561), .O(gate179inter8));
  nand2 gate1410(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1411(.a(s_123), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1412(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1413(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1414(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1835(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1836(.a(gate180inter0), .b(s_184), .O(gate180inter1));
  and2  gate1837(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1838(.a(s_184), .O(gate180inter3));
  inv1  gate1839(.a(s_185), .O(gate180inter4));
  nand2 gate1840(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1841(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1842(.a(G507), .O(gate180inter7));
  inv1  gate1843(.a(G561), .O(gate180inter8));
  nand2 gate1844(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1845(.a(s_185), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1846(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1847(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1848(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1933(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1934(.a(gate183inter0), .b(s_198), .O(gate183inter1));
  and2  gate1935(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1936(.a(s_198), .O(gate183inter3));
  inv1  gate1937(.a(s_199), .O(gate183inter4));
  nand2 gate1938(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1939(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1940(.a(G516), .O(gate183inter7));
  inv1  gate1941(.a(G567), .O(gate183inter8));
  nand2 gate1942(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1943(.a(s_199), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1944(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1945(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1946(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2549(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2550(.a(gate185inter0), .b(s_286), .O(gate185inter1));
  and2  gate2551(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2552(.a(s_286), .O(gate185inter3));
  inv1  gate2553(.a(s_287), .O(gate185inter4));
  nand2 gate2554(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2555(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2556(.a(G570), .O(gate185inter7));
  inv1  gate2557(.a(G571), .O(gate185inter8));
  nand2 gate2558(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2559(.a(s_287), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2560(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2561(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2562(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate575(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate576(.a(gate186inter0), .b(s_4), .O(gate186inter1));
  and2  gate577(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate578(.a(s_4), .O(gate186inter3));
  inv1  gate579(.a(s_5), .O(gate186inter4));
  nand2 gate580(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate581(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate582(.a(G572), .O(gate186inter7));
  inv1  gate583(.a(G573), .O(gate186inter8));
  nand2 gate584(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate585(.a(s_5), .b(gate186inter3), .O(gate186inter10));
  nor2  gate586(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate587(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate588(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2801(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2802(.a(gate188inter0), .b(s_322), .O(gate188inter1));
  and2  gate2803(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2804(.a(s_322), .O(gate188inter3));
  inv1  gate2805(.a(s_323), .O(gate188inter4));
  nand2 gate2806(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2807(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2808(.a(G576), .O(gate188inter7));
  inv1  gate2809(.a(G577), .O(gate188inter8));
  nand2 gate2810(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2811(.a(s_323), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2812(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2813(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2814(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate953(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate954(.a(gate189inter0), .b(s_58), .O(gate189inter1));
  and2  gate955(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate956(.a(s_58), .O(gate189inter3));
  inv1  gate957(.a(s_59), .O(gate189inter4));
  nand2 gate958(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate959(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate960(.a(G578), .O(gate189inter7));
  inv1  gate961(.a(G579), .O(gate189inter8));
  nand2 gate962(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate963(.a(s_59), .b(gate189inter3), .O(gate189inter10));
  nor2  gate964(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate965(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate966(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2227(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2228(.a(gate193inter0), .b(s_240), .O(gate193inter1));
  and2  gate2229(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2230(.a(s_240), .O(gate193inter3));
  inv1  gate2231(.a(s_241), .O(gate193inter4));
  nand2 gate2232(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2233(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2234(.a(G586), .O(gate193inter7));
  inv1  gate2235(.a(G587), .O(gate193inter8));
  nand2 gate2236(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2237(.a(s_241), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2238(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2239(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2240(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2843(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2844(.a(gate195inter0), .b(s_328), .O(gate195inter1));
  and2  gate2845(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2846(.a(s_328), .O(gate195inter3));
  inv1  gate2847(.a(s_329), .O(gate195inter4));
  nand2 gate2848(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2849(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2850(.a(G590), .O(gate195inter7));
  inv1  gate2851(.a(G591), .O(gate195inter8));
  nand2 gate2852(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2853(.a(s_329), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2854(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2855(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2856(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1009(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1010(.a(gate202inter0), .b(s_66), .O(gate202inter1));
  and2  gate1011(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1012(.a(s_66), .O(gate202inter3));
  inv1  gate1013(.a(s_67), .O(gate202inter4));
  nand2 gate1014(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1015(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1016(.a(G612), .O(gate202inter7));
  inv1  gate1017(.a(G617), .O(gate202inter8));
  nand2 gate1018(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1019(.a(s_67), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1020(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1021(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1022(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate995(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate996(.a(gate203inter0), .b(s_64), .O(gate203inter1));
  and2  gate997(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate998(.a(s_64), .O(gate203inter3));
  inv1  gate999(.a(s_65), .O(gate203inter4));
  nand2 gate1000(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1001(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1002(.a(G602), .O(gate203inter7));
  inv1  gate1003(.a(G612), .O(gate203inter8));
  nand2 gate1004(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1005(.a(s_65), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1006(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1007(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1008(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1989(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1990(.a(gate205inter0), .b(s_206), .O(gate205inter1));
  and2  gate1991(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1992(.a(s_206), .O(gate205inter3));
  inv1  gate1993(.a(s_207), .O(gate205inter4));
  nand2 gate1994(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1995(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1996(.a(G622), .O(gate205inter7));
  inv1  gate1997(.a(G627), .O(gate205inter8));
  nand2 gate1998(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1999(.a(s_207), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2000(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2001(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2002(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2829(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2830(.a(gate211inter0), .b(s_326), .O(gate211inter1));
  and2  gate2831(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2832(.a(s_326), .O(gate211inter3));
  inv1  gate2833(.a(s_327), .O(gate211inter4));
  nand2 gate2834(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2835(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2836(.a(G612), .O(gate211inter7));
  inv1  gate2837(.a(G669), .O(gate211inter8));
  nand2 gate2838(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2839(.a(s_327), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2840(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2841(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2842(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2577(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2578(.a(gate212inter0), .b(s_290), .O(gate212inter1));
  and2  gate2579(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2580(.a(s_290), .O(gate212inter3));
  inv1  gate2581(.a(s_291), .O(gate212inter4));
  nand2 gate2582(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2583(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2584(.a(G617), .O(gate212inter7));
  inv1  gate2585(.a(G669), .O(gate212inter8));
  nand2 gate2586(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2587(.a(s_291), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2588(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2589(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2590(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1443(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1444(.a(gate216inter0), .b(s_128), .O(gate216inter1));
  and2  gate1445(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1446(.a(s_128), .O(gate216inter3));
  inv1  gate1447(.a(s_129), .O(gate216inter4));
  nand2 gate1448(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1449(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1450(.a(G617), .O(gate216inter7));
  inv1  gate1451(.a(G675), .O(gate216inter8));
  nand2 gate1452(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1453(.a(s_129), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1454(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1455(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1456(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate617(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate618(.a(gate225inter0), .b(s_10), .O(gate225inter1));
  and2  gate619(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate620(.a(s_10), .O(gate225inter3));
  inv1  gate621(.a(s_11), .O(gate225inter4));
  nand2 gate622(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate623(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate624(.a(G690), .O(gate225inter7));
  inv1  gate625(.a(G691), .O(gate225inter8));
  nand2 gate626(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate627(.a(s_11), .b(gate225inter3), .O(gate225inter10));
  nor2  gate628(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate629(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate630(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1317(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1318(.a(gate226inter0), .b(s_110), .O(gate226inter1));
  and2  gate1319(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1320(.a(s_110), .O(gate226inter3));
  inv1  gate1321(.a(s_111), .O(gate226inter4));
  nand2 gate1322(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1323(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1324(.a(G692), .O(gate226inter7));
  inv1  gate1325(.a(G693), .O(gate226inter8));
  nand2 gate1326(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1327(.a(s_111), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1328(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1329(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1330(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2325(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2326(.a(gate229inter0), .b(s_254), .O(gate229inter1));
  and2  gate2327(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2328(.a(s_254), .O(gate229inter3));
  inv1  gate2329(.a(s_255), .O(gate229inter4));
  nand2 gate2330(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2331(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2332(.a(G698), .O(gate229inter7));
  inv1  gate2333(.a(G699), .O(gate229inter8));
  nand2 gate2334(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2335(.a(s_255), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2336(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2337(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2338(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate939(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate940(.a(gate232inter0), .b(s_56), .O(gate232inter1));
  and2  gate941(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate942(.a(s_56), .O(gate232inter3));
  inv1  gate943(.a(s_57), .O(gate232inter4));
  nand2 gate944(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate945(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate946(.a(G704), .O(gate232inter7));
  inv1  gate947(.a(G705), .O(gate232inter8));
  nand2 gate948(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate949(.a(s_57), .b(gate232inter3), .O(gate232inter10));
  nor2  gate950(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate951(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate952(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2717(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2718(.a(gate237inter0), .b(s_310), .O(gate237inter1));
  and2  gate2719(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2720(.a(s_310), .O(gate237inter3));
  inv1  gate2721(.a(s_311), .O(gate237inter4));
  nand2 gate2722(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2723(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2724(.a(G254), .O(gate237inter7));
  inv1  gate2725(.a(G706), .O(gate237inter8));
  nand2 gate2726(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2727(.a(s_311), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2728(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2729(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2730(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate897(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate898(.a(gate238inter0), .b(s_50), .O(gate238inter1));
  and2  gate899(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate900(.a(s_50), .O(gate238inter3));
  inv1  gate901(.a(s_51), .O(gate238inter4));
  nand2 gate902(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate903(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate904(.a(G257), .O(gate238inter7));
  inv1  gate905(.a(G709), .O(gate238inter8));
  nand2 gate906(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate907(.a(s_51), .b(gate238inter3), .O(gate238inter10));
  nor2  gate908(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate909(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate910(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1947(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1948(.a(gate240inter0), .b(s_200), .O(gate240inter1));
  and2  gate1949(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1950(.a(s_200), .O(gate240inter3));
  inv1  gate1951(.a(s_201), .O(gate240inter4));
  nand2 gate1952(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1953(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1954(.a(G263), .O(gate240inter7));
  inv1  gate1955(.a(G715), .O(gate240inter8));
  nand2 gate1956(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1957(.a(s_201), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1958(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1959(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1960(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1555(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1556(.a(gate241inter0), .b(s_144), .O(gate241inter1));
  and2  gate1557(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1558(.a(s_144), .O(gate241inter3));
  inv1  gate1559(.a(s_145), .O(gate241inter4));
  nand2 gate1560(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1561(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1562(.a(G242), .O(gate241inter7));
  inv1  gate1563(.a(G730), .O(gate241inter8));
  nand2 gate1564(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1565(.a(s_145), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1566(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1567(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1568(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1135(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1136(.a(gate242inter0), .b(s_84), .O(gate242inter1));
  and2  gate1137(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1138(.a(s_84), .O(gate242inter3));
  inv1  gate1139(.a(s_85), .O(gate242inter4));
  nand2 gate1140(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1141(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1142(.a(G718), .O(gate242inter7));
  inv1  gate1143(.a(G730), .O(gate242inter8));
  nand2 gate1144(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1145(.a(s_85), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1146(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1147(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1148(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1429(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1430(.a(gate246inter0), .b(s_126), .O(gate246inter1));
  and2  gate1431(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1432(.a(s_126), .O(gate246inter3));
  inv1  gate1433(.a(s_127), .O(gate246inter4));
  nand2 gate1434(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1435(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1436(.a(G724), .O(gate246inter7));
  inv1  gate1437(.a(G736), .O(gate246inter8));
  nand2 gate1438(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1439(.a(s_127), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1440(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1441(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1442(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1485(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1486(.a(gate247inter0), .b(s_134), .O(gate247inter1));
  and2  gate1487(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1488(.a(s_134), .O(gate247inter3));
  inv1  gate1489(.a(s_135), .O(gate247inter4));
  nand2 gate1490(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1491(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1492(.a(G251), .O(gate247inter7));
  inv1  gate1493(.a(G739), .O(gate247inter8));
  nand2 gate1494(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1495(.a(s_135), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1496(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1497(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1498(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2479(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2480(.a(gate249inter0), .b(s_276), .O(gate249inter1));
  and2  gate2481(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2482(.a(s_276), .O(gate249inter3));
  inv1  gate2483(.a(s_277), .O(gate249inter4));
  nand2 gate2484(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2485(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2486(.a(G254), .O(gate249inter7));
  inv1  gate2487(.a(G742), .O(gate249inter8));
  nand2 gate2488(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2489(.a(s_277), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2490(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2491(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2492(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1877(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1878(.a(gate255inter0), .b(s_190), .O(gate255inter1));
  and2  gate1879(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1880(.a(s_190), .O(gate255inter3));
  inv1  gate1881(.a(s_191), .O(gate255inter4));
  nand2 gate1882(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1883(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1884(.a(G263), .O(gate255inter7));
  inv1  gate1885(.a(G751), .O(gate255inter8));
  nand2 gate1886(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1887(.a(s_191), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1888(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1889(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1890(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate2073(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2074(.a(gate256inter0), .b(s_218), .O(gate256inter1));
  and2  gate2075(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2076(.a(s_218), .O(gate256inter3));
  inv1  gate2077(.a(s_219), .O(gate256inter4));
  nand2 gate2078(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2079(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2080(.a(G715), .O(gate256inter7));
  inv1  gate2081(.a(G751), .O(gate256inter8));
  nand2 gate2082(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2083(.a(s_219), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2084(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2085(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2086(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1653(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1654(.a(gate261inter0), .b(s_158), .O(gate261inter1));
  and2  gate1655(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1656(.a(s_158), .O(gate261inter3));
  inv1  gate1657(.a(s_159), .O(gate261inter4));
  nand2 gate1658(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1659(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1660(.a(G762), .O(gate261inter7));
  inv1  gate1661(.a(G763), .O(gate261inter8));
  nand2 gate1662(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1663(.a(s_159), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1664(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1665(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1666(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate967(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate968(.a(gate263inter0), .b(s_60), .O(gate263inter1));
  and2  gate969(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate970(.a(s_60), .O(gate263inter3));
  inv1  gate971(.a(s_61), .O(gate263inter4));
  nand2 gate972(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate973(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate974(.a(G766), .O(gate263inter7));
  inv1  gate975(.a(G767), .O(gate263inter8));
  nand2 gate976(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate977(.a(s_61), .b(gate263inter3), .O(gate263inter10));
  nor2  gate978(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate979(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate980(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2857(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2858(.a(gate264inter0), .b(s_330), .O(gate264inter1));
  and2  gate2859(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2860(.a(s_330), .O(gate264inter3));
  inv1  gate2861(.a(s_331), .O(gate264inter4));
  nand2 gate2862(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2863(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2864(.a(G768), .O(gate264inter7));
  inv1  gate2865(.a(G769), .O(gate264inter8));
  nand2 gate2866(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2867(.a(s_331), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2868(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2869(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2870(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2213(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2214(.a(gate268inter0), .b(s_238), .O(gate268inter1));
  and2  gate2215(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2216(.a(s_238), .O(gate268inter3));
  inv1  gate2217(.a(s_239), .O(gate268inter4));
  nand2 gate2218(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2219(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2220(.a(G651), .O(gate268inter7));
  inv1  gate2221(.a(G779), .O(gate268inter8));
  nand2 gate2222(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2223(.a(s_239), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2224(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2225(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2226(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate701(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate702(.a(gate270inter0), .b(s_22), .O(gate270inter1));
  and2  gate703(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate704(.a(s_22), .O(gate270inter3));
  inv1  gate705(.a(s_23), .O(gate270inter4));
  nand2 gate706(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate707(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate708(.a(G657), .O(gate270inter7));
  inv1  gate709(.a(G785), .O(gate270inter8));
  nand2 gate710(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate711(.a(s_23), .b(gate270inter3), .O(gate270inter10));
  nor2  gate712(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate713(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate714(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1569(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1570(.a(gate271inter0), .b(s_146), .O(gate271inter1));
  and2  gate1571(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1572(.a(s_146), .O(gate271inter3));
  inv1  gate1573(.a(s_147), .O(gate271inter4));
  nand2 gate1574(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1575(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1576(.a(G660), .O(gate271inter7));
  inv1  gate1577(.a(G788), .O(gate271inter8));
  nand2 gate1578(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1579(.a(s_147), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1580(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1581(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1582(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2059(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2060(.a(gate277inter0), .b(s_216), .O(gate277inter1));
  and2  gate2061(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2062(.a(s_216), .O(gate277inter3));
  inv1  gate2063(.a(s_217), .O(gate277inter4));
  nand2 gate2064(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2065(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2066(.a(G648), .O(gate277inter7));
  inv1  gate2067(.a(G800), .O(gate277inter8));
  nand2 gate2068(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2069(.a(s_217), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2070(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2071(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2072(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate2619(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2620(.a(gate278inter0), .b(s_296), .O(gate278inter1));
  and2  gate2621(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2622(.a(s_296), .O(gate278inter3));
  inv1  gate2623(.a(s_297), .O(gate278inter4));
  nand2 gate2624(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2625(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2626(.a(G776), .O(gate278inter7));
  inv1  gate2627(.a(G800), .O(gate278inter8));
  nand2 gate2628(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2629(.a(s_297), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2630(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2631(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2632(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2759(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2760(.a(gate280inter0), .b(s_316), .O(gate280inter1));
  and2  gate2761(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2762(.a(s_316), .O(gate280inter3));
  inv1  gate2763(.a(s_317), .O(gate280inter4));
  nand2 gate2764(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2765(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2766(.a(G779), .O(gate280inter7));
  inv1  gate2767(.a(G803), .O(gate280inter8));
  nand2 gate2768(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2769(.a(s_317), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2770(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2771(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2772(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate631(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate632(.a(gate289inter0), .b(s_12), .O(gate289inter1));
  and2  gate633(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate634(.a(s_12), .O(gate289inter3));
  inv1  gate635(.a(s_13), .O(gate289inter4));
  nand2 gate636(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate637(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate638(.a(G818), .O(gate289inter7));
  inv1  gate639(.a(G819), .O(gate289inter8));
  nand2 gate640(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate641(.a(s_13), .b(gate289inter3), .O(gate289inter10));
  nor2  gate642(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate643(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate644(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2129(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2130(.a(gate291inter0), .b(s_226), .O(gate291inter1));
  and2  gate2131(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2132(.a(s_226), .O(gate291inter3));
  inv1  gate2133(.a(s_227), .O(gate291inter4));
  nand2 gate2134(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2135(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2136(.a(G822), .O(gate291inter7));
  inv1  gate2137(.a(G823), .O(gate291inter8));
  nand2 gate2138(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2139(.a(s_227), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2140(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2141(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2142(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1681(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1682(.a(gate391inter0), .b(s_162), .O(gate391inter1));
  and2  gate1683(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1684(.a(s_162), .O(gate391inter3));
  inv1  gate1685(.a(s_163), .O(gate391inter4));
  nand2 gate1686(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1687(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1688(.a(G5), .O(gate391inter7));
  inv1  gate1689(.a(G1048), .O(gate391inter8));
  nand2 gate1690(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1691(.a(s_163), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1692(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1693(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1694(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2689(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2690(.a(gate393inter0), .b(s_306), .O(gate393inter1));
  and2  gate2691(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2692(.a(s_306), .O(gate393inter3));
  inv1  gate2693(.a(s_307), .O(gate393inter4));
  nand2 gate2694(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2695(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2696(.a(G7), .O(gate393inter7));
  inv1  gate2697(.a(G1054), .O(gate393inter8));
  nand2 gate2698(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2699(.a(s_307), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2700(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2701(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2702(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate589(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate590(.a(gate396inter0), .b(s_6), .O(gate396inter1));
  and2  gate591(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate592(.a(s_6), .O(gate396inter3));
  inv1  gate593(.a(s_7), .O(gate396inter4));
  nand2 gate594(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate595(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate596(.a(G10), .O(gate396inter7));
  inv1  gate597(.a(G1063), .O(gate396inter8));
  nand2 gate598(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate599(.a(s_7), .b(gate396inter3), .O(gate396inter10));
  nor2  gate600(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate601(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate602(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate2675(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2676(.a(gate397inter0), .b(s_304), .O(gate397inter1));
  and2  gate2677(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2678(.a(s_304), .O(gate397inter3));
  inv1  gate2679(.a(s_305), .O(gate397inter4));
  nand2 gate2680(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2681(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2682(.a(G11), .O(gate397inter7));
  inv1  gate2683(.a(G1066), .O(gate397inter8));
  nand2 gate2684(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2685(.a(s_305), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2686(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2687(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2688(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1163(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1164(.a(gate398inter0), .b(s_88), .O(gate398inter1));
  and2  gate1165(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1166(.a(s_88), .O(gate398inter3));
  inv1  gate1167(.a(s_89), .O(gate398inter4));
  nand2 gate1168(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1169(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1170(.a(G12), .O(gate398inter7));
  inv1  gate1171(.a(G1069), .O(gate398inter8));
  nand2 gate1172(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1173(.a(s_89), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1174(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1175(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1176(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1373(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1374(.a(gate402inter0), .b(s_118), .O(gate402inter1));
  and2  gate1375(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1376(.a(s_118), .O(gate402inter3));
  inv1  gate1377(.a(s_119), .O(gate402inter4));
  nand2 gate1378(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1379(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1380(.a(G16), .O(gate402inter7));
  inv1  gate1381(.a(G1081), .O(gate402inter8));
  nand2 gate1382(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1383(.a(s_119), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1384(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1385(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1386(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1275(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1276(.a(gate403inter0), .b(s_104), .O(gate403inter1));
  and2  gate1277(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1278(.a(s_104), .O(gate403inter3));
  inv1  gate1279(.a(s_105), .O(gate403inter4));
  nand2 gate1280(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1281(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1282(.a(G17), .O(gate403inter7));
  inv1  gate1283(.a(G1084), .O(gate403inter8));
  nand2 gate1284(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1285(.a(s_105), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1286(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1287(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1288(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate561(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate562(.a(gate404inter0), .b(s_2), .O(gate404inter1));
  and2  gate563(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate564(.a(s_2), .O(gate404inter3));
  inv1  gate565(.a(s_3), .O(gate404inter4));
  nand2 gate566(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate567(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate568(.a(G18), .O(gate404inter7));
  inv1  gate569(.a(G1087), .O(gate404inter8));
  nand2 gate570(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate571(.a(s_3), .b(gate404inter3), .O(gate404inter10));
  nor2  gate572(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate573(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate574(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1597(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1598(.a(gate410inter0), .b(s_150), .O(gate410inter1));
  and2  gate1599(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1600(.a(s_150), .O(gate410inter3));
  inv1  gate1601(.a(s_151), .O(gate410inter4));
  nand2 gate1602(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1603(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1604(.a(G24), .O(gate410inter7));
  inv1  gate1605(.a(G1105), .O(gate410inter8));
  nand2 gate1606(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1607(.a(s_151), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1608(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1609(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1610(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2731(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2732(.a(gate412inter0), .b(s_312), .O(gate412inter1));
  and2  gate2733(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2734(.a(s_312), .O(gate412inter3));
  inv1  gate2735(.a(s_313), .O(gate412inter4));
  nand2 gate2736(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2737(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2738(.a(G26), .O(gate412inter7));
  inv1  gate2739(.a(G1111), .O(gate412inter8));
  nand2 gate2740(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2741(.a(s_313), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2742(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2743(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2744(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1583(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1584(.a(gate416inter0), .b(s_148), .O(gate416inter1));
  and2  gate1585(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1586(.a(s_148), .O(gate416inter3));
  inv1  gate1587(.a(s_149), .O(gate416inter4));
  nand2 gate1588(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1589(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1590(.a(G30), .O(gate416inter7));
  inv1  gate1591(.a(G1123), .O(gate416inter8));
  nand2 gate1592(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1593(.a(s_149), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1594(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1595(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1596(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate659(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate660(.a(gate422inter0), .b(s_16), .O(gate422inter1));
  and2  gate661(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate662(.a(s_16), .O(gate422inter3));
  inv1  gate663(.a(s_17), .O(gate422inter4));
  nand2 gate664(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate665(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate666(.a(G1039), .O(gate422inter7));
  inv1  gate667(.a(G1135), .O(gate422inter8));
  nand2 gate668(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate669(.a(s_17), .b(gate422inter3), .O(gate422inter10));
  nor2  gate670(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate671(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate672(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1079(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1080(.a(gate423inter0), .b(s_76), .O(gate423inter1));
  and2  gate1081(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1082(.a(s_76), .O(gate423inter3));
  inv1  gate1083(.a(s_77), .O(gate423inter4));
  nand2 gate1084(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1085(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1086(.a(G3), .O(gate423inter7));
  inv1  gate1087(.a(G1138), .O(gate423inter8));
  nand2 gate1088(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1089(.a(s_77), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1090(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1091(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1092(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1121(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1122(.a(gate425inter0), .b(s_82), .O(gate425inter1));
  and2  gate1123(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1124(.a(s_82), .O(gate425inter3));
  inv1  gate1125(.a(s_83), .O(gate425inter4));
  nand2 gate1126(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1127(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1128(.a(G4), .O(gate425inter7));
  inv1  gate1129(.a(G1141), .O(gate425inter8));
  nand2 gate1130(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1131(.a(s_83), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1132(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1133(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1134(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1821(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1822(.a(gate427inter0), .b(s_182), .O(gate427inter1));
  and2  gate1823(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1824(.a(s_182), .O(gate427inter3));
  inv1  gate1825(.a(s_183), .O(gate427inter4));
  nand2 gate1826(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1827(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1828(.a(G5), .O(gate427inter7));
  inv1  gate1829(.a(G1144), .O(gate427inter8));
  nand2 gate1830(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1831(.a(s_183), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1832(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1833(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1834(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1863(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1864(.a(gate428inter0), .b(s_188), .O(gate428inter1));
  and2  gate1865(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1866(.a(s_188), .O(gate428inter3));
  inv1  gate1867(.a(s_189), .O(gate428inter4));
  nand2 gate1868(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1869(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1870(.a(G1048), .O(gate428inter7));
  inv1  gate1871(.a(G1144), .O(gate428inter8));
  nand2 gate1872(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1873(.a(s_189), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1874(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1875(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1876(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1667(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1668(.a(gate431inter0), .b(s_160), .O(gate431inter1));
  and2  gate1669(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1670(.a(s_160), .O(gate431inter3));
  inv1  gate1671(.a(s_161), .O(gate431inter4));
  nand2 gate1672(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1673(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1674(.a(G7), .O(gate431inter7));
  inv1  gate1675(.a(G1150), .O(gate431inter8));
  nand2 gate1676(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1677(.a(s_161), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1678(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1679(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1680(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1919(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1920(.a(gate433inter0), .b(s_196), .O(gate433inter1));
  and2  gate1921(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1922(.a(s_196), .O(gate433inter3));
  inv1  gate1923(.a(s_197), .O(gate433inter4));
  nand2 gate1924(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1925(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1926(.a(G8), .O(gate433inter7));
  inv1  gate1927(.a(G1153), .O(gate433inter8));
  nand2 gate1928(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1929(.a(s_197), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1930(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1931(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1932(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1289(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1290(.a(gate434inter0), .b(s_106), .O(gate434inter1));
  and2  gate1291(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1292(.a(s_106), .O(gate434inter3));
  inv1  gate1293(.a(s_107), .O(gate434inter4));
  nand2 gate1294(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1295(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1296(.a(G1057), .O(gate434inter7));
  inv1  gate1297(.a(G1153), .O(gate434inter8));
  nand2 gate1298(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1299(.a(s_107), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1300(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1301(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1302(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2185(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2186(.a(gate442inter0), .b(s_234), .O(gate442inter1));
  and2  gate2187(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2188(.a(s_234), .O(gate442inter3));
  inv1  gate2189(.a(s_235), .O(gate442inter4));
  nand2 gate2190(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2191(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2192(.a(G1069), .O(gate442inter7));
  inv1  gate2193(.a(G1165), .O(gate442inter8));
  nand2 gate2194(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2195(.a(s_235), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2196(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2197(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2198(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate687(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate688(.a(gate444inter0), .b(s_20), .O(gate444inter1));
  and2  gate689(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate690(.a(s_20), .O(gate444inter3));
  inv1  gate691(.a(s_21), .O(gate444inter4));
  nand2 gate692(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate693(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate694(.a(G1072), .O(gate444inter7));
  inv1  gate695(.a(G1168), .O(gate444inter8));
  nand2 gate696(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate697(.a(s_21), .b(gate444inter3), .O(gate444inter10));
  nor2  gate698(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate699(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate700(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1191(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1192(.a(gate446inter0), .b(s_92), .O(gate446inter1));
  and2  gate1193(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1194(.a(s_92), .O(gate446inter3));
  inv1  gate1195(.a(s_93), .O(gate446inter4));
  nand2 gate1196(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1197(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1198(.a(G1075), .O(gate446inter7));
  inv1  gate1199(.a(G1171), .O(gate446inter8));
  nand2 gate1200(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1201(.a(s_93), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1202(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1203(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1204(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1793(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1794(.a(gate448inter0), .b(s_178), .O(gate448inter1));
  and2  gate1795(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1796(.a(s_178), .O(gate448inter3));
  inv1  gate1797(.a(s_179), .O(gate448inter4));
  nand2 gate1798(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1799(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1800(.a(G1078), .O(gate448inter7));
  inv1  gate1801(.a(G1174), .O(gate448inter8));
  nand2 gate1802(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1803(.a(s_179), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1804(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1805(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1806(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1051(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1052(.a(gate451inter0), .b(s_72), .O(gate451inter1));
  and2  gate1053(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1054(.a(s_72), .O(gate451inter3));
  inv1  gate1055(.a(s_73), .O(gate451inter4));
  nand2 gate1056(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1057(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1058(.a(G17), .O(gate451inter7));
  inv1  gate1059(.a(G1180), .O(gate451inter8));
  nand2 gate1060(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1061(.a(s_73), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1062(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1063(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1064(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1723(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1724(.a(gate453inter0), .b(s_168), .O(gate453inter1));
  and2  gate1725(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1726(.a(s_168), .O(gate453inter3));
  inv1  gate1727(.a(s_169), .O(gate453inter4));
  nand2 gate1728(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1729(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1730(.a(G18), .O(gate453inter7));
  inv1  gate1731(.a(G1183), .O(gate453inter8));
  nand2 gate1732(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1733(.a(s_169), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1734(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1735(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1736(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2703(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2704(.a(gate456inter0), .b(s_308), .O(gate456inter1));
  and2  gate2705(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2706(.a(s_308), .O(gate456inter3));
  inv1  gate2707(.a(s_309), .O(gate456inter4));
  nand2 gate2708(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2709(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2710(.a(G1090), .O(gate456inter7));
  inv1  gate2711(.a(G1186), .O(gate456inter8));
  nand2 gate2712(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2713(.a(s_309), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2714(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2715(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2716(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1177(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1178(.a(gate457inter0), .b(s_90), .O(gate457inter1));
  and2  gate1179(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1180(.a(s_90), .O(gate457inter3));
  inv1  gate1181(.a(s_91), .O(gate457inter4));
  nand2 gate1182(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1183(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1184(.a(G20), .O(gate457inter7));
  inv1  gate1185(.a(G1189), .O(gate457inter8));
  nand2 gate1186(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1187(.a(s_91), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1188(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1189(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1190(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1023(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1024(.a(gate461inter0), .b(s_68), .O(gate461inter1));
  and2  gate1025(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1026(.a(s_68), .O(gate461inter3));
  inv1  gate1027(.a(s_69), .O(gate461inter4));
  nand2 gate1028(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1029(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1030(.a(G22), .O(gate461inter7));
  inv1  gate1031(.a(G1195), .O(gate461inter8));
  nand2 gate1032(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1033(.a(s_69), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1034(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1035(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1036(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1359(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1360(.a(gate465inter0), .b(s_116), .O(gate465inter1));
  and2  gate1361(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1362(.a(s_116), .O(gate465inter3));
  inv1  gate1363(.a(s_117), .O(gate465inter4));
  nand2 gate1364(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1365(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1366(.a(G24), .O(gate465inter7));
  inv1  gate1367(.a(G1201), .O(gate465inter8));
  nand2 gate1368(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1369(.a(s_117), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1370(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1371(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1372(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1219(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1220(.a(gate470inter0), .b(s_96), .O(gate470inter1));
  and2  gate1221(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1222(.a(s_96), .O(gate470inter3));
  inv1  gate1223(.a(s_97), .O(gate470inter4));
  nand2 gate1224(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1225(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1226(.a(G1111), .O(gate470inter7));
  inv1  gate1227(.a(G1207), .O(gate470inter8));
  nand2 gate1228(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1229(.a(s_97), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1230(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1231(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1232(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate771(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate772(.a(gate471inter0), .b(s_32), .O(gate471inter1));
  and2  gate773(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate774(.a(s_32), .O(gate471inter3));
  inv1  gate775(.a(s_33), .O(gate471inter4));
  nand2 gate776(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate777(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate778(.a(G27), .O(gate471inter7));
  inv1  gate779(.a(G1210), .O(gate471inter8));
  nand2 gate780(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate781(.a(s_33), .b(gate471inter3), .O(gate471inter10));
  nor2  gate782(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate783(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate784(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1709(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1710(.a(gate473inter0), .b(s_166), .O(gate473inter1));
  and2  gate1711(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1712(.a(s_166), .O(gate473inter3));
  inv1  gate1713(.a(s_167), .O(gate473inter4));
  nand2 gate1714(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1715(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1716(.a(G28), .O(gate473inter7));
  inv1  gate1717(.a(G1213), .O(gate473inter8));
  nand2 gate1718(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1719(.a(s_167), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1720(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1721(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1722(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2143(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2144(.a(gate475inter0), .b(s_228), .O(gate475inter1));
  and2  gate2145(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2146(.a(s_228), .O(gate475inter3));
  inv1  gate2147(.a(s_229), .O(gate475inter4));
  nand2 gate2148(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2149(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2150(.a(G29), .O(gate475inter7));
  inv1  gate2151(.a(G1216), .O(gate475inter8));
  nand2 gate2152(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2153(.a(s_229), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2154(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2155(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2156(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate547(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate548(.a(gate479inter0), .b(s_0), .O(gate479inter1));
  and2  gate549(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate550(.a(s_0), .O(gate479inter3));
  inv1  gate551(.a(s_1), .O(gate479inter4));
  nand2 gate552(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate553(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate554(.a(G31), .O(gate479inter7));
  inv1  gate555(.a(G1222), .O(gate479inter8));
  nand2 gate556(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate557(.a(s_1), .b(gate479inter3), .O(gate479inter10));
  nor2  gate558(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate559(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate560(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1107(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1108(.a(gate480inter0), .b(s_80), .O(gate480inter1));
  and2  gate1109(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1110(.a(s_80), .O(gate480inter3));
  inv1  gate1111(.a(s_81), .O(gate480inter4));
  nand2 gate1112(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1113(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1114(.a(G1126), .O(gate480inter7));
  inv1  gate1115(.a(G1222), .O(gate480inter8));
  nand2 gate1116(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1117(.a(s_81), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1118(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1119(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1120(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2199(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2200(.a(gate482inter0), .b(s_236), .O(gate482inter1));
  and2  gate2201(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2202(.a(s_236), .O(gate482inter3));
  inv1  gate2203(.a(s_237), .O(gate482inter4));
  nand2 gate2204(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2205(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2206(.a(G1129), .O(gate482inter7));
  inv1  gate2207(.a(G1225), .O(gate482inter8));
  nand2 gate2208(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2209(.a(s_237), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2210(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2211(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2212(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1975(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1976(.a(gate484inter0), .b(s_204), .O(gate484inter1));
  and2  gate1977(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1978(.a(s_204), .O(gate484inter3));
  inv1  gate1979(.a(s_205), .O(gate484inter4));
  nand2 gate1980(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1981(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1982(.a(G1230), .O(gate484inter7));
  inv1  gate1983(.a(G1231), .O(gate484inter8));
  nand2 gate1984(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1985(.a(s_205), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1986(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1987(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1988(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2465(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2466(.a(gate488inter0), .b(s_274), .O(gate488inter1));
  and2  gate2467(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2468(.a(s_274), .O(gate488inter3));
  inv1  gate2469(.a(s_275), .O(gate488inter4));
  nand2 gate2470(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2471(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2472(.a(G1238), .O(gate488inter7));
  inv1  gate2473(.a(G1239), .O(gate488inter8));
  nand2 gate2474(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2475(.a(s_275), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2476(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2477(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2478(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate2367(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2368(.a(gate489inter0), .b(s_260), .O(gate489inter1));
  and2  gate2369(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2370(.a(s_260), .O(gate489inter3));
  inv1  gate2371(.a(s_261), .O(gate489inter4));
  nand2 gate2372(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2373(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2374(.a(G1240), .O(gate489inter7));
  inv1  gate2375(.a(G1241), .O(gate489inter8));
  nand2 gate2376(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2377(.a(s_261), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2378(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2379(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2380(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2031(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2032(.a(gate491inter0), .b(s_212), .O(gate491inter1));
  and2  gate2033(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2034(.a(s_212), .O(gate491inter3));
  inv1  gate2035(.a(s_213), .O(gate491inter4));
  nand2 gate2036(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2037(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2038(.a(G1244), .O(gate491inter7));
  inv1  gate2039(.a(G1245), .O(gate491inter8));
  nand2 gate2040(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2041(.a(s_213), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2042(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2043(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2044(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate603(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate604(.a(gate492inter0), .b(s_8), .O(gate492inter1));
  and2  gate605(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate606(.a(s_8), .O(gate492inter3));
  inv1  gate607(.a(s_9), .O(gate492inter4));
  nand2 gate608(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate609(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate610(.a(G1246), .O(gate492inter7));
  inv1  gate611(.a(G1247), .O(gate492inter8));
  nand2 gate612(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate613(.a(s_9), .b(gate492inter3), .O(gate492inter10));
  nor2  gate614(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate615(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate616(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1037(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1038(.a(gate493inter0), .b(s_70), .O(gate493inter1));
  and2  gate1039(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1040(.a(s_70), .O(gate493inter3));
  inv1  gate1041(.a(s_71), .O(gate493inter4));
  nand2 gate1042(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1043(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1044(.a(G1248), .O(gate493inter7));
  inv1  gate1045(.a(G1249), .O(gate493inter8));
  nand2 gate1046(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1047(.a(s_71), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1048(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1049(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1050(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate869(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate870(.a(gate494inter0), .b(s_46), .O(gate494inter1));
  and2  gate871(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate872(.a(s_46), .O(gate494inter3));
  inv1  gate873(.a(s_47), .O(gate494inter4));
  nand2 gate874(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate875(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate876(.a(G1250), .O(gate494inter7));
  inv1  gate877(.a(G1251), .O(gate494inter8));
  nand2 gate878(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate879(.a(s_47), .b(gate494inter3), .O(gate494inter10));
  nor2  gate880(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate881(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate882(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2003(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2004(.a(gate496inter0), .b(s_208), .O(gate496inter1));
  and2  gate2005(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2006(.a(s_208), .O(gate496inter3));
  inv1  gate2007(.a(s_209), .O(gate496inter4));
  nand2 gate2008(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2009(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2010(.a(G1254), .O(gate496inter7));
  inv1  gate2011(.a(G1255), .O(gate496inter8));
  nand2 gate2012(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2013(.a(s_209), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2014(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2015(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2016(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate813(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate814(.a(gate498inter0), .b(s_38), .O(gate498inter1));
  and2  gate815(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate816(.a(s_38), .O(gate498inter3));
  inv1  gate817(.a(s_39), .O(gate498inter4));
  nand2 gate818(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate819(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate820(.a(G1258), .O(gate498inter7));
  inv1  gate821(.a(G1259), .O(gate498inter8));
  nand2 gate822(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate823(.a(s_39), .b(gate498inter3), .O(gate498inter10));
  nor2  gate824(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate825(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate826(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1807(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1808(.a(gate499inter0), .b(s_180), .O(gate499inter1));
  and2  gate1809(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1810(.a(s_180), .O(gate499inter3));
  inv1  gate1811(.a(s_181), .O(gate499inter4));
  nand2 gate1812(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1813(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1814(.a(G1260), .O(gate499inter7));
  inv1  gate1815(.a(G1261), .O(gate499inter8));
  nand2 gate1816(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1817(.a(s_181), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1818(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1819(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1820(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1261(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1262(.a(gate503inter0), .b(s_102), .O(gate503inter1));
  and2  gate1263(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1264(.a(s_102), .O(gate503inter3));
  inv1  gate1265(.a(s_103), .O(gate503inter4));
  nand2 gate1266(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1267(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1268(.a(G1268), .O(gate503inter7));
  inv1  gate1269(.a(G1269), .O(gate503inter8));
  nand2 gate1270(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1271(.a(s_103), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1272(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1273(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1274(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate1513(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1514(.a(gate504inter0), .b(s_138), .O(gate504inter1));
  and2  gate1515(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1516(.a(s_138), .O(gate504inter3));
  inv1  gate1517(.a(s_139), .O(gate504inter4));
  nand2 gate1518(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1519(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1520(.a(G1270), .O(gate504inter7));
  inv1  gate1521(.a(G1271), .O(gate504inter8));
  nand2 gate1522(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1523(.a(s_139), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1524(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1525(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1526(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1345(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1346(.a(gate506inter0), .b(s_114), .O(gate506inter1));
  and2  gate1347(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1348(.a(s_114), .O(gate506inter3));
  inv1  gate1349(.a(s_115), .O(gate506inter4));
  nand2 gate1350(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1351(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1352(.a(G1274), .O(gate506inter7));
  inv1  gate1353(.a(G1275), .O(gate506inter8));
  nand2 gate1354(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1355(.a(s_115), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1356(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1357(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1358(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate2241(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2242(.a(gate507inter0), .b(s_242), .O(gate507inter1));
  and2  gate2243(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2244(.a(s_242), .O(gate507inter3));
  inv1  gate2245(.a(s_243), .O(gate507inter4));
  nand2 gate2246(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2247(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2248(.a(G1276), .O(gate507inter7));
  inv1  gate2249(.a(G1277), .O(gate507inter8));
  nand2 gate2250(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2251(.a(s_243), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2252(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2253(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2254(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate981(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate982(.a(gate508inter0), .b(s_62), .O(gate508inter1));
  and2  gate983(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate984(.a(s_62), .O(gate508inter3));
  inv1  gate985(.a(s_63), .O(gate508inter4));
  nand2 gate986(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate987(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate988(.a(G1278), .O(gate508inter7));
  inv1  gate989(.a(G1279), .O(gate508inter8));
  nand2 gate990(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate991(.a(s_63), .b(gate508inter3), .O(gate508inter10));
  nor2  gate992(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate993(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate994(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1233(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1234(.a(gate513inter0), .b(s_98), .O(gate513inter1));
  and2  gate1235(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1236(.a(s_98), .O(gate513inter3));
  inv1  gate1237(.a(s_99), .O(gate513inter4));
  nand2 gate1238(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1239(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1240(.a(G1288), .O(gate513inter7));
  inv1  gate1241(.a(G1289), .O(gate513inter8));
  nand2 gate1242(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1243(.a(s_99), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1244(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1245(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1246(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule