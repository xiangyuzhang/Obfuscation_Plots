module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1737(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1738(.a(gate10inter0), .b(s_170), .O(gate10inter1));
  and2  gate1739(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1740(.a(s_170), .O(gate10inter3));
  inv1  gate1741(.a(s_171), .O(gate10inter4));
  nand2 gate1742(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1743(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1744(.a(G3), .O(gate10inter7));
  inv1  gate1745(.a(G4), .O(gate10inter8));
  nand2 gate1746(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1747(.a(s_171), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1748(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1749(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1750(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1695(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1696(.a(gate16inter0), .b(s_164), .O(gate16inter1));
  and2  gate1697(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1698(.a(s_164), .O(gate16inter3));
  inv1  gate1699(.a(s_165), .O(gate16inter4));
  nand2 gate1700(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1701(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1702(.a(G15), .O(gate16inter7));
  inv1  gate1703(.a(G16), .O(gate16inter8));
  nand2 gate1704(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1705(.a(s_165), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1706(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1707(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1708(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1639(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1640(.a(gate20inter0), .b(s_156), .O(gate20inter1));
  and2  gate1641(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1642(.a(s_156), .O(gate20inter3));
  inv1  gate1643(.a(s_157), .O(gate20inter4));
  nand2 gate1644(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1645(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1646(.a(G23), .O(gate20inter7));
  inv1  gate1647(.a(G24), .O(gate20inter8));
  nand2 gate1648(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1649(.a(s_157), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1650(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1651(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1652(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1863(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1864(.a(gate29inter0), .b(s_188), .O(gate29inter1));
  and2  gate1865(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1866(.a(s_188), .O(gate29inter3));
  inv1  gate1867(.a(s_189), .O(gate29inter4));
  nand2 gate1868(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1869(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1870(.a(G3), .O(gate29inter7));
  inv1  gate1871(.a(G7), .O(gate29inter8));
  nand2 gate1872(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1873(.a(s_189), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1874(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1875(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1876(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate785(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate786(.a(gate31inter0), .b(s_34), .O(gate31inter1));
  and2  gate787(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate788(.a(s_34), .O(gate31inter3));
  inv1  gate789(.a(s_35), .O(gate31inter4));
  nand2 gate790(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate791(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate792(.a(G4), .O(gate31inter7));
  inv1  gate793(.a(G8), .O(gate31inter8));
  nand2 gate794(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate795(.a(s_35), .b(gate31inter3), .O(gate31inter10));
  nor2  gate796(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate797(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate798(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1513(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1514(.a(gate32inter0), .b(s_138), .O(gate32inter1));
  and2  gate1515(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1516(.a(s_138), .O(gate32inter3));
  inv1  gate1517(.a(s_139), .O(gate32inter4));
  nand2 gate1518(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1519(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1520(.a(G12), .O(gate32inter7));
  inv1  gate1521(.a(G16), .O(gate32inter8));
  nand2 gate1522(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1523(.a(s_139), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1524(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1525(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1526(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2213(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2214(.a(gate34inter0), .b(s_238), .O(gate34inter1));
  and2  gate2215(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2216(.a(s_238), .O(gate34inter3));
  inv1  gate2217(.a(s_239), .O(gate34inter4));
  nand2 gate2218(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2219(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2220(.a(G25), .O(gate34inter7));
  inv1  gate2221(.a(G29), .O(gate34inter8));
  nand2 gate2222(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2223(.a(s_239), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2224(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2225(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2226(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate981(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate982(.a(gate35inter0), .b(s_62), .O(gate35inter1));
  and2  gate983(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate984(.a(s_62), .O(gate35inter3));
  inv1  gate985(.a(s_63), .O(gate35inter4));
  nand2 gate986(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate987(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate988(.a(G18), .O(gate35inter7));
  inv1  gate989(.a(G22), .O(gate35inter8));
  nand2 gate990(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate991(.a(s_63), .b(gate35inter3), .O(gate35inter10));
  nor2  gate992(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate993(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate994(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1527(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1528(.a(gate40inter0), .b(s_140), .O(gate40inter1));
  and2  gate1529(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1530(.a(s_140), .O(gate40inter3));
  inv1  gate1531(.a(s_141), .O(gate40inter4));
  nand2 gate1532(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1533(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1534(.a(G28), .O(gate40inter7));
  inv1  gate1535(.a(G32), .O(gate40inter8));
  nand2 gate1536(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1537(.a(s_141), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1538(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1539(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1540(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1821(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1822(.a(gate42inter0), .b(s_182), .O(gate42inter1));
  and2  gate1823(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1824(.a(s_182), .O(gate42inter3));
  inv1  gate1825(.a(s_183), .O(gate42inter4));
  nand2 gate1826(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1827(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1828(.a(G2), .O(gate42inter7));
  inv1  gate1829(.a(G266), .O(gate42inter8));
  nand2 gate1830(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1831(.a(s_183), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1832(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1833(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1834(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1107(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1108(.a(gate45inter0), .b(s_80), .O(gate45inter1));
  and2  gate1109(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1110(.a(s_80), .O(gate45inter3));
  inv1  gate1111(.a(s_81), .O(gate45inter4));
  nand2 gate1112(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1113(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1114(.a(G5), .O(gate45inter7));
  inv1  gate1115(.a(G272), .O(gate45inter8));
  nand2 gate1116(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1117(.a(s_81), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1118(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1119(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1120(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate2157(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2158(.a(gate46inter0), .b(s_230), .O(gate46inter1));
  and2  gate2159(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2160(.a(s_230), .O(gate46inter3));
  inv1  gate2161(.a(s_231), .O(gate46inter4));
  nand2 gate2162(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2163(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2164(.a(G6), .O(gate46inter7));
  inv1  gate2165(.a(G272), .O(gate46inter8));
  nand2 gate2166(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2167(.a(s_231), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2168(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2169(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2170(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate911(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate912(.a(gate48inter0), .b(s_52), .O(gate48inter1));
  and2  gate913(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate914(.a(s_52), .O(gate48inter3));
  inv1  gate915(.a(s_53), .O(gate48inter4));
  nand2 gate916(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate917(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate918(.a(G8), .O(gate48inter7));
  inv1  gate919(.a(G275), .O(gate48inter8));
  nand2 gate920(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate921(.a(s_53), .b(gate48inter3), .O(gate48inter10));
  nor2  gate922(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate923(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate924(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate589(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate590(.a(gate49inter0), .b(s_6), .O(gate49inter1));
  and2  gate591(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate592(.a(s_6), .O(gate49inter3));
  inv1  gate593(.a(s_7), .O(gate49inter4));
  nand2 gate594(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate595(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate596(.a(G9), .O(gate49inter7));
  inv1  gate597(.a(G278), .O(gate49inter8));
  nand2 gate598(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate599(.a(s_7), .b(gate49inter3), .O(gate49inter10));
  nor2  gate600(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate601(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate602(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1247(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1248(.a(gate51inter0), .b(s_100), .O(gate51inter1));
  and2  gate1249(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1250(.a(s_100), .O(gate51inter3));
  inv1  gate1251(.a(s_101), .O(gate51inter4));
  nand2 gate1252(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1253(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1254(.a(G11), .O(gate51inter7));
  inv1  gate1255(.a(G281), .O(gate51inter8));
  nand2 gate1256(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1257(.a(s_101), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1258(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1259(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1260(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1121(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1122(.a(gate57inter0), .b(s_82), .O(gate57inter1));
  and2  gate1123(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1124(.a(s_82), .O(gate57inter3));
  inv1  gate1125(.a(s_83), .O(gate57inter4));
  nand2 gate1126(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1127(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1128(.a(G17), .O(gate57inter7));
  inv1  gate1129(.a(G290), .O(gate57inter8));
  nand2 gate1130(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1131(.a(s_83), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1132(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1133(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1134(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1471(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1472(.a(gate62inter0), .b(s_132), .O(gate62inter1));
  and2  gate1473(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1474(.a(s_132), .O(gate62inter3));
  inv1  gate1475(.a(s_133), .O(gate62inter4));
  nand2 gate1476(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1477(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1478(.a(G22), .O(gate62inter7));
  inv1  gate1479(.a(G296), .O(gate62inter8));
  nand2 gate1480(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1481(.a(s_133), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1482(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1483(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1484(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate715(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate716(.a(gate66inter0), .b(s_24), .O(gate66inter1));
  and2  gate717(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate718(.a(s_24), .O(gate66inter3));
  inv1  gate719(.a(s_25), .O(gate66inter4));
  nand2 gate720(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate721(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate722(.a(G26), .O(gate66inter7));
  inv1  gate723(.a(G302), .O(gate66inter8));
  nand2 gate724(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate725(.a(s_25), .b(gate66inter3), .O(gate66inter10));
  nor2  gate726(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate727(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate728(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate897(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate898(.a(gate70inter0), .b(s_50), .O(gate70inter1));
  and2  gate899(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate900(.a(s_50), .O(gate70inter3));
  inv1  gate901(.a(s_51), .O(gate70inter4));
  nand2 gate902(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate903(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate904(.a(G30), .O(gate70inter7));
  inv1  gate905(.a(G308), .O(gate70inter8));
  nand2 gate906(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate907(.a(s_51), .b(gate70inter3), .O(gate70inter10));
  nor2  gate908(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate909(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate910(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1975(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1976(.a(gate71inter0), .b(s_204), .O(gate71inter1));
  and2  gate1977(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1978(.a(s_204), .O(gate71inter3));
  inv1  gate1979(.a(s_205), .O(gate71inter4));
  nand2 gate1980(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1981(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1982(.a(G31), .O(gate71inter7));
  inv1  gate1983(.a(G311), .O(gate71inter8));
  nand2 gate1984(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1985(.a(s_205), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1986(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1987(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1988(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2115(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2116(.a(gate72inter0), .b(s_224), .O(gate72inter1));
  and2  gate2117(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2118(.a(s_224), .O(gate72inter3));
  inv1  gate2119(.a(s_225), .O(gate72inter4));
  nand2 gate2120(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2121(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2122(.a(G32), .O(gate72inter7));
  inv1  gate2123(.a(G311), .O(gate72inter8));
  nand2 gate2124(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2125(.a(s_225), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2126(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2127(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2128(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1877(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1878(.a(gate73inter0), .b(s_190), .O(gate73inter1));
  and2  gate1879(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1880(.a(s_190), .O(gate73inter3));
  inv1  gate1881(.a(s_191), .O(gate73inter4));
  nand2 gate1882(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1883(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1884(.a(G1), .O(gate73inter7));
  inv1  gate1885(.a(G314), .O(gate73inter8));
  nand2 gate1886(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1887(.a(s_191), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1888(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1889(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1890(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate673(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate674(.a(gate74inter0), .b(s_18), .O(gate74inter1));
  and2  gate675(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate676(.a(s_18), .O(gate74inter3));
  inv1  gate677(.a(s_19), .O(gate74inter4));
  nand2 gate678(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate679(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate680(.a(G5), .O(gate74inter7));
  inv1  gate681(.a(G314), .O(gate74inter8));
  nand2 gate682(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate683(.a(s_19), .b(gate74inter3), .O(gate74inter10));
  nor2  gate684(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate685(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate686(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1905(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1906(.a(gate76inter0), .b(s_194), .O(gate76inter1));
  and2  gate1907(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1908(.a(s_194), .O(gate76inter3));
  inv1  gate1909(.a(s_195), .O(gate76inter4));
  nand2 gate1910(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1911(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1912(.a(G13), .O(gate76inter7));
  inv1  gate1913(.a(G317), .O(gate76inter8));
  nand2 gate1914(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1915(.a(s_195), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1916(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1917(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1918(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate617(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate618(.a(gate78inter0), .b(s_10), .O(gate78inter1));
  and2  gate619(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate620(.a(s_10), .O(gate78inter3));
  inv1  gate621(.a(s_11), .O(gate78inter4));
  nand2 gate622(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate623(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate624(.a(G6), .O(gate78inter7));
  inv1  gate625(.a(G320), .O(gate78inter8));
  nand2 gate626(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate627(.a(s_11), .b(gate78inter3), .O(gate78inter10));
  nor2  gate628(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate629(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate630(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1779(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1780(.a(gate80inter0), .b(s_176), .O(gate80inter1));
  and2  gate1781(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1782(.a(s_176), .O(gate80inter3));
  inv1  gate1783(.a(s_177), .O(gate80inter4));
  nand2 gate1784(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1785(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1786(.a(G14), .O(gate80inter7));
  inv1  gate1787(.a(G323), .O(gate80inter8));
  nand2 gate1788(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1789(.a(s_177), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1790(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1791(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1792(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1149(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1150(.a(gate81inter0), .b(s_86), .O(gate81inter1));
  and2  gate1151(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1152(.a(s_86), .O(gate81inter3));
  inv1  gate1153(.a(s_87), .O(gate81inter4));
  nand2 gate1154(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1155(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1156(.a(G3), .O(gate81inter7));
  inv1  gate1157(.a(G326), .O(gate81inter8));
  nand2 gate1158(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1159(.a(s_87), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1160(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1161(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1162(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate2045(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2046(.a(gate82inter0), .b(s_214), .O(gate82inter1));
  and2  gate2047(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2048(.a(s_214), .O(gate82inter3));
  inv1  gate2049(.a(s_215), .O(gate82inter4));
  nand2 gate2050(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2051(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2052(.a(G7), .O(gate82inter7));
  inv1  gate2053(.a(G326), .O(gate82inter8));
  nand2 gate2054(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2055(.a(s_215), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2056(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2057(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2058(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1289(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1290(.a(gate86inter0), .b(s_106), .O(gate86inter1));
  and2  gate1291(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1292(.a(s_106), .O(gate86inter3));
  inv1  gate1293(.a(s_107), .O(gate86inter4));
  nand2 gate1294(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1295(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1296(.a(G8), .O(gate86inter7));
  inv1  gate1297(.a(G332), .O(gate86inter8));
  nand2 gate1298(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1299(.a(s_107), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1300(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1301(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1302(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1177(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1178(.a(gate87inter0), .b(s_90), .O(gate87inter1));
  and2  gate1179(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1180(.a(s_90), .O(gate87inter3));
  inv1  gate1181(.a(s_91), .O(gate87inter4));
  nand2 gate1182(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1183(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1184(.a(G12), .O(gate87inter7));
  inv1  gate1185(.a(G335), .O(gate87inter8));
  nand2 gate1186(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1187(.a(s_91), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1188(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1189(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1190(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2297(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2298(.a(gate95inter0), .b(s_250), .O(gate95inter1));
  and2  gate2299(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2300(.a(s_250), .O(gate95inter3));
  inv1  gate2301(.a(s_251), .O(gate95inter4));
  nand2 gate2302(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2303(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2304(.a(G26), .O(gate95inter7));
  inv1  gate2305(.a(G347), .O(gate95inter8));
  nand2 gate2306(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2307(.a(s_251), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2308(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2309(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2310(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1205(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1206(.a(gate98inter0), .b(s_94), .O(gate98inter1));
  and2  gate1207(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1208(.a(s_94), .O(gate98inter3));
  inv1  gate1209(.a(s_95), .O(gate98inter4));
  nand2 gate1210(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1211(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1212(.a(G23), .O(gate98inter7));
  inv1  gate1213(.a(G350), .O(gate98inter8));
  nand2 gate1214(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1215(.a(s_95), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1216(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1217(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1218(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2367(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2368(.a(gate100inter0), .b(s_260), .O(gate100inter1));
  and2  gate2369(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2370(.a(s_260), .O(gate100inter3));
  inv1  gate2371(.a(s_261), .O(gate100inter4));
  nand2 gate2372(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2373(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2374(.a(G31), .O(gate100inter7));
  inv1  gate2375(.a(G353), .O(gate100inter8));
  nand2 gate2376(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2377(.a(s_261), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2378(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2379(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2380(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1681(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1682(.a(gate102inter0), .b(s_162), .O(gate102inter1));
  and2  gate1683(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1684(.a(s_162), .O(gate102inter3));
  inv1  gate1685(.a(s_163), .O(gate102inter4));
  nand2 gate1686(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1687(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1688(.a(G24), .O(gate102inter7));
  inv1  gate1689(.a(G356), .O(gate102inter8));
  nand2 gate1690(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1691(.a(s_163), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1692(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1693(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1694(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2129(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2130(.a(gate107inter0), .b(s_226), .O(gate107inter1));
  and2  gate2131(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2132(.a(s_226), .O(gate107inter3));
  inv1  gate2133(.a(s_227), .O(gate107inter4));
  nand2 gate2134(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2135(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2136(.a(G366), .O(gate107inter7));
  inv1  gate2137(.a(G367), .O(gate107inter8));
  nand2 gate2138(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2139(.a(s_227), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2140(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2141(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2142(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2437(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2438(.a(gate110inter0), .b(s_270), .O(gate110inter1));
  and2  gate2439(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2440(.a(s_270), .O(gate110inter3));
  inv1  gate2441(.a(s_271), .O(gate110inter4));
  nand2 gate2442(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2443(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2444(.a(G372), .O(gate110inter7));
  inv1  gate2445(.a(G373), .O(gate110inter8));
  nand2 gate2446(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2447(.a(s_271), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2448(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2449(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2450(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1233(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1234(.a(gate111inter0), .b(s_98), .O(gate111inter1));
  and2  gate1235(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1236(.a(s_98), .O(gate111inter3));
  inv1  gate1237(.a(s_99), .O(gate111inter4));
  nand2 gate1238(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1239(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1240(.a(G374), .O(gate111inter7));
  inv1  gate1241(.a(G375), .O(gate111inter8));
  nand2 gate1242(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1243(.a(s_99), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1244(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1245(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1246(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate827(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate828(.a(gate121inter0), .b(s_40), .O(gate121inter1));
  and2  gate829(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate830(.a(s_40), .O(gate121inter3));
  inv1  gate831(.a(s_41), .O(gate121inter4));
  nand2 gate832(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate833(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate834(.a(G394), .O(gate121inter7));
  inv1  gate835(.a(G395), .O(gate121inter8));
  nand2 gate836(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate837(.a(s_41), .b(gate121inter3), .O(gate121inter10));
  nor2  gate838(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate839(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate840(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1569(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1570(.a(gate123inter0), .b(s_146), .O(gate123inter1));
  and2  gate1571(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1572(.a(s_146), .O(gate123inter3));
  inv1  gate1573(.a(s_147), .O(gate123inter4));
  nand2 gate1574(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1575(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1576(.a(G398), .O(gate123inter7));
  inv1  gate1577(.a(G399), .O(gate123inter8));
  nand2 gate1578(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1579(.a(s_147), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1580(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1581(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1582(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1373(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1374(.a(gate124inter0), .b(s_118), .O(gate124inter1));
  and2  gate1375(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1376(.a(s_118), .O(gate124inter3));
  inv1  gate1377(.a(s_119), .O(gate124inter4));
  nand2 gate1378(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1379(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1380(.a(G400), .O(gate124inter7));
  inv1  gate1381(.a(G401), .O(gate124inter8));
  nand2 gate1382(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1383(.a(s_119), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1384(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1385(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1386(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate2171(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2172(.a(gate125inter0), .b(s_232), .O(gate125inter1));
  and2  gate2173(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2174(.a(s_232), .O(gate125inter3));
  inv1  gate2175(.a(s_233), .O(gate125inter4));
  nand2 gate2176(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2177(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2178(.a(G402), .O(gate125inter7));
  inv1  gate2179(.a(G403), .O(gate125inter8));
  nand2 gate2180(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2181(.a(s_233), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2182(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2183(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2184(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2255(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2256(.a(gate128inter0), .b(s_244), .O(gate128inter1));
  and2  gate2257(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2258(.a(s_244), .O(gate128inter3));
  inv1  gate2259(.a(s_245), .O(gate128inter4));
  nand2 gate2260(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2261(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2262(.a(G408), .O(gate128inter7));
  inv1  gate2263(.a(G409), .O(gate128inter8));
  nand2 gate2264(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2265(.a(s_245), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2266(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2267(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2268(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1359(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1360(.a(gate136inter0), .b(s_116), .O(gate136inter1));
  and2  gate1361(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1362(.a(s_116), .O(gate136inter3));
  inv1  gate1363(.a(s_117), .O(gate136inter4));
  nand2 gate1364(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1365(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1366(.a(G424), .O(gate136inter7));
  inv1  gate1367(.a(G425), .O(gate136inter8));
  nand2 gate1368(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1369(.a(s_117), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1370(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1371(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1372(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1443(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1444(.a(gate146inter0), .b(s_128), .O(gate146inter1));
  and2  gate1445(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1446(.a(s_128), .O(gate146inter3));
  inv1  gate1447(.a(s_129), .O(gate146inter4));
  nand2 gate1448(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1449(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1450(.a(G480), .O(gate146inter7));
  inv1  gate1451(.a(G483), .O(gate146inter8));
  nand2 gate1452(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1453(.a(s_129), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1454(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1455(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1456(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2227(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2228(.a(gate152inter0), .b(s_240), .O(gate152inter1));
  and2  gate2229(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2230(.a(s_240), .O(gate152inter3));
  inv1  gate2231(.a(s_241), .O(gate152inter4));
  nand2 gate2232(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2233(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2234(.a(G516), .O(gate152inter7));
  inv1  gate2235(.a(G519), .O(gate152inter8));
  nand2 gate2236(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2237(.a(s_241), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2238(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2239(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2240(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate1457(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1458(.a(gate153inter0), .b(s_130), .O(gate153inter1));
  and2  gate1459(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1460(.a(s_130), .O(gate153inter3));
  inv1  gate1461(.a(s_131), .O(gate153inter4));
  nand2 gate1462(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1463(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1464(.a(G426), .O(gate153inter7));
  inv1  gate1465(.a(G522), .O(gate153inter8));
  nand2 gate1466(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1467(.a(s_131), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1468(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1469(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1470(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1499(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1500(.a(gate159inter0), .b(s_136), .O(gate159inter1));
  and2  gate1501(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1502(.a(s_136), .O(gate159inter3));
  inv1  gate1503(.a(s_137), .O(gate159inter4));
  nand2 gate1504(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1505(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1506(.a(G444), .O(gate159inter7));
  inv1  gate1507(.a(G531), .O(gate159inter8));
  nand2 gate1508(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1509(.a(s_137), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1510(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1511(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1512(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1093(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1094(.a(gate163inter0), .b(s_78), .O(gate163inter1));
  and2  gate1095(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1096(.a(s_78), .O(gate163inter3));
  inv1  gate1097(.a(s_79), .O(gate163inter4));
  nand2 gate1098(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1099(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1100(.a(G456), .O(gate163inter7));
  inv1  gate1101(.a(G537), .O(gate163inter8));
  nand2 gate1102(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1103(.a(s_79), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1104(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1105(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1106(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate883(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate884(.a(gate167inter0), .b(s_48), .O(gate167inter1));
  and2  gate885(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate886(.a(s_48), .O(gate167inter3));
  inv1  gate887(.a(s_49), .O(gate167inter4));
  nand2 gate888(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate889(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate890(.a(G468), .O(gate167inter7));
  inv1  gate891(.a(G543), .O(gate167inter8));
  nand2 gate892(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate893(.a(s_49), .b(gate167inter3), .O(gate167inter10));
  nor2  gate894(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate895(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate896(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1317(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1318(.a(gate169inter0), .b(s_110), .O(gate169inter1));
  and2  gate1319(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1320(.a(s_110), .O(gate169inter3));
  inv1  gate1321(.a(s_111), .O(gate169inter4));
  nand2 gate1322(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1323(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1324(.a(G474), .O(gate169inter7));
  inv1  gate1325(.a(G546), .O(gate169inter8));
  nand2 gate1326(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1327(.a(s_111), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1328(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1329(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1330(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate659(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate660(.a(gate171inter0), .b(s_16), .O(gate171inter1));
  and2  gate661(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate662(.a(s_16), .O(gate171inter3));
  inv1  gate663(.a(s_17), .O(gate171inter4));
  nand2 gate664(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate665(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate666(.a(G480), .O(gate171inter7));
  inv1  gate667(.a(G549), .O(gate171inter8));
  nand2 gate668(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate669(.a(s_17), .b(gate171inter3), .O(gate171inter10));
  nor2  gate670(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate671(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate672(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2143(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2144(.a(gate172inter0), .b(s_228), .O(gate172inter1));
  and2  gate2145(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2146(.a(s_228), .O(gate172inter3));
  inv1  gate2147(.a(s_229), .O(gate172inter4));
  nand2 gate2148(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2149(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2150(.a(G483), .O(gate172inter7));
  inv1  gate2151(.a(G549), .O(gate172inter8));
  nand2 gate2152(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2153(.a(s_229), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2154(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2155(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2156(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2073(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2074(.a(gate173inter0), .b(s_218), .O(gate173inter1));
  and2  gate2075(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2076(.a(s_218), .O(gate173inter3));
  inv1  gate2077(.a(s_219), .O(gate173inter4));
  nand2 gate2078(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2079(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2080(.a(G486), .O(gate173inter7));
  inv1  gate2081(.a(G552), .O(gate173inter8));
  nand2 gate2082(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2083(.a(s_219), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2084(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2085(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2086(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2031(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2032(.a(gate176inter0), .b(s_212), .O(gate176inter1));
  and2  gate2033(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2034(.a(s_212), .O(gate176inter3));
  inv1  gate2035(.a(s_213), .O(gate176inter4));
  nand2 gate2036(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2037(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2038(.a(G495), .O(gate176inter7));
  inv1  gate2039(.a(G555), .O(gate176inter8));
  nand2 gate2040(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2041(.a(s_213), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2042(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2043(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2044(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate743(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate744(.a(gate178inter0), .b(s_28), .O(gate178inter1));
  and2  gate745(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate746(.a(s_28), .O(gate178inter3));
  inv1  gate747(.a(s_29), .O(gate178inter4));
  nand2 gate748(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate749(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate750(.a(G501), .O(gate178inter7));
  inv1  gate751(.a(G558), .O(gate178inter8));
  nand2 gate752(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate753(.a(s_29), .b(gate178inter3), .O(gate178inter10));
  nor2  gate754(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate755(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate756(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1835(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1836(.a(gate181inter0), .b(s_184), .O(gate181inter1));
  and2  gate1837(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1838(.a(s_184), .O(gate181inter3));
  inv1  gate1839(.a(s_185), .O(gate181inter4));
  nand2 gate1840(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1841(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1842(.a(G510), .O(gate181inter7));
  inv1  gate1843(.a(G564), .O(gate181inter8));
  nand2 gate1844(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1845(.a(s_185), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1846(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1847(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1848(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2269(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2270(.a(gate182inter0), .b(s_246), .O(gate182inter1));
  and2  gate2271(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2272(.a(s_246), .O(gate182inter3));
  inv1  gate2273(.a(s_247), .O(gate182inter4));
  nand2 gate2274(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2275(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2276(.a(G513), .O(gate182inter7));
  inv1  gate2277(.a(G564), .O(gate182inter8));
  nand2 gate2278(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2279(.a(s_247), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2280(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2281(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2282(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate939(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate940(.a(gate183inter0), .b(s_56), .O(gate183inter1));
  and2  gate941(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate942(.a(s_56), .O(gate183inter3));
  inv1  gate943(.a(s_57), .O(gate183inter4));
  nand2 gate944(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate945(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate946(.a(G516), .O(gate183inter7));
  inv1  gate947(.a(G567), .O(gate183inter8));
  nand2 gate948(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate949(.a(s_57), .b(gate183inter3), .O(gate183inter10));
  nor2  gate950(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate951(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate952(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate701(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate702(.a(gate189inter0), .b(s_22), .O(gate189inter1));
  and2  gate703(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate704(.a(s_22), .O(gate189inter3));
  inv1  gate705(.a(s_23), .O(gate189inter4));
  nand2 gate706(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate707(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate708(.a(G578), .O(gate189inter7));
  inv1  gate709(.a(G579), .O(gate189inter8));
  nand2 gate710(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate711(.a(s_23), .b(gate189inter3), .O(gate189inter10));
  nor2  gate712(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate713(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate714(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate855(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate856(.a(gate195inter0), .b(s_44), .O(gate195inter1));
  and2  gate857(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate858(.a(s_44), .O(gate195inter3));
  inv1  gate859(.a(s_45), .O(gate195inter4));
  nand2 gate860(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate861(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate862(.a(G590), .O(gate195inter7));
  inv1  gate863(.a(G591), .O(gate195inter8));
  nand2 gate864(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate865(.a(s_45), .b(gate195inter3), .O(gate195inter10));
  nor2  gate866(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate867(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate868(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate645(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate646(.a(gate197inter0), .b(s_14), .O(gate197inter1));
  and2  gate647(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate648(.a(s_14), .O(gate197inter3));
  inv1  gate649(.a(s_15), .O(gate197inter4));
  nand2 gate650(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate651(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate652(.a(G594), .O(gate197inter7));
  inv1  gate653(.a(G595), .O(gate197inter8));
  nand2 gate654(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate655(.a(s_15), .b(gate197inter3), .O(gate197inter10));
  nor2  gate656(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate657(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate658(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2381(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2382(.a(gate200inter0), .b(s_262), .O(gate200inter1));
  and2  gate2383(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2384(.a(s_262), .O(gate200inter3));
  inv1  gate2385(.a(s_263), .O(gate200inter4));
  nand2 gate2386(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2387(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2388(.a(G600), .O(gate200inter7));
  inv1  gate2389(.a(G601), .O(gate200inter8));
  nand2 gate2390(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2391(.a(s_263), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2392(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2393(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2394(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1583(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1584(.a(gate214inter0), .b(s_148), .O(gate214inter1));
  and2  gate1585(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1586(.a(s_148), .O(gate214inter3));
  inv1  gate1587(.a(s_149), .O(gate214inter4));
  nand2 gate1588(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1589(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1590(.a(G612), .O(gate214inter7));
  inv1  gate1591(.a(G672), .O(gate214inter8));
  nand2 gate1592(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1593(.a(s_149), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1594(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1595(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1596(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1303(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1304(.a(gate216inter0), .b(s_108), .O(gate216inter1));
  and2  gate1305(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1306(.a(s_108), .O(gate216inter3));
  inv1  gate1307(.a(s_109), .O(gate216inter4));
  nand2 gate1308(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1309(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1310(.a(G617), .O(gate216inter7));
  inv1  gate1311(.a(G675), .O(gate216inter8));
  nand2 gate1312(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1313(.a(s_109), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1314(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1315(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1316(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1723(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1724(.a(gate218inter0), .b(s_168), .O(gate218inter1));
  and2  gate1725(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1726(.a(s_168), .O(gate218inter3));
  inv1  gate1727(.a(s_169), .O(gate218inter4));
  nand2 gate1728(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1729(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1730(.a(G627), .O(gate218inter7));
  inv1  gate1731(.a(G678), .O(gate218inter8));
  nand2 gate1732(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1733(.a(s_169), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1734(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1735(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1736(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1611(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1612(.a(gate223inter0), .b(s_152), .O(gate223inter1));
  and2  gate1613(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1614(.a(s_152), .O(gate223inter3));
  inv1  gate1615(.a(s_153), .O(gate223inter4));
  nand2 gate1616(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1617(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1618(.a(G627), .O(gate223inter7));
  inv1  gate1619(.a(G687), .O(gate223inter8));
  nand2 gate1620(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1621(.a(s_153), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1622(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1623(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1624(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1401(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1402(.a(gate224inter0), .b(s_122), .O(gate224inter1));
  and2  gate1403(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1404(.a(s_122), .O(gate224inter3));
  inv1  gate1405(.a(s_123), .O(gate224inter4));
  nand2 gate1406(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1407(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1408(.a(G637), .O(gate224inter7));
  inv1  gate1409(.a(G687), .O(gate224inter8));
  nand2 gate1410(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1411(.a(s_123), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1412(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1413(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1414(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1933(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1934(.a(gate227inter0), .b(s_198), .O(gate227inter1));
  and2  gate1935(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1936(.a(s_198), .O(gate227inter3));
  inv1  gate1937(.a(s_199), .O(gate227inter4));
  nand2 gate1938(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1939(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1940(.a(G694), .O(gate227inter7));
  inv1  gate1941(.a(G695), .O(gate227inter8));
  nand2 gate1942(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1943(.a(s_199), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1944(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1945(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1946(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1261(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1262(.a(gate229inter0), .b(s_102), .O(gate229inter1));
  and2  gate1263(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1264(.a(s_102), .O(gate229inter3));
  inv1  gate1265(.a(s_103), .O(gate229inter4));
  nand2 gate1266(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1267(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1268(.a(G698), .O(gate229inter7));
  inv1  gate1269(.a(G699), .O(gate229inter8));
  nand2 gate1270(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1271(.a(s_103), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1272(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1273(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1274(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate799(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate800(.a(gate231inter0), .b(s_36), .O(gate231inter1));
  and2  gate801(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate802(.a(s_36), .O(gate231inter3));
  inv1  gate803(.a(s_37), .O(gate231inter4));
  nand2 gate804(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate805(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate806(.a(G702), .O(gate231inter7));
  inv1  gate807(.a(G703), .O(gate231inter8));
  nand2 gate808(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate809(.a(s_37), .b(gate231inter3), .O(gate231inter10));
  nor2  gate810(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate811(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate812(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1667(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1668(.a(gate234inter0), .b(s_160), .O(gate234inter1));
  and2  gate1669(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1670(.a(s_160), .O(gate234inter3));
  inv1  gate1671(.a(s_161), .O(gate234inter4));
  nand2 gate1672(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1673(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1674(.a(G245), .O(gate234inter7));
  inv1  gate1675(.a(G721), .O(gate234inter8));
  nand2 gate1676(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1677(.a(s_161), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1678(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1679(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1680(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1429(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1430(.a(gate237inter0), .b(s_126), .O(gate237inter1));
  and2  gate1431(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1432(.a(s_126), .O(gate237inter3));
  inv1  gate1433(.a(s_127), .O(gate237inter4));
  nand2 gate1434(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1435(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1436(.a(G254), .O(gate237inter7));
  inv1  gate1437(.a(G706), .O(gate237inter8));
  nand2 gate1438(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1439(.a(s_127), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1440(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1441(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1442(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1597(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1598(.a(gate238inter0), .b(s_150), .O(gate238inter1));
  and2  gate1599(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1600(.a(s_150), .O(gate238inter3));
  inv1  gate1601(.a(s_151), .O(gate238inter4));
  nand2 gate1602(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1603(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1604(.a(G257), .O(gate238inter7));
  inv1  gate1605(.a(G709), .O(gate238inter8));
  nand2 gate1606(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1607(.a(s_151), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1608(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1609(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1610(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1891(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1892(.a(gate239inter0), .b(s_192), .O(gate239inter1));
  and2  gate1893(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1894(.a(s_192), .O(gate239inter3));
  inv1  gate1895(.a(s_193), .O(gate239inter4));
  nand2 gate1896(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1897(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1898(.a(G260), .O(gate239inter7));
  inv1  gate1899(.a(G712), .O(gate239inter8));
  nand2 gate1900(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1901(.a(s_193), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1902(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1903(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1904(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2353(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2354(.a(gate243inter0), .b(s_258), .O(gate243inter1));
  and2  gate2355(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2356(.a(s_258), .O(gate243inter3));
  inv1  gate2357(.a(s_259), .O(gate243inter4));
  nand2 gate2358(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2359(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2360(.a(G245), .O(gate243inter7));
  inv1  gate2361(.a(G733), .O(gate243inter8));
  nand2 gate2362(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2363(.a(s_259), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2364(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2365(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2366(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1947(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1948(.a(gate253inter0), .b(s_200), .O(gate253inter1));
  and2  gate1949(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1950(.a(s_200), .O(gate253inter3));
  inv1  gate1951(.a(s_201), .O(gate253inter4));
  nand2 gate1952(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1953(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1954(.a(G260), .O(gate253inter7));
  inv1  gate1955(.a(G748), .O(gate253inter8));
  nand2 gate1956(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1957(.a(s_201), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1958(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1959(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1960(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate925(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate926(.a(gate254inter0), .b(s_54), .O(gate254inter1));
  and2  gate927(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate928(.a(s_54), .O(gate254inter3));
  inv1  gate929(.a(s_55), .O(gate254inter4));
  nand2 gate930(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate931(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate932(.a(G712), .O(gate254inter7));
  inv1  gate933(.a(G748), .O(gate254inter8));
  nand2 gate934(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate935(.a(s_55), .b(gate254inter3), .O(gate254inter10));
  nor2  gate936(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate937(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate938(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1653(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1654(.a(gate255inter0), .b(s_158), .O(gate255inter1));
  and2  gate1655(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1656(.a(s_158), .O(gate255inter3));
  inv1  gate1657(.a(s_159), .O(gate255inter4));
  nand2 gate1658(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1659(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1660(.a(G263), .O(gate255inter7));
  inv1  gate1661(.a(G751), .O(gate255inter8));
  nand2 gate1662(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1663(.a(s_159), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1664(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1665(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1666(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1065(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1066(.a(gate260inter0), .b(s_74), .O(gate260inter1));
  and2  gate1067(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1068(.a(s_74), .O(gate260inter3));
  inv1  gate1069(.a(s_75), .O(gate260inter4));
  nand2 gate1070(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1071(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1072(.a(G760), .O(gate260inter7));
  inv1  gate1073(.a(G761), .O(gate260inter8));
  nand2 gate1074(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1075(.a(s_75), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1076(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1077(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1078(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate547(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate548(.a(gate265inter0), .b(s_0), .O(gate265inter1));
  and2  gate549(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate550(.a(s_0), .O(gate265inter3));
  inv1  gate551(.a(s_1), .O(gate265inter4));
  nand2 gate552(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate553(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate554(.a(G642), .O(gate265inter7));
  inv1  gate555(.a(G770), .O(gate265inter8));
  nand2 gate556(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate557(.a(s_1), .b(gate265inter3), .O(gate265inter10));
  nor2  gate558(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate559(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate560(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1807(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1808(.a(gate266inter0), .b(s_180), .O(gate266inter1));
  and2  gate1809(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1810(.a(s_180), .O(gate266inter3));
  inv1  gate1811(.a(s_181), .O(gate266inter4));
  nand2 gate1812(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1813(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1814(.a(G645), .O(gate266inter7));
  inv1  gate1815(.a(G773), .O(gate266inter8));
  nand2 gate1816(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1817(.a(s_181), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1818(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1819(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1820(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate771(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate772(.a(gate267inter0), .b(s_32), .O(gate267inter1));
  and2  gate773(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate774(.a(s_32), .O(gate267inter3));
  inv1  gate775(.a(s_33), .O(gate267inter4));
  nand2 gate776(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate777(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate778(.a(G648), .O(gate267inter7));
  inv1  gate779(.a(G776), .O(gate267inter8));
  nand2 gate780(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate781(.a(s_33), .b(gate267inter3), .O(gate267inter10));
  nor2  gate782(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate783(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate784(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2395(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2396(.a(gate269inter0), .b(s_264), .O(gate269inter1));
  and2  gate2397(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2398(.a(s_264), .O(gate269inter3));
  inv1  gate2399(.a(s_265), .O(gate269inter4));
  nand2 gate2400(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2401(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2402(.a(G654), .O(gate269inter7));
  inv1  gate2403(.a(G782), .O(gate269inter8));
  nand2 gate2404(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2405(.a(s_265), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2406(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2407(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2408(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1275(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1276(.a(gate272inter0), .b(s_104), .O(gate272inter1));
  and2  gate1277(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1278(.a(s_104), .O(gate272inter3));
  inv1  gate1279(.a(s_105), .O(gate272inter4));
  nand2 gate1280(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1281(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1282(.a(G663), .O(gate272inter7));
  inv1  gate1283(.a(G791), .O(gate272inter8));
  nand2 gate1284(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1285(.a(s_105), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1286(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1287(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1288(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1079(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1080(.a(gate274inter0), .b(s_76), .O(gate274inter1));
  and2  gate1081(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1082(.a(s_76), .O(gate274inter3));
  inv1  gate1083(.a(s_77), .O(gate274inter4));
  nand2 gate1084(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1085(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1086(.a(G770), .O(gate274inter7));
  inv1  gate1087(.a(G794), .O(gate274inter8));
  nand2 gate1088(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1089(.a(s_77), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1090(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1091(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1092(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1219(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1220(.a(gate275inter0), .b(s_96), .O(gate275inter1));
  and2  gate1221(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1222(.a(s_96), .O(gate275inter3));
  inv1  gate1223(.a(s_97), .O(gate275inter4));
  nand2 gate1224(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1225(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1226(.a(G645), .O(gate275inter7));
  inv1  gate1227(.a(G797), .O(gate275inter8));
  nand2 gate1228(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1229(.a(s_97), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1230(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1231(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1232(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1541(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1542(.a(gate277inter0), .b(s_142), .O(gate277inter1));
  and2  gate1543(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1544(.a(s_142), .O(gate277inter3));
  inv1  gate1545(.a(s_143), .O(gate277inter4));
  nand2 gate1546(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1547(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1548(.a(G648), .O(gate277inter7));
  inv1  gate1549(.a(G800), .O(gate277inter8));
  nand2 gate1550(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1551(.a(s_143), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1552(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1553(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1554(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate841(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate842(.a(gate278inter0), .b(s_42), .O(gate278inter1));
  and2  gate843(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate844(.a(s_42), .O(gate278inter3));
  inv1  gate845(.a(s_43), .O(gate278inter4));
  nand2 gate846(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate847(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate848(.a(G776), .O(gate278inter7));
  inv1  gate849(.a(G800), .O(gate278inter8));
  nand2 gate850(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate851(.a(s_43), .b(gate278inter3), .O(gate278inter10));
  nor2  gate852(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate853(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate854(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1331(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1332(.a(gate290inter0), .b(s_112), .O(gate290inter1));
  and2  gate1333(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1334(.a(s_112), .O(gate290inter3));
  inv1  gate1335(.a(s_113), .O(gate290inter4));
  nand2 gate1336(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1337(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1338(.a(G820), .O(gate290inter7));
  inv1  gate1339(.a(G821), .O(gate290inter8));
  nand2 gate1340(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1341(.a(s_113), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1342(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1343(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1344(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2003(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2004(.a(gate292inter0), .b(s_208), .O(gate292inter1));
  and2  gate2005(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2006(.a(s_208), .O(gate292inter3));
  inv1  gate2007(.a(s_209), .O(gate292inter4));
  nand2 gate2008(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2009(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2010(.a(G824), .O(gate292inter7));
  inv1  gate2011(.a(G825), .O(gate292inter8));
  nand2 gate2012(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2013(.a(s_209), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2014(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2015(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2016(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2311(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2312(.a(gate294inter0), .b(s_252), .O(gate294inter1));
  and2  gate2313(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2314(.a(s_252), .O(gate294inter3));
  inv1  gate2315(.a(s_253), .O(gate294inter4));
  nand2 gate2316(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2317(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2318(.a(G832), .O(gate294inter7));
  inv1  gate2319(.a(G833), .O(gate294inter8));
  nand2 gate2320(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2321(.a(s_253), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2322(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2323(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2324(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1709(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1710(.a(gate387inter0), .b(s_166), .O(gate387inter1));
  and2  gate1711(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1712(.a(s_166), .O(gate387inter3));
  inv1  gate1713(.a(s_167), .O(gate387inter4));
  nand2 gate1714(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1715(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1716(.a(G1), .O(gate387inter7));
  inv1  gate1717(.a(G1036), .O(gate387inter8));
  nand2 gate1718(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1719(.a(s_167), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1720(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1721(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1722(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2199(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2200(.a(gate393inter0), .b(s_236), .O(gate393inter1));
  and2  gate2201(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2202(.a(s_236), .O(gate393inter3));
  inv1  gate2203(.a(s_237), .O(gate393inter4));
  nand2 gate2204(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2205(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2206(.a(G7), .O(gate393inter7));
  inv1  gate2207(.a(G1054), .O(gate393inter8));
  nand2 gate2208(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2209(.a(s_237), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2210(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2211(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2212(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1765(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1766(.a(gate395inter0), .b(s_174), .O(gate395inter1));
  and2  gate1767(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1768(.a(s_174), .O(gate395inter3));
  inv1  gate1769(.a(s_175), .O(gate395inter4));
  nand2 gate1770(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1771(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1772(.a(G9), .O(gate395inter7));
  inv1  gate1773(.a(G1060), .O(gate395inter8));
  nand2 gate1774(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1775(.a(s_175), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1776(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1777(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1778(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1555(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1556(.a(gate397inter0), .b(s_144), .O(gate397inter1));
  and2  gate1557(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1558(.a(s_144), .O(gate397inter3));
  inv1  gate1559(.a(s_145), .O(gate397inter4));
  nand2 gate1560(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1561(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1562(.a(G11), .O(gate397inter7));
  inv1  gate1563(.a(G1066), .O(gate397inter8));
  nand2 gate1564(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1565(.a(s_145), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1566(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1567(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1568(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1051(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1052(.a(gate398inter0), .b(s_72), .O(gate398inter1));
  and2  gate1053(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1054(.a(s_72), .O(gate398inter3));
  inv1  gate1055(.a(s_73), .O(gate398inter4));
  nand2 gate1056(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1057(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1058(.a(G12), .O(gate398inter7));
  inv1  gate1059(.a(G1069), .O(gate398inter8));
  nand2 gate1060(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1061(.a(s_73), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1062(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1063(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1064(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2087(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2088(.a(gate401inter0), .b(s_220), .O(gate401inter1));
  and2  gate2089(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2090(.a(s_220), .O(gate401inter3));
  inv1  gate2091(.a(s_221), .O(gate401inter4));
  nand2 gate2092(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2093(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2094(.a(G15), .O(gate401inter7));
  inv1  gate2095(.a(G1078), .O(gate401inter8));
  nand2 gate2096(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2097(.a(s_221), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2098(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2099(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2100(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1009(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1010(.a(gate402inter0), .b(s_66), .O(gate402inter1));
  and2  gate1011(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1012(.a(s_66), .O(gate402inter3));
  inv1  gate1013(.a(s_67), .O(gate402inter4));
  nand2 gate1014(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1015(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1016(.a(G16), .O(gate402inter7));
  inv1  gate1017(.a(G1081), .O(gate402inter8));
  nand2 gate1018(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1019(.a(s_67), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1020(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1021(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1022(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1415(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1416(.a(gate403inter0), .b(s_124), .O(gate403inter1));
  and2  gate1417(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1418(.a(s_124), .O(gate403inter3));
  inv1  gate1419(.a(s_125), .O(gate403inter4));
  nand2 gate1420(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1421(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1422(.a(G17), .O(gate403inter7));
  inv1  gate1423(.a(G1084), .O(gate403inter8));
  nand2 gate1424(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1425(.a(s_125), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1426(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1427(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1428(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1849(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1850(.a(gate407inter0), .b(s_186), .O(gate407inter1));
  and2  gate1851(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1852(.a(s_186), .O(gate407inter3));
  inv1  gate1853(.a(s_187), .O(gate407inter4));
  nand2 gate1854(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1855(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1856(.a(G21), .O(gate407inter7));
  inv1  gate1857(.a(G1096), .O(gate407inter8));
  nand2 gate1858(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1859(.a(s_187), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1860(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1861(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1862(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate967(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate968(.a(gate409inter0), .b(s_60), .O(gate409inter1));
  and2  gate969(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate970(.a(s_60), .O(gate409inter3));
  inv1  gate971(.a(s_61), .O(gate409inter4));
  nand2 gate972(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate973(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate974(.a(G23), .O(gate409inter7));
  inv1  gate975(.a(G1102), .O(gate409inter8));
  nand2 gate976(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate977(.a(s_61), .b(gate409inter3), .O(gate409inter10));
  nor2  gate978(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate979(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate980(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2017(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2018(.a(gate415inter0), .b(s_210), .O(gate415inter1));
  and2  gate2019(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2020(.a(s_210), .O(gate415inter3));
  inv1  gate2021(.a(s_211), .O(gate415inter4));
  nand2 gate2022(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2023(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2024(.a(G29), .O(gate415inter7));
  inv1  gate2025(.a(G1120), .O(gate415inter8));
  nand2 gate2026(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2027(.a(s_211), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2028(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2029(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2030(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1163(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1164(.a(gate422inter0), .b(s_88), .O(gate422inter1));
  and2  gate1165(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1166(.a(s_88), .O(gate422inter3));
  inv1  gate1167(.a(s_89), .O(gate422inter4));
  nand2 gate1168(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1169(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1170(.a(G1039), .O(gate422inter7));
  inv1  gate1171(.a(G1135), .O(gate422inter8));
  nand2 gate1172(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1173(.a(s_89), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1174(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1175(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1176(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate2339(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2340(.a(gate423inter0), .b(s_256), .O(gate423inter1));
  and2  gate2341(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2342(.a(s_256), .O(gate423inter3));
  inv1  gate2343(.a(s_257), .O(gate423inter4));
  nand2 gate2344(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2345(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2346(.a(G3), .O(gate423inter7));
  inv1  gate2347(.a(G1138), .O(gate423inter8));
  nand2 gate2348(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2349(.a(s_257), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2350(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2351(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2352(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate687(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate688(.a(gate425inter0), .b(s_20), .O(gate425inter1));
  and2  gate689(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate690(.a(s_20), .O(gate425inter3));
  inv1  gate691(.a(s_21), .O(gate425inter4));
  nand2 gate692(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate693(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate694(.a(G4), .O(gate425inter7));
  inv1  gate695(.a(G1141), .O(gate425inter8));
  nand2 gate696(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate697(.a(s_21), .b(gate425inter3), .O(gate425inter10));
  nor2  gate698(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate699(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate700(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2325(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2326(.a(gate428inter0), .b(s_254), .O(gate428inter1));
  and2  gate2327(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2328(.a(s_254), .O(gate428inter3));
  inv1  gate2329(.a(s_255), .O(gate428inter4));
  nand2 gate2330(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2331(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2332(.a(G1048), .O(gate428inter7));
  inv1  gate2333(.a(G1144), .O(gate428inter8));
  nand2 gate2334(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2335(.a(s_255), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2336(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2337(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2338(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate869(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate870(.a(gate430inter0), .b(s_46), .O(gate430inter1));
  and2  gate871(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate872(.a(s_46), .O(gate430inter3));
  inv1  gate873(.a(s_47), .O(gate430inter4));
  nand2 gate874(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate875(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate876(.a(G1051), .O(gate430inter7));
  inv1  gate877(.a(G1147), .O(gate430inter8));
  nand2 gate878(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate879(.a(s_47), .b(gate430inter3), .O(gate430inter10));
  nor2  gate880(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate881(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate882(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2059(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2060(.a(gate431inter0), .b(s_216), .O(gate431inter1));
  and2  gate2061(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2062(.a(s_216), .O(gate431inter3));
  inv1  gate2063(.a(s_217), .O(gate431inter4));
  nand2 gate2064(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2065(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2066(.a(G7), .O(gate431inter7));
  inv1  gate2067(.a(G1150), .O(gate431inter8));
  nand2 gate2068(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2069(.a(s_217), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2070(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2071(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2072(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate757(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate758(.a(gate434inter0), .b(s_30), .O(gate434inter1));
  and2  gate759(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate760(.a(s_30), .O(gate434inter3));
  inv1  gate761(.a(s_31), .O(gate434inter4));
  nand2 gate762(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate763(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate764(.a(G1057), .O(gate434inter7));
  inv1  gate765(.a(G1153), .O(gate434inter8));
  nand2 gate766(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate767(.a(s_31), .b(gate434inter3), .O(gate434inter10));
  nor2  gate768(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate769(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate770(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2101(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2102(.a(gate438inter0), .b(s_222), .O(gate438inter1));
  and2  gate2103(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2104(.a(s_222), .O(gate438inter3));
  inv1  gate2105(.a(s_223), .O(gate438inter4));
  nand2 gate2106(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2107(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2108(.a(G1063), .O(gate438inter7));
  inv1  gate2109(.a(G1159), .O(gate438inter8));
  nand2 gate2110(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2111(.a(s_223), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2112(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2113(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2114(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2241(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2242(.a(gate444inter0), .b(s_242), .O(gate444inter1));
  and2  gate2243(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2244(.a(s_242), .O(gate444inter3));
  inv1  gate2245(.a(s_243), .O(gate444inter4));
  nand2 gate2246(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2247(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2248(.a(G1072), .O(gate444inter7));
  inv1  gate2249(.a(G1168), .O(gate444inter8));
  nand2 gate2250(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2251(.a(s_243), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2252(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2253(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2254(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1793(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1794(.a(gate447inter0), .b(s_178), .O(gate447inter1));
  and2  gate1795(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1796(.a(s_178), .O(gate447inter3));
  inv1  gate1797(.a(s_179), .O(gate447inter4));
  nand2 gate1798(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1799(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1800(.a(G15), .O(gate447inter7));
  inv1  gate1801(.a(G1174), .O(gate447inter8));
  nand2 gate1802(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1803(.a(s_179), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1804(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1805(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1806(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate561(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate562(.a(gate449inter0), .b(s_2), .O(gate449inter1));
  and2  gate563(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate564(.a(s_2), .O(gate449inter3));
  inv1  gate565(.a(s_3), .O(gate449inter4));
  nand2 gate566(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate567(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate568(.a(G16), .O(gate449inter7));
  inv1  gate569(.a(G1177), .O(gate449inter8));
  nand2 gate570(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate571(.a(s_3), .b(gate449inter3), .O(gate449inter10));
  nor2  gate572(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate573(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate574(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1191(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1192(.a(gate450inter0), .b(s_92), .O(gate450inter1));
  and2  gate1193(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1194(.a(s_92), .O(gate450inter3));
  inv1  gate1195(.a(s_93), .O(gate450inter4));
  nand2 gate1196(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1197(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1198(.a(G1081), .O(gate450inter7));
  inv1  gate1199(.a(G1177), .O(gate450inter8));
  nand2 gate1200(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1201(.a(s_93), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1202(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1203(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1204(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1387(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1388(.a(gate460inter0), .b(s_120), .O(gate460inter1));
  and2  gate1389(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1390(.a(s_120), .O(gate460inter3));
  inv1  gate1391(.a(s_121), .O(gate460inter4));
  nand2 gate1392(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1393(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1394(.a(G1096), .O(gate460inter7));
  inv1  gate1395(.a(G1192), .O(gate460inter8));
  nand2 gate1396(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1397(.a(s_121), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1398(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1399(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1400(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1625(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1626(.a(gate462inter0), .b(s_154), .O(gate462inter1));
  and2  gate1627(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1628(.a(s_154), .O(gate462inter3));
  inv1  gate1629(.a(s_155), .O(gate462inter4));
  nand2 gate1630(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1631(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1632(.a(G1099), .O(gate462inter7));
  inv1  gate1633(.a(G1195), .O(gate462inter8));
  nand2 gate1634(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1635(.a(s_155), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1636(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1637(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1638(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate729(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate730(.a(gate464inter0), .b(s_26), .O(gate464inter1));
  and2  gate731(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate732(.a(s_26), .O(gate464inter3));
  inv1  gate733(.a(s_27), .O(gate464inter4));
  nand2 gate734(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate735(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate736(.a(G1102), .O(gate464inter7));
  inv1  gate737(.a(G1198), .O(gate464inter8));
  nand2 gate738(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate739(.a(s_27), .b(gate464inter3), .O(gate464inter10));
  nor2  gate740(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate741(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate742(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2409(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2410(.a(gate465inter0), .b(s_266), .O(gate465inter1));
  and2  gate2411(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2412(.a(s_266), .O(gate465inter3));
  inv1  gate2413(.a(s_267), .O(gate465inter4));
  nand2 gate2414(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2415(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2416(.a(G24), .O(gate465inter7));
  inv1  gate2417(.a(G1201), .O(gate465inter8));
  nand2 gate2418(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2419(.a(s_267), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2420(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2421(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2422(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate813(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate814(.a(gate466inter0), .b(s_38), .O(gate466inter1));
  and2  gate815(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate816(.a(s_38), .O(gate466inter3));
  inv1  gate817(.a(s_39), .O(gate466inter4));
  nand2 gate818(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate819(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate820(.a(G1105), .O(gate466inter7));
  inv1  gate821(.a(G1201), .O(gate466inter8));
  nand2 gate822(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate823(.a(s_39), .b(gate466inter3), .O(gate466inter10));
  nor2  gate824(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate825(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate826(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1023(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1024(.a(gate473inter0), .b(s_68), .O(gate473inter1));
  and2  gate1025(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1026(.a(s_68), .O(gate473inter3));
  inv1  gate1027(.a(s_69), .O(gate473inter4));
  nand2 gate1028(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1029(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1030(.a(G28), .O(gate473inter7));
  inv1  gate1031(.a(G1213), .O(gate473inter8));
  nand2 gate1032(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1033(.a(s_69), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1034(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1035(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1036(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1135(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1136(.a(gate476inter0), .b(s_84), .O(gate476inter1));
  and2  gate1137(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1138(.a(s_84), .O(gate476inter3));
  inv1  gate1139(.a(s_85), .O(gate476inter4));
  nand2 gate1140(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1141(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1142(.a(G1120), .O(gate476inter7));
  inv1  gate1143(.a(G1216), .O(gate476inter8));
  nand2 gate1144(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1145(.a(s_85), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1146(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1147(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1148(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate631(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate632(.a(gate479inter0), .b(s_12), .O(gate479inter1));
  and2  gate633(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate634(.a(s_12), .O(gate479inter3));
  inv1  gate635(.a(s_13), .O(gate479inter4));
  nand2 gate636(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate637(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate638(.a(G31), .O(gate479inter7));
  inv1  gate639(.a(G1222), .O(gate479inter8));
  nand2 gate640(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate641(.a(s_13), .b(gate479inter3), .O(gate479inter10));
  nor2  gate642(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate643(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate644(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1961(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1962(.a(gate481inter0), .b(s_202), .O(gate481inter1));
  and2  gate1963(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1964(.a(s_202), .O(gate481inter3));
  inv1  gate1965(.a(s_203), .O(gate481inter4));
  nand2 gate1966(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1967(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1968(.a(G32), .O(gate481inter7));
  inv1  gate1969(.a(G1225), .O(gate481inter8));
  nand2 gate1970(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1971(.a(s_203), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1972(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1973(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1974(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1919(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1920(.a(gate482inter0), .b(s_196), .O(gate482inter1));
  and2  gate1921(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1922(.a(s_196), .O(gate482inter3));
  inv1  gate1923(.a(s_197), .O(gate482inter4));
  nand2 gate1924(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1925(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1926(.a(G1129), .O(gate482inter7));
  inv1  gate1927(.a(G1225), .O(gate482inter8));
  nand2 gate1928(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1929(.a(s_197), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1930(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1931(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1932(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1485(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1486(.a(gate483inter0), .b(s_134), .O(gate483inter1));
  and2  gate1487(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1488(.a(s_134), .O(gate483inter3));
  inv1  gate1489(.a(s_135), .O(gate483inter4));
  nand2 gate1490(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1491(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1492(.a(G1228), .O(gate483inter7));
  inv1  gate1493(.a(G1229), .O(gate483inter8));
  nand2 gate1494(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1495(.a(s_135), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1496(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1497(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1498(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1751(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1752(.a(gate484inter0), .b(s_172), .O(gate484inter1));
  and2  gate1753(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1754(.a(s_172), .O(gate484inter3));
  inv1  gate1755(.a(s_173), .O(gate484inter4));
  nand2 gate1756(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1757(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1758(.a(G1230), .O(gate484inter7));
  inv1  gate1759(.a(G1231), .O(gate484inter8));
  nand2 gate1760(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1761(.a(s_173), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1762(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1763(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1764(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1345(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1346(.a(gate486inter0), .b(s_114), .O(gate486inter1));
  and2  gate1347(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1348(.a(s_114), .O(gate486inter3));
  inv1  gate1349(.a(s_115), .O(gate486inter4));
  nand2 gate1350(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1351(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1352(.a(G1234), .O(gate486inter7));
  inv1  gate1353(.a(G1235), .O(gate486inter8));
  nand2 gate1354(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1355(.a(s_115), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1356(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1357(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1358(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2283(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2284(.a(gate493inter0), .b(s_248), .O(gate493inter1));
  and2  gate2285(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2286(.a(s_248), .O(gate493inter3));
  inv1  gate2287(.a(s_249), .O(gate493inter4));
  nand2 gate2288(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2289(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2290(.a(G1248), .O(gate493inter7));
  inv1  gate2291(.a(G1249), .O(gate493inter8));
  nand2 gate2292(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2293(.a(s_249), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2294(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2295(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2296(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate995(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate996(.a(gate495inter0), .b(s_64), .O(gate495inter1));
  and2  gate997(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate998(.a(s_64), .O(gate495inter3));
  inv1  gate999(.a(s_65), .O(gate495inter4));
  nand2 gate1000(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1001(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1002(.a(G1252), .O(gate495inter7));
  inv1  gate1003(.a(G1253), .O(gate495inter8));
  nand2 gate1004(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1005(.a(s_65), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1006(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1007(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1008(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate575(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate576(.a(gate500inter0), .b(s_4), .O(gate500inter1));
  and2  gate577(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate578(.a(s_4), .O(gate500inter3));
  inv1  gate579(.a(s_5), .O(gate500inter4));
  nand2 gate580(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate581(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate582(.a(G1262), .O(gate500inter7));
  inv1  gate583(.a(G1263), .O(gate500inter8));
  nand2 gate584(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate585(.a(s_5), .b(gate500inter3), .O(gate500inter10));
  nor2  gate586(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate587(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate588(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2185(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2186(.a(gate501inter0), .b(s_234), .O(gate501inter1));
  and2  gate2187(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2188(.a(s_234), .O(gate501inter3));
  inv1  gate2189(.a(s_235), .O(gate501inter4));
  nand2 gate2190(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2191(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2192(.a(G1264), .O(gate501inter7));
  inv1  gate2193(.a(G1265), .O(gate501inter8));
  nand2 gate2194(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2195(.a(s_235), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2196(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2197(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2198(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2423(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2424(.a(gate502inter0), .b(s_268), .O(gate502inter1));
  and2  gate2425(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2426(.a(s_268), .O(gate502inter3));
  inv1  gate2427(.a(s_269), .O(gate502inter4));
  nand2 gate2428(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2429(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2430(.a(G1266), .O(gate502inter7));
  inv1  gate2431(.a(G1267), .O(gate502inter8));
  nand2 gate2432(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2433(.a(s_269), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2434(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2435(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2436(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate603(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate604(.a(gate504inter0), .b(s_8), .O(gate504inter1));
  and2  gate605(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate606(.a(s_8), .O(gate504inter3));
  inv1  gate607(.a(s_9), .O(gate504inter4));
  nand2 gate608(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate609(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate610(.a(G1270), .O(gate504inter7));
  inv1  gate611(.a(G1271), .O(gate504inter8));
  nand2 gate612(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate613(.a(s_9), .b(gate504inter3), .O(gate504inter10));
  nor2  gate614(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate615(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate616(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1037(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1038(.a(gate505inter0), .b(s_70), .O(gate505inter1));
  and2  gate1039(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1040(.a(s_70), .O(gate505inter3));
  inv1  gate1041(.a(s_71), .O(gate505inter4));
  nand2 gate1042(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1043(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1044(.a(G1272), .O(gate505inter7));
  inv1  gate1045(.a(G1273), .O(gate505inter8));
  nand2 gate1046(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1047(.a(s_71), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1048(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1049(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1050(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1989(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1990(.a(gate506inter0), .b(s_206), .O(gate506inter1));
  and2  gate1991(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1992(.a(s_206), .O(gate506inter3));
  inv1  gate1993(.a(s_207), .O(gate506inter4));
  nand2 gate1994(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1995(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1996(.a(G1274), .O(gate506inter7));
  inv1  gate1997(.a(G1275), .O(gate506inter8));
  nand2 gate1998(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1999(.a(s_207), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2000(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2001(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2002(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate953(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate954(.a(gate513inter0), .b(s_58), .O(gate513inter1));
  and2  gate955(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate956(.a(s_58), .O(gate513inter3));
  inv1  gate957(.a(s_59), .O(gate513inter4));
  nand2 gate958(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate959(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate960(.a(G1288), .O(gate513inter7));
  inv1  gate961(.a(G1289), .O(gate513inter8));
  nand2 gate962(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate963(.a(s_59), .b(gate513inter3), .O(gate513inter10));
  nor2  gate964(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate965(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate966(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule