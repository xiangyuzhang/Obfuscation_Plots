module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate547(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate548(.a(gate11inter0), .b(s_0), .O(gate11inter1));
  and2  gate549(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate550(.a(s_0), .O(gate11inter3));
  inv1  gate551(.a(s_1), .O(gate11inter4));
  nand2 gate552(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate553(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate554(.a(G5), .O(gate11inter7));
  inv1  gate555(.a(G6), .O(gate11inter8));
  nand2 gate556(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate557(.a(s_1), .b(gate11inter3), .O(gate11inter10));
  nor2  gate558(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate559(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate560(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate785(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate786(.a(gate17inter0), .b(s_34), .O(gate17inter1));
  and2  gate787(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate788(.a(s_34), .O(gate17inter3));
  inv1  gate789(.a(s_35), .O(gate17inter4));
  nand2 gate790(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate791(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate792(.a(G17), .O(gate17inter7));
  inv1  gate793(.a(G18), .O(gate17inter8));
  nand2 gate794(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate795(.a(s_35), .b(gate17inter3), .O(gate17inter10));
  nor2  gate796(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate797(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate798(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate645(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate646(.a(gate19inter0), .b(s_14), .O(gate19inter1));
  and2  gate647(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate648(.a(s_14), .O(gate19inter3));
  inv1  gate649(.a(s_15), .O(gate19inter4));
  nand2 gate650(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate651(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate652(.a(G21), .O(gate19inter7));
  inv1  gate653(.a(G22), .O(gate19inter8));
  nand2 gate654(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate655(.a(s_15), .b(gate19inter3), .O(gate19inter10));
  nor2  gate656(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate657(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate658(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1387(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1388(.a(gate20inter0), .b(s_120), .O(gate20inter1));
  and2  gate1389(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1390(.a(s_120), .O(gate20inter3));
  inv1  gate1391(.a(s_121), .O(gate20inter4));
  nand2 gate1392(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1393(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1394(.a(G23), .O(gate20inter7));
  inv1  gate1395(.a(G24), .O(gate20inter8));
  nand2 gate1396(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1397(.a(s_121), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1398(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1399(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1400(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate687(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate688(.a(gate33inter0), .b(s_20), .O(gate33inter1));
  and2  gate689(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate690(.a(s_20), .O(gate33inter3));
  inv1  gate691(.a(s_21), .O(gate33inter4));
  nand2 gate692(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate693(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate694(.a(G17), .O(gate33inter7));
  inv1  gate695(.a(G21), .O(gate33inter8));
  nand2 gate696(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate697(.a(s_21), .b(gate33inter3), .O(gate33inter10));
  nor2  gate698(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate699(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate700(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate953(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate954(.a(gate41inter0), .b(s_58), .O(gate41inter1));
  and2  gate955(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate956(.a(s_58), .O(gate41inter3));
  inv1  gate957(.a(s_59), .O(gate41inter4));
  nand2 gate958(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate959(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate960(.a(G1), .O(gate41inter7));
  inv1  gate961(.a(G266), .O(gate41inter8));
  nand2 gate962(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate963(.a(s_59), .b(gate41inter3), .O(gate41inter10));
  nor2  gate964(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate965(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate966(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1499(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1500(.a(gate42inter0), .b(s_136), .O(gate42inter1));
  and2  gate1501(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1502(.a(s_136), .O(gate42inter3));
  inv1  gate1503(.a(s_137), .O(gate42inter4));
  nand2 gate1504(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1505(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1506(.a(G2), .O(gate42inter7));
  inv1  gate1507(.a(G266), .O(gate42inter8));
  nand2 gate1508(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1509(.a(s_137), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1510(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1511(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1512(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate967(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate968(.a(gate47inter0), .b(s_60), .O(gate47inter1));
  and2  gate969(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate970(.a(s_60), .O(gate47inter3));
  inv1  gate971(.a(s_61), .O(gate47inter4));
  nand2 gate972(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate973(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate974(.a(G7), .O(gate47inter7));
  inv1  gate975(.a(G275), .O(gate47inter8));
  nand2 gate976(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate977(.a(s_61), .b(gate47inter3), .O(gate47inter10));
  nor2  gate978(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate979(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate980(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate715(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate716(.a(gate49inter0), .b(s_24), .O(gate49inter1));
  and2  gate717(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate718(.a(s_24), .O(gate49inter3));
  inv1  gate719(.a(s_25), .O(gate49inter4));
  nand2 gate720(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate721(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate722(.a(G9), .O(gate49inter7));
  inv1  gate723(.a(G278), .O(gate49inter8));
  nand2 gate724(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate725(.a(s_25), .b(gate49inter3), .O(gate49inter10));
  nor2  gate726(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate727(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate728(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1107(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1108(.a(gate54inter0), .b(s_80), .O(gate54inter1));
  and2  gate1109(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1110(.a(s_80), .O(gate54inter3));
  inv1  gate1111(.a(s_81), .O(gate54inter4));
  nand2 gate1112(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1113(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1114(.a(G14), .O(gate54inter7));
  inv1  gate1115(.a(G284), .O(gate54inter8));
  nand2 gate1116(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1117(.a(s_81), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1118(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1119(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1120(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1093(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1094(.a(gate56inter0), .b(s_78), .O(gate56inter1));
  and2  gate1095(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1096(.a(s_78), .O(gate56inter3));
  inv1  gate1097(.a(s_79), .O(gate56inter4));
  nand2 gate1098(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1099(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1100(.a(G16), .O(gate56inter7));
  inv1  gate1101(.a(G287), .O(gate56inter8));
  nand2 gate1102(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1103(.a(s_79), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1104(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1105(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1106(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate897(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate898(.a(gate57inter0), .b(s_50), .O(gate57inter1));
  and2  gate899(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate900(.a(s_50), .O(gate57inter3));
  inv1  gate901(.a(s_51), .O(gate57inter4));
  nand2 gate902(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate903(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate904(.a(G17), .O(gate57inter7));
  inv1  gate905(.a(G290), .O(gate57inter8));
  nand2 gate906(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate907(.a(s_51), .b(gate57inter3), .O(gate57inter10));
  nor2  gate908(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate909(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate910(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1443(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1444(.a(gate60inter0), .b(s_128), .O(gate60inter1));
  and2  gate1445(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1446(.a(s_128), .O(gate60inter3));
  inv1  gate1447(.a(s_129), .O(gate60inter4));
  nand2 gate1448(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1449(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1450(.a(G20), .O(gate60inter7));
  inv1  gate1451(.a(G293), .O(gate60inter8));
  nand2 gate1452(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1453(.a(s_129), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1454(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1455(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1456(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1331(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1332(.a(gate75inter0), .b(s_112), .O(gate75inter1));
  and2  gate1333(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1334(.a(s_112), .O(gate75inter3));
  inv1  gate1335(.a(s_113), .O(gate75inter4));
  nand2 gate1336(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1337(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1338(.a(G9), .O(gate75inter7));
  inv1  gate1339(.a(G317), .O(gate75inter8));
  nand2 gate1340(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1341(.a(s_113), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1342(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1343(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1344(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1471(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1472(.a(gate78inter0), .b(s_132), .O(gate78inter1));
  and2  gate1473(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1474(.a(s_132), .O(gate78inter3));
  inv1  gate1475(.a(s_133), .O(gate78inter4));
  nand2 gate1476(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1477(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1478(.a(G6), .O(gate78inter7));
  inv1  gate1479(.a(G320), .O(gate78inter8));
  nand2 gate1480(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1481(.a(s_133), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1482(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1483(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1484(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1527(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1528(.a(gate86inter0), .b(s_140), .O(gate86inter1));
  and2  gate1529(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1530(.a(s_140), .O(gate86inter3));
  inv1  gate1531(.a(s_141), .O(gate86inter4));
  nand2 gate1532(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1533(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1534(.a(G8), .O(gate86inter7));
  inv1  gate1535(.a(G332), .O(gate86inter8));
  nand2 gate1536(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1537(.a(s_141), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1538(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1539(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1540(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1065(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1066(.a(gate87inter0), .b(s_74), .O(gate87inter1));
  and2  gate1067(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1068(.a(s_74), .O(gate87inter3));
  inv1  gate1069(.a(s_75), .O(gate87inter4));
  nand2 gate1070(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1071(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1072(.a(G12), .O(gate87inter7));
  inv1  gate1073(.a(G335), .O(gate87inter8));
  nand2 gate1074(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1075(.a(s_75), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1076(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1077(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1078(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1317(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1318(.a(gate88inter0), .b(s_110), .O(gate88inter1));
  and2  gate1319(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1320(.a(s_110), .O(gate88inter3));
  inv1  gate1321(.a(s_111), .O(gate88inter4));
  nand2 gate1322(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1323(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1324(.a(G16), .O(gate88inter7));
  inv1  gate1325(.a(G335), .O(gate88inter8));
  nand2 gate1326(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1327(.a(s_111), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1328(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1329(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1330(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1205(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1206(.a(gate89inter0), .b(s_94), .O(gate89inter1));
  and2  gate1207(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1208(.a(s_94), .O(gate89inter3));
  inv1  gate1209(.a(s_95), .O(gate89inter4));
  nand2 gate1210(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1211(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1212(.a(G17), .O(gate89inter7));
  inv1  gate1213(.a(G338), .O(gate89inter8));
  nand2 gate1214(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1215(.a(s_95), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1216(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1217(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1218(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1303(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1304(.a(gate92inter0), .b(s_108), .O(gate92inter1));
  and2  gate1305(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1306(.a(s_108), .O(gate92inter3));
  inv1  gate1307(.a(s_109), .O(gate92inter4));
  nand2 gate1308(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1309(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1310(.a(G29), .O(gate92inter7));
  inv1  gate1311(.a(G341), .O(gate92inter8));
  nand2 gate1312(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1313(.a(s_109), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1314(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1315(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1316(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate911(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate912(.a(gate102inter0), .b(s_52), .O(gate102inter1));
  and2  gate913(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate914(.a(s_52), .O(gate102inter3));
  inv1  gate915(.a(s_53), .O(gate102inter4));
  nand2 gate916(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate917(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate918(.a(G24), .O(gate102inter7));
  inv1  gate919(.a(G356), .O(gate102inter8));
  nand2 gate920(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate921(.a(s_53), .b(gate102inter3), .O(gate102inter10));
  nor2  gate922(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate923(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate924(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate771(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate772(.a(gate110inter0), .b(s_32), .O(gate110inter1));
  and2  gate773(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate774(.a(s_32), .O(gate110inter3));
  inv1  gate775(.a(s_33), .O(gate110inter4));
  nand2 gate776(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate777(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate778(.a(G372), .O(gate110inter7));
  inv1  gate779(.a(G373), .O(gate110inter8));
  nand2 gate780(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate781(.a(s_33), .b(gate110inter3), .O(gate110inter10));
  nor2  gate782(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate783(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate784(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate659(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate660(.a(gate112inter0), .b(s_16), .O(gate112inter1));
  and2  gate661(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate662(.a(s_16), .O(gate112inter3));
  inv1  gate663(.a(s_17), .O(gate112inter4));
  nand2 gate664(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate665(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate666(.a(G376), .O(gate112inter7));
  inv1  gate667(.a(G377), .O(gate112inter8));
  nand2 gate668(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate669(.a(s_17), .b(gate112inter3), .O(gate112inter10));
  nor2  gate670(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate671(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate672(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1079(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1080(.a(gate115inter0), .b(s_76), .O(gate115inter1));
  and2  gate1081(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1082(.a(s_76), .O(gate115inter3));
  inv1  gate1083(.a(s_77), .O(gate115inter4));
  nand2 gate1084(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1085(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1086(.a(G382), .O(gate115inter7));
  inv1  gate1087(.a(G383), .O(gate115inter8));
  nand2 gate1088(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1089(.a(s_77), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1090(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1091(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1092(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1261(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1262(.a(gate117inter0), .b(s_102), .O(gate117inter1));
  and2  gate1263(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1264(.a(s_102), .O(gate117inter3));
  inv1  gate1265(.a(s_103), .O(gate117inter4));
  nand2 gate1266(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1267(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1268(.a(G386), .O(gate117inter7));
  inv1  gate1269(.a(G387), .O(gate117inter8));
  nand2 gate1270(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1271(.a(s_103), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1272(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1273(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1274(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1373(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1374(.a(gate120inter0), .b(s_118), .O(gate120inter1));
  and2  gate1375(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1376(.a(s_118), .O(gate120inter3));
  inv1  gate1377(.a(s_119), .O(gate120inter4));
  nand2 gate1378(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1379(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1380(.a(G392), .O(gate120inter7));
  inv1  gate1381(.a(G393), .O(gate120inter8));
  nand2 gate1382(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1383(.a(s_119), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1384(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1385(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1386(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate729(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate730(.a(gate127inter0), .b(s_26), .O(gate127inter1));
  and2  gate731(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate732(.a(s_26), .O(gate127inter3));
  inv1  gate733(.a(s_27), .O(gate127inter4));
  nand2 gate734(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate735(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate736(.a(G406), .O(gate127inter7));
  inv1  gate737(.a(G407), .O(gate127inter8));
  nand2 gate738(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate739(.a(s_27), .b(gate127inter3), .O(gate127inter10));
  nor2  gate740(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate741(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate742(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1555(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1556(.a(gate133inter0), .b(s_144), .O(gate133inter1));
  and2  gate1557(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1558(.a(s_144), .O(gate133inter3));
  inv1  gate1559(.a(s_145), .O(gate133inter4));
  nand2 gate1560(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1561(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1562(.a(G418), .O(gate133inter7));
  inv1  gate1563(.a(G419), .O(gate133inter8));
  nand2 gate1564(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1565(.a(s_145), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1566(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1567(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1568(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1569(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1570(.a(gate155inter0), .b(s_146), .O(gate155inter1));
  and2  gate1571(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1572(.a(s_146), .O(gate155inter3));
  inv1  gate1573(.a(s_147), .O(gate155inter4));
  nand2 gate1574(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1575(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1576(.a(G432), .O(gate155inter7));
  inv1  gate1577(.a(G525), .O(gate155inter8));
  nand2 gate1578(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1579(.a(s_147), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1580(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1581(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1582(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1457(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1458(.a(gate158inter0), .b(s_130), .O(gate158inter1));
  and2  gate1459(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1460(.a(s_130), .O(gate158inter3));
  inv1  gate1461(.a(s_131), .O(gate158inter4));
  nand2 gate1462(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1463(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1464(.a(G441), .O(gate158inter7));
  inv1  gate1465(.a(G528), .O(gate158inter8));
  nand2 gate1466(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1467(.a(s_131), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1468(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1469(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1470(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1121(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1122(.a(gate165inter0), .b(s_82), .O(gate165inter1));
  and2  gate1123(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1124(.a(s_82), .O(gate165inter3));
  inv1  gate1125(.a(s_83), .O(gate165inter4));
  nand2 gate1126(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1127(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1128(.a(G462), .O(gate165inter7));
  inv1  gate1129(.a(G540), .O(gate165inter8));
  nand2 gate1130(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1131(.a(s_83), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1132(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1133(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1134(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate575(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate576(.a(gate166inter0), .b(s_4), .O(gate166inter1));
  and2  gate577(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate578(.a(s_4), .O(gate166inter3));
  inv1  gate579(.a(s_5), .O(gate166inter4));
  nand2 gate580(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate581(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate582(.a(G465), .O(gate166inter7));
  inv1  gate583(.a(G540), .O(gate166inter8));
  nand2 gate584(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate585(.a(s_5), .b(gate166inter3), .O(gate166inter10));
  nor2  gate586(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate587(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate588(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate855(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate856(.a(gate171inter0), .b(s_44), .O(gate171inter1));
  and2  gate857(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate858(.a(s_44), .O(gate171inter3));
  inv1  gate859(.a(s_45), .O(gate171inter4));
  nand2 gate860(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate861(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate862(.a(G480), .O(gate171inter7));
  inv1  gate863(.a(G549), .O(gate171inter8));
  nand2 gate864(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate865(.a(s_45), .b(gate171inter3), .O(gate171inter10));
  nor2  gate866(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate867(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate868(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate981(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate982(.a(gate177inter0), .b(s_62), .O(gate177inter1));
  and2  gate983(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate984(.a(s_62), .O(gate177inter3));
  inv1  gate985(.a(s_63), .O(gate177inter4));
  nand2 gate986(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate987(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate988(.a(G498), .O(gate177inter7));
  inv1  gate989(.a(G558), .O(gate177inter8));
  nand2 gate990(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate991(.a(s_63), .b(gate177inter3), .O(gate177inter10));
  nor2  gate992(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate993(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate994(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1359(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1360(.a(gate178inter0), .b(s_116), .O(gate178inter1));
  and2  gate1361(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1362(.a(s_116), .O(gate178inter3));
  inv1  gate1363(.a(s_117), .O(gate178inter4));
  nand2 gate1364(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1365(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1366(.a(G501), .O(gate178inter7));
  inv1  gate1367(.a(G558), .O(gate178inter8));
  nand2 gate1368(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1369(.a(s_117), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1370(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1371(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1372(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate813(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate814(.a(gate180inter0), .b(s_38), .O(gate180inter1));
  and2  gate815(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate816(.a(s_38), .O(gate180inter3));
  inv1  gate817(.a(s_39), .O(gate180inter4));
  nand2 gate818(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate819(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate820(.a(G507), .O(gate180inter7));
  inv1  gate821(.a(G561), .O(gate180inter8));
  nand2 gate822(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate823(.a(s_39), .b(gate180inter3), .O(gate180inter10));
  nor2  gate824(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate825(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate826(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1485(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1486(.a(gate194inter0), .b(s_134), .O(gate194inter1));
  and2  gate1487(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1488(.a(s_134), .O(gate194inter3));
  inv1  gate1489(.a(s_135), .O(gate194inter4));
  nand2 gate1490(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1491(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1492(.a(G588), .O(gate194inter7));
  inv1  gate1493(.a(G589), .O(gate194inter8));
  nand2 gate1494(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1495(.a(s_135), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1496(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1497(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1498(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1625(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1626(.a(gate195inter0), .b(s_154), .O(gate195inter1));
  and2  gate1627(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1628(.a(s_154), .O(gate195inter3));
  inv1  gate1629(.a(s_155), .O(gate195inter4));
  nand2 gate1630(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1631(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1632(.a(G590), .O(gate195inter7));
  inv1  gate1633(.a(G591), .O(gate195inter8));
  nand2 gate1634(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1635(.a(s_155), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1636(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1637(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1638(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate925(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate926(.a(gate204inter0), .b(s_54), .O(gate204inter1));
  and2  gate927(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate928(.a(s_54), .O(gate204inter3));
  inv1  gate929(.a(s_55), .O(gate204inter4));
  nand2 gate930(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate931(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate932(.a(G607), .O(gate204inter7));
  inv1  gate933(.a(G617), .O(gate204inter8));
  nand2 gate934(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate935(.a(s_55), .b(gate204inter3), .O(gate204inter10));
  nor2  gate936(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate937(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate938(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1037(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1038(.a(gate205inter0), .b(s_70), .O(gate205inter1));
  and2  gate1039(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1040(.a(s_70), .O(gate205inter3));
  inv1  gate1041(.a(s_71), .O(gate205inter4));
  nand2 gate1042(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1043(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1044(.a(G622), .O(gate205inter7));
  inv1  gate1045(.a(G627), .O(gate205inter8));
  nand2 gate1046(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1047(.a(s_71), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1048(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1049(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1050(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1513(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1514(.a(gate206inter0), .b(s_138), .O(gate206inter1));
  and2  gate1515(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1516(.a(s_138), .O(gate206inter3));
  inv1  gate1517(.a(s_139), .O(gate206inter4));
  nand2 gate1518(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1519(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1520(.a(G632), .O(gate206inter7));
  inv1  gate1521(.a(G637), .O(gate206inter8));
  nand2 gate1522(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1523(.a(s_139), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1524(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1525(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1526(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate841(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate842(.a(gate207inter0), .b(s_42), .O(gate207inter1));
  and2  gate843(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate844(.a(s_42), .O(gate207inter3));
  inv1  gate845(.a(s_43), .O(gate207inter4));
  nand2 gate846(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate847(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate848(.a(G622), .O(gate207inter7));
  inv1  gate849(.a(G632), .O(gate207inter8));
  nand2 gate850(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate851(.a(s_43), .b(gate207inter3), .O(gate207inter10));
  nor2  gate852(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate853(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate854(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate743(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate744(.a(gate208inter0), .b(s_28), .O(gate208inter1));
  and2  gate745(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate746(.a(s_28), .O(gate208inter3));
  inv1  gate747(.a(s_29), .O(gate208inter4));
  nand2 gate748(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate749(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate750(.a(G627), .O(gate208inter7));
  inv1  gate751(.a(G637), .O(gate208inter8));
  nand2 gate752(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate753(.a(s_29), .b(gate208inter3), .O(gate208inter10));
  nor2  gate754(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate755(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate756(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1149(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1150(.a(gate209inter0), .b(s_86), .O(gate209inter1));
  and2  gate1151(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1152(.a(s_86), .O(gate209inter3));
  inv1  gate1153(.a(s_87), .O(gate209inter4));
  nand2 gate1154(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1155(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1156(.a(G602), .O(gate209inter7));
  inv1  gate1157(.a(G666), .O(gate209inter8));
  nand2 gate1158(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1159(.a(s_87), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1160(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1161(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1162(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1583(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1584(.a(gate211inter0), .b(s_148), .O(gate211inter1));
  and2  gate1585(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1586(.a(s_148), .O(gate211inter3));
  inv1  gate1587(.a(s_149), .O(gate211inter4));
  nand2 gate1588(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1589(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1590(.a(G612), .O(gate211inter7));
  inv1  gate1591(.a(G669), .O(gate211inter8));
  nand2 gate1592(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1593(.a(s_149), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1594(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1595(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1596(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1597(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1598(.a(gate214inter0), .b(s_150), .O(gate214inter1));
  and2  gate1599(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1600(.a(s_150), .O(gate214inter3));
  inv1  gate1601(.a(s_151), .O(gate214inter4));
  nand2 gate1602(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1603(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1604(.a(G612), .O(gate214inter7));
  inv1  gate1605(.a(G672), .O(gate214inter8));
  nand2 gate1606(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1607(.a(s_151), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1608(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1609(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1610(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1289(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1290(.a(gate220inter0), .b(s_106), .O(gate220inter1));
  and2  gate1291(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1292(.a(s_106), .O(gate220inter3));
  inv1  gate1293(.a(s_107), .O(gate220inter4));
  nand2 gate1294(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1295(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1296(.a(G637), .O(gate220inter7));
  inv1  gate1297(.a(G681), .O(gate220inter8));
  nand2 gate1298(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1299(.a(s_107), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1300(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1301(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1302(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate799(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate800(.a(gate224inter0), .b(s_36), .O(gate224inter1));
  and2  gate801(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate802(.a(s_36), .O(gate224inter3));
  inv1  gate803(.a(s_37), .O(gate224inter4));
  nand2 gate804(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate805(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate806(.a(G637), .O(gate224inter7));
  inv1  gate807(.a(G687), .O(gate224inter8));
  nand2 gate808(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate809(.a(s_37), .b(gate224inter3), .O(gate224inter10));
  nor2  gate810(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate811(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate812(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1219(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1220(.a(gate233inter0), .b(s_96), .O(gate233inter1));
  and2  gate1221(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1222(.a(s_96), .O(gate233inter3));
  inv1  gate1223(.a(s_97), .O(gate233inter4));
  nand2 gate1224(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1225(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1226(.a(G242), .O(gate233inter7));
  inv1  gate1227(.a(G718), .O(gate233inter8));
  nand2 gate1228(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1229(.a(s_97), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1230(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1231(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1232(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1163(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1164(.a(gate248inter0), .b(s_88), .O(gate248inter1));
  and2  gate1165(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1166(.a(s_88), .O(gate248inter3));
  inv1  gate1167(.a(s_89), .O(gate248inter4));
  nand2 gate1168(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1169(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1170(.a(G727), .O(gate248inter7));
  inv1  gate1171(.a(G739), .O(gate248inter8));
  nand2 gate1172(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1173(.a(s_89), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1174(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1175(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1176(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1415(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1416(.a(gate253inter0), .b(s_124), .O(gate253inter1));
  and2  gate1417(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1418(.a(s_124), .O(gate253inter3));
  inv1  gate1419(.a(s_125), .O(gate253inter4));
  nand2 gate1420(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1421(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1422(.a(G260), .O(gate253inter7));
  inv1  gate1423(.a(G748), .O(gate253inter8));
  nand2 gate1424(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1425(.a(s_125), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1426(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1427(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1428(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1135(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1136(.a(gate254inter0), .b(s_84), .O(gate254inter1));
  and2  gate1137(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1138(.a(s_84), .O(gate254inter3));
  inv1  gate1139(.a(s_85), .O(gate254inter4));
  nand2 gate1140(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1141(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1142(.a(G712), .O(gate254inter7));
  inv1  gate1143(.a(G748), .O(gate254inter8));
  nand2 gate1144(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1145(.a(s_85), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1146(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1147(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1148(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1611(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1612(.a(gate270inter0), .b(s_152), .O(gate270inter1));
  and2  gate1613(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1614(.a(s_152), .O(gate270inter3));
  inv1  gate1615(.a(s_153), .O(gate270inter4));
  nand2 gate1616(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1617(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1618(.a(G657), .O(gate270inter7));
  inv1  gate1619(.a(G785), .O(gate270inter8));
  nand2 gate1620(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1621(.a(s_153), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1622(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1623(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1624(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate869(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate870(.a(gate280inter0), .b(s_46), .O(gate280inter1));
  and2  gate871(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate872(.a(s_46), .O(gate280inter3));
  inv1  gate873(.a(s_47), .O(gate280inter4));
  nand2 gate874(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate875(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate876(.a(G779), .O(gate280inter7));
  inv1  gate877(.a(G803), .O(gate280inter8));
  nand2 gate878(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate879(.a(s_47), .b(gate280inter3), .O(gate280inter10));
  nor2  gate880(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate881(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate882(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1653(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1654(.a(gate281inter0), .b(s_158), .O(gate281inter1));
  and2  gate1655(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1656(.a(s_158), .O(gate281inter3));
  inv1  gate1657(.a(s_159), .O(gate281inter4));
  nand2 gate1658(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1659(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1660(.a(G654), .O(gate281inter7));
  inv1  gate1661(.a(G806), .O(gate281inter8));
  nand2 gate1662(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1663(.a(s_159), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1664(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1665(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1666(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1191(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1192(.a(gate283inter0), .b(s_92), .O(gate283inter1));
  and2  gate1193(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1194(.a(s_92), .O(gate283inter3));
  inv1  gate1195(.a(s_93), .O(gate283inter4));
  nand2 gate1196(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1197(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1198(.a(G657), .O(gate283inter7));
  inv1  gate1199(.a(G809), .O(gate283inter8));
  nand2 gate1200(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1201(.a(s_93), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1202(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1203(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1204(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate631(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate632(.a(gate285inter0), .b(s_12), .O(gate285inter1));
  and2  gate633(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate634(.a(s_12), .O(gate285inter3));
  inv1  gate635(.a(s_13), .O(gate285inter4));
  nand2 gate636(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate637(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate638(.a(G660), .O(gate285inter7));
  inv1  gate639(.a(G812), .O(gate285inter8));
  nand2 gate640(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate641(.a(s_13), .b(gate285inter3), .O(gate285inter10));
  nor2  gate642(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate643(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate644(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate603(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate604(.a(gate288inter0), .b(s_8), .O(gate288inter1));
  and2  gate605(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate606(.a(s_8), .O(gate288inter3));
  inv1  gate607(.a(s_9), .O(gate288inter4));
  nand2 gate608(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate609(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate610(.a(G791), .O(gate288inter7));
  inv1  gate611(.a(G815), .O(gate288inter8));
  nand2 gate612(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate613(.a(s_9), .b(gate288inter3), .O(gate288inter10));
  nor2  gate614(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate615(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate616(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1009(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1010(.a(gate293inter0), .b(s_66), .O(gate293inter1));
  and2  gate1011(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1012(.a(s_66), .O(gate293inter3));
  inv1  gate1013(.a(s_67), .O(gate293inter4));
  nand2 gate1014(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1015(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1016(.a(G828), .O(gate293inter7));
  inv1  gate1017(.a(G829), .O(gate293inter8));
  nand2 gate1018(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1019(.a(s_67), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1020(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1021(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1022(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1639(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1640(.a(gate294inter0), .b(s_156), .O(gate294inter1));
  and2  gate1641(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1642(.a(s_156), .O(gate294inter3));
  inv1  gate1643(.a(s_157), .O(gate294inter4));
  nand2 gate1644(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1645(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1646(.a(G832), .O(gate294inter7));
  inv1  gate1647(.a(G833), .O(gate294inter8));
  nand2 gate1648(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1649(.a(s_157), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1650(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1651(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1652(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1541(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1542(.a(gate389inter0), .b(s_142), .O(gate389inter1));
  and2  gate1543(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1544(.a(s_142), .O(gate389inter3));
  inv1  gate1545(.a(s_143), .O(gate389inter4));
  nand2 gate1546(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1547(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1548(.a(G3), .O(gate389inter7));
  inv1  gate1549(.a(G1042), .O(gate389inter8));
  nand2 gate1550(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1551(.a(s_143), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1552(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1553(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1554(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1051(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1052(.a(gate391inter0), .b(s_72), .O(gate391inter1));
  and2  gate1053(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1054(.a(s_72), .O(gate391inter3));
  inv1  gate1055(.a(s_73), .O(gate391inter4));
  nand2 gate1056(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1057(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1058(.a(G5), .O(gate391inter7));
  inv1  gate1059(.a(G1048), .O(gate391inter8));
  nand2 gate1060(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1061(.a(s_73), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1062(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1063(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1064(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate701(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate702(.a(gate394inter0), .b(s_22), .O(gate394inter1));
  and2  gate703(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate704(.a(s_22), .O(gate394inter3));
  inv1  gate705(.a(s_23), .O(gate394inter4));
  nand2 gate706(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate707(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate708(.a(G8), .O(gate394inter7));
  inv1  gate709(.a(G1057), .O(gate394inter8));
  nand2 gate710(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate711(.a(s_23), .b(gate394inter3), .O(gate394inter10));
  nor2  gate712(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate713(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate714(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1429(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1430(.a(gate397inter0), .b(s_126), .O(gate397inter1));
  and2  gate1431(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1432(.a(s_126), .O(gate397inter3));
  inv1  gate1433(.a(s_127), .O(gate397inter4));
  nand2 gate1434(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1435(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1436(.a(G11), .O(gate397inter7));
  inv1  gate1437(.a(G1066), .O(gate397inter8));
  nand2 gate1438(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1439(.a(s_127), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1440(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1441(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1442(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate883(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate884(.a(gate405inter0), .b(s_48), .O(gate405inter1));
  and2  gate885(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate886(.a(s_48), .O(gate405inter3));
  inv1  gate887(.a(s_49), .O(gate405inter4));
  nand2 gate888(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate889(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate890(.a(G19), .O(gate405inter7));
  inv1  gate891(.a(G1090), .O(gate405inter8));
  nand2 gate892(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate893(.a(s_49), .b(gate405inter3), .O(gate405inter10));
  nor2  gate894(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate895(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate896(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1401(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1402(.a(gate410inter0), .b(s_122), .O(gate410inter1));
  and2  gate1403(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1404(.a(s_122), .O(gate410inter3));
  inv1  gate1405(.a(s_123), .O(gate410inter4));
  nand2 gate1406(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1407(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1408(.a(G24), .O(gate410inter7));
  inv1  gate1409(.a(G1105), .O(gate410inter8));
  nand2 gate1410(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1411(.a(s_123), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1412(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1413(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1414(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1247(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1248(.a(gate412inter0), .b(s_100), .O(gate412inter1));
  and2  gate1249(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1250(.a(s_100), .O(gate412inter3));
  inv1  gate1251(.a(s_101), .O(gate412inter4));
  nand2 gate1252(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1253(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1254(.a(G26), .O(gate412inter7));
  inv1  gate1255(.a(G1111), .O(gate412inter8));
  nand2 gate1256(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1257(.a(s_101), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1258(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1259(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1260(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1233(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1234(.a(gate417inter0), .b(s_98), .O(gate417inter1));
  and2  gate1235(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1236(.a(s_98), .O(gate417inter3));
  inv1  gate1237(.a(s_99), .O(gate417inter4));
  nand2 gate1238(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1239(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1240(.a(G31), .O(gate417inter7));
  inv1  gate1241(.a(G1126), .O(gate417inter8));
  nand2 gate1242(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1243(.a(s_99), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1244(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1245(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1246(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate995(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate996(.a(gate421inter0), .b(s_64), .O(gate421inter1));
  and2  gate997(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate998(.a(s_64), .O(gate421inter3));
  inv1  gate999(.a(s_65), .O(gate421inter4));
  nand2 gate1000(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1001(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1002(.a(G2), .O(gate421inter7));
  inv1  gate1003(.a(G1135), .O(gate421inter8));
  nand2 gate1004(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1005(.a(s_65), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1006(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1007(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1008(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1275(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1276(.a(gate428inter0), .b(s_104), .O(gate428inter1));
  and2  gate1277(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1278(.a(s_104), .O(gate428inter3));
  inv1  gate1279(.a(s_105), .O(gate428inter4));
  nand2 gate1280(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1281(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1282(.a(G1048), .O(gate428inter7));
  inv1  gate1283(.a(G1144), .O(gate428inter8));
  nand2 gate1284(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1285(.a(s_105), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1286(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1287(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1288(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate939(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate940(.a(gate440inter0), .b(s_56), .O(gate440inter1));
  and2  gate941(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate942(.a(s_56), .O(gate440inter3));
  inv1  gate943(.a(s_57), .O(gate440inter4));
  nand2 gate944(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate945(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate946(.a(G1066), .O(gate440inter7));
  inv1  gate947(.a(G1162), .O(gate440inter8));
  nand2 gate948(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate949(.a(s_57), .b(gate440inter3), .O(gate440inter10));
  nor2  gate950(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate951(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate952(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1177(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1178(.a(gate449inter0), .b(s_90), .O(gate449inter1));
  and2  gate1179(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1180(.a(s_90), .O(gate449inter3));
  inv1  gate1181(.a(s_91), .O(gate449inter4));
  nand2 gate1182(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1183(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1184(.a(G16), .O(gate449inter7));
  inv1  gate1185(.a(G1177), .O(gate449inter8));
  nand2 gate1186(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1187(.a(s_91), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1188(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1189(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1190(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate827(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate828(.a(gate452inter0), .b(s_40), .O(gate452inter1));
  and2  gate829(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate830(.a(s_40), .O(gate452inter3));
  inv1  gate831(.a(s_41), .O(gate452inter4));
  nand2 gate832(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate833(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate834(.a(G1084), .O(gate452inter7));
  inv1  gate835(.a(G1180), .O(gate452inter8));
  nand2 gate836(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate837(.a(s_41), .b(gate452inter3), .O(gate452inter10));
  nor2  gate838(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate839(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate840(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1667(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1668(.a(gate457inter0), .b(s_160), .O(gate457inter1));
  and2  gate1669(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1670(.a(s_160), .O(gate457inter3));
  inv1  gate1671(.a(s_161), .O(gate457inter4));
  nand2 gate1672(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1673(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1674(.a(G20), .O(gate457inter7));
  inv1  gate1675(.a(G1189), .O(gate457inter8));
  nand2 gate1676(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1677(.a(s_161), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1678(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1679(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1680(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate561(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate562(.a(gate466inter0), .b(s_2), .O(gate466inter1));
  and2  gate563(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate564(.a(s_2), .O(gate466inter3));
  inv1  gate565(.a(s_3), .O(gate466inter4));
  nand2 gate566(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate567(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate568(.a(G1105), .O(gate466inter7));
  inv1  gate569(.a(G1201), .O(gate466inter8));
  nand2 gate570(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate571(.a(s_3), .b(gate466inter3), .O(gate466inter10));
  nor2  gate572(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate573(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate574(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate673(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate674(.a(gate482inter0), .b(s_18), .O(gate482inter1));
  and2  gate675(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate676(.a(s_18), .O(gate482inter3));
  inv1  gate677(.a(s_19), .O(gate482inter4));
  nand2 gate678(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate679(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate680(.a(G1129), .O(gate482inter7));
  inv1  gate681(.a(G1225), .O(gate482inter8));
  nand2 gate682(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate683(.a(s_19), .b(gate482inter3), .O(gate482inter10));
  nor2  gate684(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate685(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate686(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate589(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate590(.a(gate492inter0), .b(s_6), .O(gate492inter1));
  and2  gate591(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate592(.a(s_6), .O(gate492inter3));
  inv1  gate593(.a(s_7), .O(gate492inter4));
  nand2 gate594(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate595(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate596(.a(G1246), .O(gate492inter7));
  inv1  gate597(.a(G1247), .O(gate492inter8));
  nand2 gate598(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate599(.a(s_7), .b(gate492inter3), .O(gate492inter10));
  nor2  gate600(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate601(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate602(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1023(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1024(.a(gate501inter0), .b(s_68), .O(gate501inter1));
  and2  gate1025(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1026(.a(s_68), .O(gate501inter3));
  inv1  gate1027(.a(s_69), .O(gate501inter4));
  nand2 gate1028(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1029(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1030(.a(G1264), .O(gate501inter7));
  inv1  gate1031(.a(G1265), .O(gate501inter8));
  nand2 gate1032(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1033(.a(s_69), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1034(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1035(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1036(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate617(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate618(.a(gate502inter0), .b(s_10), .O(gate502inter1));
  and2  gate619(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate620(.a(s_10), .O(gate502inter3));
  inv1  gate621(.a(s_11), .O(gate502inter4));
  nand2 gate622(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate623(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate624(.a(G1266), .O(gate502inter7));
  inv1  gate625(.a(G1267), .O(gate502inter8));
  nand2 gate626(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate627(.a(s_11), .b(gate502inter3), .O(gate502inter10));
  nor2  gate628(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate629(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate630(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate757(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate758(.a(gate504inter0), .b(s_30), .O(gate504inter1));
  and2  gate759(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate760(.a(s_30), .O(gate504inter3));
  inv1  gate761(.a(s_31), .O(gate504inter4));
  nand2 gate762(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate763(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate764(.a(G1270), .O(gate504inter7));
  inv1  gate765(.a(G1271), .O(gate504inter8));
  nand2 gate766(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate767(.a(s_31), .b(gate504inter3), .O(gate504inter10));
  nor2  gate768(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate769(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate770(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1345(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1346(.a(gate508inter0), .b(s_114), .O(gate508inter1));
  and2  gate1347(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1348(.a(s_114), .O(gate508inter3));
  inv1  gate1349(.a(s_115), .O(gate508inter4));
  nand2 gate1350(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1351(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1352(.a(G1278), .O(gate508inter7));
  inv1  gate1353(.a(G1279), .O(gate508inter8));
  nand2 gate1354(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1355(.a(s_115), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1356(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1357(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1358(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule