module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1653(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1654(.a(gate18inter0), .b(s_158), .O(gate18inter1));
  and2  gate1655(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1656(.a(s_158), .O(gate18inter3));
  inv1  gate1657(.a(s_159), .O(gate18inter4));
  nand2 gate1658(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1659(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1660(.a(G19), .O(gate18inter7));
  inv1  gate1661(.a(G20), .O(gate18inter8));
  nand2 gate1662(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1663(.a(s_159), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1664(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1665(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1666(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1079(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1080(.a(gate21inter0), .b(s_76), .O(gate21inter1));
  and2  gate1081(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1082(.a(s_76), .O(gate21inter3));
  inv1  gate1083(.a(s_77), .O(gate21inter4));
  nand2 gate1084(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1085(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1086(.a(G25), .O(gate21inter7));
  inv1  gate1087(.a(G26), .O(gate21inter8));
  nand2 gate1088(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1089(.a(s_77), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1090(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1091(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1092(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1261(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1262(.a(gate33inter0), .b(s_102), .O(gate33inter1));
  and2  gate1263(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1264(.a(s_102), .O(gate33inter3));
  inv1  gate1265(.a(s_103), .O(gate33inter4));
  nand2 gate1266(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1267(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1268(.a(G17), .O(gate33inter7));
  inv1  gate1269(.a(G21), .O(gate33inter8));
  nand2 gate1270(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1271(.a(s_103), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1272(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1273(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1274(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1555(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1556(.a(gate42inter0), .b(s_144), .O(gate42inter1));
  and2  gate1557(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1558(.a(s_144), .O(gate42inter3));
  inv1  gate1559(.a(s_145), .O(gate42inter4));
  nand2 gate1560(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1561(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1562(.a(G2), .O(gate42inter7));
  inv1  gate1563(.a(G266), .O(gate42inter8));
  nand2 gate1564(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1565(.a(s_145), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1566(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1567(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1568(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate799(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate800(.a(gate48inter0), .b(s_36), .O(gate48inter1));
  and2  gate801(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate802(.a(s_36), .O(gate48inter3));
  inv1  gate803(.a(s_37), .O(gate48inter4));
  nand2 gate804(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate805(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate806(.a(G8), .O(gate48inter7));
  inv1  gate807(.a(G275), .O(gate48inter8));
  nand2 gate808(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate809(.a(s_37), .b(gate48inter3), .O(gate48inter10));
  nor2  gate810(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate811(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate812(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1709(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1710(.a(gate54inter0), .b(s_166), .O(gate54inter1));
  and2  gate1711(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1712(.a(s_166), .O(gate54inter3));
  inv1  gate1713(.a(s_167), .O(gate54inter4));
  nand2 gate1714(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1715(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1716(.a(G14), .O(gate54inter7));
  inv1  gate1717(.a(G284), .O(gate54inter8));
  nand2 gate1718(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1719(.a(s_167), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1720(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1721(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1722(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1723(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1724(.a(gate55inter0), .b(s_168), .O(gate55inter1));
  and2  gate1725(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1726(.a(s_168), .O(gate55inter3));
  inv1  gate1727(.a(s_169), .O(gate55inter4));
  nand2 gate1728(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1729(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1730(.a(G15), .O(gate55inter7));
  inv1  gate1731(.a(G287), .O(gate55inter8));
  nand2 gate1732(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1733(.a(s_169), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1734(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1735(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1736(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1443(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1444(.a(gate57inter0), .b(s_128), .O(gate57inter1));
  and2  gate1445(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1446(.a(s_128), .O(gate57inter3));
  inv1  gate1447(.a(s_129), .O(gate57inter4));
  nand2 gate1448(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1449(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1450(.a(G17), .O(gate57inter7));
  inv1  gate1451(.a(G290), .O(gate57inter8));
  nand2 gate1452(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1453(.a(s_129), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1454(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1455(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1456(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1457(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1458(.a(gate63inter0), .b(s_130), .O(gate63inter1));
  and2  gate1459(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1460(.a(s_130), .O(gate63inter3));
  inv1  gate1461(.a(s_131), .O(gate63inter4));
  nand2 gate1462(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1463(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1464(.a(G23), .O(gate63inter7));
  inv1  gate1465(.a(G299), .O(gate63inter8));
  nand2 gate1466(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1467(.a(s_131), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1468(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1469(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1470(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate757(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate758(.a(gate70inter0), .b(s_30), .O(gate70inter1));
  and2  gate759(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate760(.a(s_30), .O(gate70inter3));
  inv1  gate761(.a(s_31), .O(gate70inter4));
  nand2 gate762(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate763(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate764(.a(G30), .O(gate70inter7));
  inv1  gate765(.a(G308), .O(gate70inter8));
  nand2 gate766(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate767(.a(s_31), .b(gate70inter3), .O(gate70inter10));
  nor2  gate768(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate769(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate770(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1401(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1402(.a(gate74inter0), .b(s_122), .O(gate74inter1));
  and2  gate1403(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1404(.a(s_122), .O(gate74inter3));
  inv1  gate1405(.a(s_123), .O(gate74inter4));
  nand2 gate1406(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1407(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1408(.a(G5), .O(gate74inter7));
  inv1  gate1409(.a(G314), .O(gate74inter8));
  nand2 gate1410(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1411(.a(s_123), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1412(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1413(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1414(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1583(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1584(.a(gate78inter0), .b(s_148), .O(gate78inter1));
  and2  gate1585(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1586(.a(s_148), .O(gate78inter3));
  inv1  gate1587(.a(s_149), .O(gate78inter4));
  nand2 gate1588(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1589(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1590(.a(G6), .O(gate78inter7));
  inv1  gate1591(.a(G320), .O(gate78inter8));
  nand2 gate1592(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1593(.a(s_149), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1594(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1595(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1596(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1611(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1612(.a(gate81inter0), .b(s_152), .O(gate81inter1));
  and2  gate1613(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1614(.a(s_152), .O(gate81inter3));
  inv1  gate1615(.a(s_153), .O(gate81inter4));
  nand2 gate1616(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1617(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1618(.a(G3), .O(gate81inter7));
  inv1  gate1619(.a(G326), .O(gate81inter8));
  nand2 gate1620(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1621(.a(s_153), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1622(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1623(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1624(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate939(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate940(.a(gate94inter0), .b(s_56), .O(gate94inter1));
  and2  gate941(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate942(.a(s_56), .O(gate94inter3));
  inv1  gate943(.a(s_57), .O(gate94inter4));
  nand2 gate944(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate945(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate946(.a(G22), .O(gate94inter7));
  inv1  gate947(.a(G344), .O(gate94inter8));
  nand2 gate948(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate949(.a(s_57), .b(gate94inter3), .O(gate94inter10));
  nor2  gate950(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate951(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate952(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate715(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate716(.a(gate97inter0), .b(s_24), .O(gate97inter1));
  and2  gate717(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate718(.a(s_24), .O(gate97inter3));
  inv1  gate719(.a(s_25), .O(gate97inter4));
  nand2 gate720(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate721(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate722(.a(G19), .O(gate97inter7));
  inv1  gate723(.a(G350), .O(gate97inter8));
  nand2 gate724(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate725(.a(s_25), .b(gate97inter3), .O(gate97inter10));
  nor2  gate726(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate727(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate728(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1275(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1276(.a(gate101inter0), .b(s_104), .O(gate101inter1));
  and2  gate1277(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1278(.a(s_104), .O(gate101inter3));
  inv1  gate1279(.a(s_105), .O(gate101inter4));
  nand2 gate1280(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1281(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1282(.a(G20), .O(gate101inter7));
  inv1  gate1283(.a(G356), .O(gate101inter8));
  nand2 gate1284(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1285(.a(s_105), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1286(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1287(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1288(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate855(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate856(.a(gate110inter0), .b(s_44), .O(gate110inter1));
  and2  gate857(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate858(.a(s_44), .O(gate110inter3));
  inv1  gate859(.a(s_45), .O(gate110inter4));
  nand2 gate860(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate861(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate862(.a(G372), .O(gate110inter7));
  inv1  gate863(.a(G373), .O(gate110inter8));
  nand2 gate864(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate865(.a(s_45), .b(gate110inter3), .O(gate110inter10));
  nor2  gate866(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate867(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate868(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1737(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1738(.a(gate116inter0), .b(s_170), .O(gate116inter1));
  and2  gate1739(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1740(.a(s_170), .O(gate116inter3));
  inv1  gate1741(.a(s_171), .O(gate116inter4));
  nand2 gate1742(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1743(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1744(.a(G384), .O(gate116inter7));
  inv1  gate1745(.a(G385), .O(gate116inter8));
  nand2 gate1746(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1747(.a(s_171), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1748(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1749(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1750(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1429(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1430(.a(gate123inter0), .b(s_126), .O(gate123inter1));
  and2  gate1431(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1432(.a(s_126), .O(gate123inter3));
  inv1  gate1433(.a(s_127), .O(gate123inter4));
  nand2 gate1434(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1435(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1436(.a(G398), .O(gate123inter7));
  inv1  gate1437(.a(G399), .O(gate123inter8));
  nand2 gate1438(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1439(.a(s_127), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1440(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1441(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1442(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1485(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1486(.a(gate142inter0), .b(s_134), .O(gate142inter1));
  and2  gate1487(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1488(.a(s_134), .O(gate142inter3));
  inv1  gate1489(.a(s_135), .O(gate142inter4));
  nand2 gate1490(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1491(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1492(.a(G456), .O(gate142inter7));
  inv1  gate1493(.a(G459), .O(gate142inter8));
  nand2 gate1494(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1495(.a(s_135), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1496(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1497(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1498(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1527(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1528(.a(gate143inter0), .b(s_140), .O(gate143inter1));
  and2  gate1529(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1530(.a(s_140), .O(gate143inter3));
  inv1  gate1531(.a(s_141), .O(gate143inter4));
  nand2 gate1532(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1533(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1534(.a(G462), .O(gate143inter7));
  inv1  gate1535(.a(G465), .O(gate143inter8));
  nand2 gate1536(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1537(.a(s_141), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1538(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1539(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1540(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate561(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate562(.a(gate144inter0), .b(s_2), .O(gate144inter1));
  and2  gate563(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate564(.a(s_2), .O(gate144inter3));
  inv1  gate565(.a(s_3), .O(gate144inter4));
  nand2 gate566(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate567(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate568(.a(G468), .O(gate144inter7));
  inv1  gate569(.a(G471), .O(gate144inter8));
  nand2 gate570(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate571(.a(s_3), .b(gate144inter3), .O(gate144inter10));
  nor2  gate572(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate573(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate574(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1051(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1052(.a(gate150inter0), .b(s_72), .O(gate150inter1));
  and2  gate1053(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1054(.a(s_72), .O(gate150inter3));
  inv1  gate1055(.a(s_73), .O(gate150inter4));
  nand2 gate1056(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1057(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1058(.a(G504), .O(gate150inter7));
  inv1  gate1059(.a(G507), .O(gate150inter8));
  nand2 gate1060(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1061(.a(s_73), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1062(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1063(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1064(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate589(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate590(.a(gate152inter0), .b(s_6), .O(gate152inter1));
  and2  gate591(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate592(.a(s_6), .O(gate152inter3));
  inv1  gate593(.a(s_7), .O(gate152inter4));
  nand2 gate594(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate595(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate596(.a(G516), .O(gate152inter7));
  inv1  gate597(.a(G519), .O(gate152inter8));
  nand2 gate598(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate599(.a(s_7), .b(gate152inter3), .O(gate152inter10));
  nor2  gate600(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate601(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate602(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate743(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate744(.a(gate156inter0), .b(s_28), .O(gate156inter1));
  and2  gate745(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate746(.a(s_28), .O(gate156inter3));
  inv1  gate747(.a(s_29), .O(gate156inter4));
  nand2 gate748(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate749(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate750(.a(G435), .O(gate156inter7));
  inv1  gate751(.a(G525), .O(gate156inter8));
  nand2 gate752(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate753(.a(s_29), .b(gate156inter3), .O(gate156inter10));
  nor2  gate754(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate755(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate756(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate841(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate842(.a(gate169inter0), .b(s_42), .O(gate169inter1));
  and2  gate843(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate844(.a(s_42), .O(gate169inter3));
  inv1  gate845(.a(s_43), .O(gate169inter4));
  nand2 gate846(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate847(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate848(.a(G474), .O(gate169inter7));
  inv1  gate849(.a(G546), .O(gate169inter8));
  nand2 gate850(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate851(.a(s_43), .b(gate169inter3), .O(gate169inter10));
  nor2  gate852(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate853(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate854(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1191(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1192(.a(gate170inter0), .b(s_92), .O(gate170inter1));
  and2  gate1193(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1194(.a(s_92), .O(gate170inter3));
  inv1  gate1195(.a(s_93), .O(gate170inter4));
  nand2 gate1196(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1197(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1198(.a(G477), .O(gate170inter7));
  inv1  gate1199(.a(G546), .O(gate170inter8));
  nand2 gate1200(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1201(.a(s_93), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1202(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1203(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1204(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate785(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate786(.a(gate179inter0), .b(s_34), .O(gate179inter1));
  and2  gate787(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate788(.a(s_34), .O(gate179inter3));
  inv1  gate789(.a(s_35), .O(gate179inter4));
  nand2 gate790(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate791(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate792(.a(G504), .O(gate179inter7));
  inv1  gate793(.a(G561), .O(gate179inter8));
  nand2 gate794(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate795(.a(s_35), .b(gate179inter3), .O(gate179inter10));
  nor2  gate796(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate797(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate798(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1345(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1346(.a(gate184inter0), .b(s_114), .O(gate184inter1));
  and2  gate1347(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1348(.a(s_114), .O(gate184inter3));
  inv1  gate1349(.a(s_115), .O(gate184inter4));
  nand2 gate1350(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1351(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1352(.a(G519), .O(gate184inter7));
  inv1  gate1353(.a(G567), .O(gate184inter8));
  nand2 gate1354(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1355(.a(s_115), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1356(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1357(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1358(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate603(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate604(.a(gate185inter0), .b(s_8), .O(gate185inter1));
  and2  gate605(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate606(.a(s_8), .O(gate185inter3));
  inv1  gate607(.a(s_9), .O(gate185inter4));
  nand2 gate608(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate609(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate610(.a(G570), .O(gate185inter7));
  inv1  gate611(.a(G571), .O(gate185inter8));
  nand2 gate612(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate613(.a(s_9), .b(gate185inter3), .O(gate185inter10));
  nor2  gate614(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate615(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate616(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1177(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1178(.a(gate186inter0), .b(s_90), .O(gate186inter1));
  and2  gate1179(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1180(.a(s_90), .O(gate186inter3));
  inv1  gate1181(.a(s_91), .O(gate186inter4));
  nand2 gate1182(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1183(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1184(.a(G572), .O(gate186inter7));
  inv1  gate1185(.a(G573), .O(gate186inter8));
  nand2 gate1186(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1187(.a(s_91), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1188(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1189(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1190(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1023(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1024(.a(gate210inter0), .b(s_68), .O(gate210inter1));
  and2  gate1025(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1026(.a(s_68), .O(gate210inter3));
  inv1  gate1027(.a(s_69), .O(gate210inter4));
  nand2 gate1028(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1029(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1030(.a(G607), .O(gate210inter7));
  inv1  gate1031(.a(G666), .O(gate210inter8));
  nand2 gate1032(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1033(.a(s_69), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1034(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1035(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1036(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1415(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1416(.a(gate214inter0), .b(s_124), .O(gate214inter1));
  and2  gate1417(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1418(.a(s_124), .O(gate214inter3));
  inv1  gate1419(.a(s_125), .O(gate214inter4));
  nand2 gate1420(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1421(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1422(.a(G612), .O(gate214inter7));
  inv1  gate1423(.a(G672), .O(gate214inter8));
  nand2 gate1424(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1425(.a(s_125), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1426(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1427(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1428(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1219(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1220(.a(gate217inter0), .b(s_96), .O(gate217inter1));
  and2  gate1221(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1222(.a(s_96), .O(gate217inter3));
  inv1  gate1223(.a(s_97), .O(gate217inter4));
  nand2 gate1224(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1225(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1226(.a(G622), .O(gate217inter7));
  inv1  gate1227(.a(G678), .O(gate217inter8));
  nand2 gate1228(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1229(.a(s_97), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1230(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1231(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1232(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate813(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate814(.a(gate219inter0), .b(s_38), .O(gate219inter1));
  and2  gate815(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate816(.a(s_38), .O(gate219inter3));
  inv1  gate817(.a(s_39), .O(gate219inter4));
  nand2 gate818(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate819(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate820(.a(G632), .O(gate219inter7));
  inv1  gate821(.a(G681), .O(gate219inter8));
  nand2 gate822(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate823(.a(s_39), .b(gate219inter3), .O(gate219inter10));
  nor2  gate824(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate825(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate826(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate547(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate548(.a(gate221inter0), .b(s_0), .O(gate221inter1));
  and2  gate549(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate550(.a(s_0), .O(gate221inter3));
  inv1  gate551(.a(s_1), .O(gate221inter4));
  nand2 gate552(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate553(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate554(.a(G622), .O(gate221inter7));
  inv1  gate555(.a(G684), .O(gate221inter8));
  nand2 gate556(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate557(.a(s_1), .b(gate221inter3), .O(gate221inter10));
  nor2  gate558(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate559(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate560(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1303(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1304(.a(gate225inter0), .b(s_108), .O(gate225inter1));
  and2  gate1305(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1306(.a(s_108), .O(gate225inter3));
  inv1  gate1307(.a(s_109), .O(gate225inter4));
  nand2 gate1308(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1309(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1310(.a(G690), .O(gate225inter7));
  inv1  gate1311(.a(G691), .O(gate225inter8));
  nand2 gate1312(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1313(.a(s_109), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1314(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1315(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1316(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1639(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1640(.a(gate228inter0), .b(s_156), .O(gate228inter1));
  and2  gate1641(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1642(.a(s_156), .O(gate228inter3));
  inv1  gate1643(.a(s_157), .O(gate228inter4));
  nand2 gate1644(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1645(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1646(.a(G696), .O(gate228inter7));
  inv1  gate1647(.a(G697), .O(gate228inter8));
  nand2 gate1648(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1649(.a(s_157), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1650(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1651(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1652(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate701(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate702(.a(gate229inter0), .b(s_22), .O(gate229inter1));
  and2  gate703(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate704(.a(s_22), .O(gate229inter3));
  inv1  gate705(.a(s_23), .O(gate229inter4));
  nand2 gate706(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate707(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate708(.a(G698), .O(gate229inter7));
  inv1  gate709(.a(G699), .O(gate229inter8));
  nand2 gate710(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate711(.a(s_23), .b(gate229inter3), .O(gate229inter10));
  nor2  gate712(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate713(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate714(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate631(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate632(.a(gate234inter0), .b(s_12), .O(gate234inter1));
  and2  gate633(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate634(.a(s_12), .O(gate234inter3));
  inv1  gate635(.a(s_13), .O(gate234inter4));
  nand2 gate636(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate637(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate638(.a(G245), .O(gate234inter7));
  inv1  gate639(.a(G721), .O(gate234inter8));
  nand2 gate640(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate641(.a(s_13), .b(gate234inter3), .O(gate234inter10));
  nor2  gate642(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate643(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate644(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate659(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate660(.a(gate236inter0), .b(s_16), .O(gate236inter1));
  and2  gate661(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate662(.a(s_16), .O(gate236inter3));
  inv1  gate663(.a(s_17), .O(gate236inter4));
  nand2 gate664(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate665(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate666(.a(G251), .O(gate236inter7));
  inv1  gate667(.a(G727), .O(gate236inter8));
  nand2 gate668(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate669(.a(s_17), .b(gate236inter3), .O(gate236inter10));
  nor2  gate670(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate671(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate672(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate617(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate618(.a(gate248inter0), .b(s_10), .O(gate248inter1));
  and2  gate619(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate620(.a(s_10), .O(gate248inter3));
  inv1  gate621(.a(s_11), .O(gate248inter4));
  nand2 gate622(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate623(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate624(.a(G727), .O(gate248inter7));
  inv1  gate625(.a(G739), .O(gate248inter8));
  nand2 gate626(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate627(.a(s_11), .b(gate248inter3), .O(gate248inter10));
  nor2  gate628(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate629(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate630(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1233(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1234(.a(gate252inter0), .b(s_98), .O(gate252inter1));
  and2  gate1235(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1236(.a(s_98), .O(gate252inter3));
  inv1  gate1237(.a(s_99), .O(gate252inter4));
  nand2 gate1238(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1239(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1240(.a(G709), .O(gate252inter7));
  inv1  gate1241(.a(G745), .O(gate252inter8));
  nand2 gate1242(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1243(.a(s_99), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1244(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1245(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1246(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1107(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1108(.a(gate263inter0), .b(s_80), .O(gate263inter1));
  and2  gate1109(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1110(.a(s_80), .O(gate263inter3));
  inv1  gate1111(.a(s_81), .O(gate263inter4));
  nand2 gate1112(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1113(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1114(.a(G766), .O(gate263inter7));
  inv1  gate1115(.a(G767), .O(gate263inter8));
  nand2 gate1116(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1117(.a(s_81), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1118(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1119(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1120(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate729(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate730(.a(gate269inter0), .b(s_26), .O(gate269inter1));
  and2  gate731(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate732(.a(s_26), .O(gate269inter3));
  inv1  gate733(.a(s_27), .O(gate269inter4));
  nand2 gate734(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate735(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate736(.a(G654), .O(gate269inter7));
  inv1  gate737(.a(G782), .O(gate269inter8));
  nand2 gate738(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate739(.a(s_27), .b(gate269inter3), .O(gate269inter10));
  nor2  gate740(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate741(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate742(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate869(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate870(.a(gate270inter0), .b(s_46), .O(gate270inter1));
  and2  gate871(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate872(.a(s_46), .O(gate270inter3));
  inv1  gate873(.a(s_47), .O(gate270inter4));
  nand2 gate874(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate875(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate876(.a(G657), .O(gate270inter7));
  inv1  gate877(.a(G785), .O(gate270inter8));
  nand2 gate878(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate879(.a(s_47), .b(gate270inter3), .O(gate270inter10));
  nor2  gate880(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate881(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate882(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate771(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate772(.a(gate277inter0), .b(s_32), .O(gate277inter1));
  and2  gate773(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate774(.a(s_32), .O(gate277inter3));
  inv1  gate775(.a(s_33), .O(gate277inter4));
  nand2 gate776(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate777(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate778(.a(G648), .O(gate277inter7));
  inv1  gate779(.a(G800), .O(gate277inter8));
  nand2 gate780(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate781(.a(s_33), .b(gate277inter3), .O(gate277inter10));
  nor2  gate782(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate783(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate784(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate953(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate954(.a(gate278inter0), .b(s_58), .O(gate278inter1));
  and2  gate955(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate956(.a(s_58), .O(gate278inter3));
  inv1  gate957(.a(s_59), .O(gate278inter4));
  nand2 gate958(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate959(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate960(.a(G776), .O(gate278inter7));
  inv1  gate961(.a(G800), .O(gate278inter8));
  nand2 gate962(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate963(.a(s_59), .b(gate278inter3), .O(gate278inter10));
  nor2  gate964(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate965(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate966(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1317(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1318(.a(gate280inter0), .b(s_110), .O(gate280inter1));
  and2  gate1319(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1320(.a(s_110), .O(gate280inter3));
  inv1  gate1321(.a(s_111), .O(gate280inter4));
  nand2 gate1322(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1323(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1324(.a(G779), .O(gate280inter7));
  inv1  gate1325(.a(G803), .O(gate280inter8));
  nand2 gate1326(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1327(.a(s_111), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1328(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1329(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1330(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1373(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1374(.a(gate281inter0), .b(s_118), .O(gate281inter1));
  and2  gate1375(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1376(.a(s_118), .O(gate281inter3));
  inv1  gate1377(.a(s_119), .O(gate281inter4));
  nand2 gate1378(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1379(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1380(.a(G654), .O(gate281inter7));
  inv1  gate1381(.a(G806), .O(gate281inter8));
  nand2 gate1382(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1383(.a(s_119), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1384(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1385(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1386(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1681(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1682(.a(gate282inter0), .b(s_162), .O(gate282inter1));
  and2  gate1683(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1684(.a(s_162), .O(gate282inter3));
  inv1  gate1685(.a(s_163), .O(gate282inter4));
  nand2 gate1686(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1687(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1688(.a(G782), .O(gate282inter7));
  inv1  gate1689(.a(G806), .O(gate282inter8));
  nand2 gate1690(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1691(.a(s_163), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1692(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1693(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1694(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1037(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1038(.a(gate284inter0), .b(s_70), .O(gate284inter1));
  and2  gate1039(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1040(.a(s_70), .O(gate284inter3));
  inv1  gate1041(.a(s_71), .O(gate284inter4));
  nand2 gate1042(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1043(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1044(.a(G785), .O(gate284inter7));
  inv1  gate1045(.a(G809), .O(gate284inter8));
  nand2 gate1046(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1047(.a(s_71), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1048(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1049(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1050(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1513(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1514(.a(gate387inter0), .b(s_138), .O(gate387inter1));
  and2  gate1515(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1516(.a(s_138), .O(gate387inter3));
  inv1  gate1517(.a(s_139), .O(gate387inter4));
  nand2 gate1518(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1519(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1520(.a(G1), .O(gate387inter7));
  inv1  gate1521(.a(G1036), .O(gate387inter8));
  nand2 gate1522(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1523(.a(s_139), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1524(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1525(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1526(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate883(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate884(.a(gate388inter0), .b(s_48), .O(gate388inter1));
  and2  gate885(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate886(.a(s_48), .O(gate388inter3));
  inv1  gate887(.a(s_49), .O(gate388inter4));
  nand2 gate888(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate889(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate890(.a(G2), .O(gate388inter7));
  inv1  gate891(.a(G1039), .O(gate388inter8));
  nand2 gate892(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate893(.a(s_49), .b(gate388inter3), .O(gate388inter10));
  nor2  gate894(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate895(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate896(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1667(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1668(.a(gate389inter0), .b(s_160), .O(gate389inter1));
  and2  gate1669(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1670(.a(s_160), .O(gate389inter3));
  inv1  gate1671(.a(s_161), .O(gate389inter4));
  nand2 gate1672(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1673(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1674(.a(G3), .O(gate389inter7));
  inv1  gate1675(.a(G1042), .O(gate389inter8));
  nand2 gate1676(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1677(.a(s_161), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1678(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1679(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1680(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1541(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1542(.a(gate391inter0), .b(s_142), .O(gate391inter1));
  and2  gate1543(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1544(.a(s_142), .O(gate391inter3));
  inv1  gate1545(.a(s_143), .O(gate391inter4));
  nand2 gate1546(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1547(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1548(.a(G5), .O(gate391inter7));
  inv1  gate1549(.a(G1048), .O(gate391inter8));
  nand2 gate1550(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1551(.a(s_143), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1552(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1553(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1554(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1289(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1290(.a(gate392inter0), .b(s_106), .O(gate392inter1));
  and2  gate1291(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1292(.a(s_106), .O(gate392inter3));
  inv1  gate1293(.a(s_107), .O(gate392inter4));
  nand2 gate1294(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1295(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1296(.a(G6), .O(gate392inter7));
  inv1  gate1297(.a(G1051), .O(gate392inter8));
  nand2 gate1298(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1299(.a(s_107), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1300(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1301(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1302(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1121(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1122(.a(gate401inter0), .b(s_82), .O(gate401inter1));
  and2  gate1123(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1124(.a(s_82), .O(gate401inter3));
  inv1  gate1125(.a(s_83), .O(gate401inter4));
  nand2 gate1126(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1127(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1128(.a(G15), .O(gate401inter7));
  inv1  gate1129(.a(G1078), .O(gate401inter8));
  nand2 gate1130(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1131(.a(s_83), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1132(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1133(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1134(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate645(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate646(.a(gate408inter0), .b(s_14), .O(gate408inter1));
  and2  gate647(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate648(.a(s_14), .O(gate408inter3));
  inv1  gate649(.a(s_15), .O(gate408inter4));
  nand2 gate650(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate651(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate652(.a(G22), .O(gate408inter7));
  inv1  gate653(.a(G1099), .O(gate408inter8));
  nand2 gate654(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate655(.a(s_15), .b(gate408inter3), .O(gate408inter10));
  nor2  gate656(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate657(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate658(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1387(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1388(.a(gate416inter0), .b(s_120), .O(gate416inter1));
  and2  gate1389(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1390(.a(s_120), .O(gate416inter3));
  inv1  gate1391(.a(s_121), .O(gate416inter4));
  nand2 gate1392(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1393(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1394(.a(G30), .O(gate416inter7));
  inv1  gate1395(.a(G1123), .O(gate416inter8));
  nand2 gate1396(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1397(.a(s_121), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1398(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1399(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1400(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1471(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1472(.a(gate422inter0), .b(s_132), .O(gate422inter1));
  and2  gate1473(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1474(.a(s_132), .O(gate422inter3));
  inv1  gate1475(.a(s_133), .O(gate422inter4));
  nand2 gate1476(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1477(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1478(.a(G1039), .O(gate422inter7));
  inv1  gate1479(.a(G1135), .O(gate422inter8));
  nand2 gate1480(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1481(.a(s_133), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1482(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1483(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1484(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1205(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1206(.a(gate425inter0), .b(s_94), .O(gate425inter1));
  and2  gate1207(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1208(.a(s_94), .O(gate425inter3));
  inv1  gate1209(.a(s_95), .O(gate425inter4));
  nand2 gate1210(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1211(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1212(.a(G4), .O(gate425inter7));
  inv1  gate1213(.a(G1141), .O(gate425inter8));
  nand2 gate1214(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1215(.a(s_95), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1216(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1217(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1218(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1163(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1164(.a(gate427inter0), .b(s_88), .O(gate427inter1));
  and2  gate1165(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1166(.a(s_88), .O(gate427inter3));
  inv1  gate1167(.a(s_89), .O(gate427inter4));
  nand2 gate1168(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1169(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1170(.a(G5), .O(gate427inter7));
  inv1  gate1171(.a(G1144), .O(gate427inter8));
  nand2 gate1172(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1173(.a(s_89), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1174(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1175(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1176(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1569(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1570(.a(gate431inter0), .b(s_146), .O(gate431inter1));
  and2  gate1571(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1572(.a(s_146), .O(gate431inter3));
  inv1  gate1573(.a(s_147), .O(gate431inter4));
  nand2 gate1574(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1575(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1576(.a(G7), .O(gate431inter7));
  inv1  gate1577(.a(G1150), .O(gate431inter8));
  nand2 gate1578(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1579(.a(s_147), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1580(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1581(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1582(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate995(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate996(.a(gate432inter0), .b(s_64), .O(gate432inter1));
  and2  gate997(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate998(.a(s_64), .O(gate432inter3));
  inv1  gate999(.a(s_65), .O(gate432inter4));
  nand2 gate1000(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1001(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1002(.a(G1054), .O(gate432inter7));
  inv1  gate1003(.a(G1150), .O(gate432inter8));
  nand2 gate1004(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1005(.a(s_65), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1006(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1007(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1008(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate827(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate828(.a(gate434inter0), .b(s_40), .O(gate434inter1));
  and2  gate829(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate830(.a(s_40), .O(gate434inter3));
  inv1  gate831(.a(s_41), .O(gate434inter4));
  nand2 gate832(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate833(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate834(.a(G1057), .O(gate434inter7));
  inv1  gate835(.a(G1153), .O(gate434inter8));
  nand2 gate836(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate837(.a(s_41), .b(gate434inter3), .O(gate434inter10));
  nor2  gate838(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate839(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate840(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate575(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate576(.a(gate438inter0), .b(s_4), .O(gate438inter1));
  and2  gate577(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate578(.a(s_4), .O(gate438inter3));
  inv1  gate579(.a(s_5), .O(gate438inter4));
  nand2 gate580(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate581(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate582(.a(G1063), .O(gate438inter7));
  inv1  gate583(.a(G1159), .O(gate438inter8));
  nand2 gate584(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate585(.a(s_5), .b(gate438inter3), .O(gate438inter10));
  nor2  gate586(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate587(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate588(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate981(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate982(.a(gate441inter0), .b(s_62), .O(gate441inter1));
  and2  gate983(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate984(.a(s_62), .O(gate441inter3));
  inv1  gate985(.a(s_63), .O(gate441inter4));
  nand2 gate986(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate987(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate988(.a(G12), .O(gate441inter7));
  inv1  gate989(.a(G1165), .O(gate441inter8));
  nand2 gate990(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate991(.a(s_63), .b(gate441inter3), .O(gate441inter10));
  nor2  gate992(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate993(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate994(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1065(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1066(.a(gate442inter0), .b(s_74), .O(gate442inter1));
  and2  gate1067(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1068(.a(s_74), .O(gate442inter3));
  inv1  gate1069(.a(s_75), .O(gate442inter4));
  nand2 gate1070(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1071(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1072(.a(G1069), .O(gate442inter7));
  inv1  gate1073(.a(G1165), .O(gate442inter8));
  nand2 gate1074(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1075(.a(s_75), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1076(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1077(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1078(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate911(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate912(.a(gate444inter0), .b(s_52), .O(gate444inter1));
  and2  gate913(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate914(.a(s_52), .O(gate444inter3));
  inv1  gate915(.a(s_53), .O(gate444inter4));
  nand2 gate916(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate917(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate918(.a(G1072), .O(gate444inter7));
  inv1  gate919(.a(G1168), .O(gate444inter8));
  nand2 gate920(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate921(.a(s_53), .b(gate444inter3), .O(gate444inter10));
  nor2  gate922(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate923(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate924(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate897(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate898(.a(gate447inter0), .b(s_50), .O(gate447inter1));
  and2  gate899(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate900(.a(s_50), .O(gate447inter3));
  inv1  gate901(.a(s_51), .O(gate447inter4));
  nand2 gate902(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate903(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate904(.a(G15), .O(gate447inter7));
  inv1  gate905(.a(G1174), .O(gate447inter8));
  nand2 gate906(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate907(.a(s_51), .b(gate447inter3), .O(gate447inter10));
  nor2  gate908(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate909(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate910(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate687(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate688(.a(gate448inter0), .b(s_20), .O(gate448inter1));
  and2  gate689(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate690(.a(s_20), .O(gate448inter3));
  inv1  gate691(.a(s_21), .O(gate448inter4));
  nand2 gate692(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate693(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate694(.a(G1078), .O(gate448inter7));
  inv1  gate695(.a(G1174), .O(gate448inter8));
  nand2 gate696(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate697(.a(s_21), .b(gate448inter3), .O(gate448inter10));
  nor2  gate698(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate699(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate700(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1359(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1360(.a(gate452inter0), .b(s_116), .O(gate452inter1));
  and2  gate1361(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1362(.a(s_116), .O(gate452inter3));
  inv1  gate1363(.a(s_117), .O(gate452inter4));
  nand2 gate1364(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1365(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1366(.a(G1084), .O(gate452inter7));
  inv1  gate1367(.a(G1180), .O(gate452inter8));
  nand2 gate1368(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1369(.a(s_117), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1370(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1371(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1372(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate673(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate674(.a(gate460inter0), .b(s_18), .O(gate460inter1));
  and2  gate675(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate676(.a(s_18), .O(gate460inter3));
  inv1  gate677(.a(s_19), .O(gate460inter4));
  nand2 gate678(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate679(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate680(.a(G1096), .O(gate460inter7));
  inv1  gate681(.a(G1192), .O(gate460inter8));
  nand2 gate682(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate683(.a(s_19), .b(gate460inter3), .O(gate460inter10));
  nor2  gate684(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate685(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate686(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1499(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1500(.a(gate473inter0), .b(s_136), .O(gate473inter1));
  and2  gate1501(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1502(.a(s_136), .O(gate473inter3));
  inv1  gate1503(.a(s_137), .O(gate473inter4));
  nand2 gate1504(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1505(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1506(.a(G28), .O(gate473inter7));
  inv1  gate1507(.a(G1213), .O(gate473inter8));
  nand2 gate1508(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1509(.a(s_137), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1510(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1511(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1512(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1597(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1598(.a(gate477inter0), .b(s_150), .O(gate477inter1));
  and2  gate1599(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1600(.a(s_150), .O(gate477inter3));
  inv1  gate1601(.a(s_151), .O(gate477inter4));
  nand2 gate1602(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1603(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1604(.a(G30), .O(gate477inter7));
  inv1  gate1605(.a(G1219), .O(gate477inter8));
  nand2 gate1606(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1607(.a(s_151), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1608(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1609(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1610(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1093(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1094(.a(gate481inter0), .b(s_78), .O(gate481inter1));
  and2  gate1095(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1096(.a(s_78), .O(gate481inter3));
  inv1  gate1097(.a(s_79), .O(gate481inter4));
  nand2 gate1098(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1099(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1100(.a(G32), .O(gate481inter7));
  inv1  gate1101(.a(G1225), .O(gate481inter8));
  nand2 gate1102(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1103(.a(s_79), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1104(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1105(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1106(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1135(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1136(.a(gate484inter0), .b(s_84), .O(gate484inter1));
  and2  gate1137(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1138(.a(s_84), .O(gate484inter3));
  inv1  gate1139(.a(s_85), .O(gate484inter4));
  nand2 gate1140(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1141(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1142(.a(G1230), .O(gate484inter7));
  inv1  gate1143(.a(G1231), .O(gate484inter8));
  nand2 gate1144(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1145(.a(s_85), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1146(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1147(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1148(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1331(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1332(.a(gate486inter0), .b(s_112), .O(gate486inter1));
  and2  gate1333(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1334(.a(s_112), .O(gate486inter3));
  inv1  gate1335(.a(s_113), .O(gate486inter4));
  nand2 gate1336(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1337(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1338(.a(G1234), .O(gate486inter7));
  inv1  gate1339(.a(G1235), .O(gate486inter8));
  nand2 gate1340(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1341(.a(s_113), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1342(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1343(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1344(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1149(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1150(.a(gate489inter0), .b(s_86), .O(gate489inter1));
  and2  gate1151(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1152(.a(s_86), .O(gate489inter3));
  inv1  gate1153(.a(s_87), .O(gate489inter4));
  nand2 gate1154(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1155(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1156(.a(G1240), .O(gate489inter7));
  inv1  gate1157(.a(G1241), .O(gate489inter8));
  nand2 gate1158(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1159(.a(s_87), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1160(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1161(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1162(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate925(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate926(.a(gate493inter0), .b(s_54), .O(gate493inter1));
  and2  gate927(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate928(.a(s_54), .O(gate493inter3));
  inv1  gate929(.a(s_55), .O(gate493inter4));
  nand2 gate930(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate931(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate932(.a(G1248), .O(gate493inter7));
  inv1  gate933(.a(G1249), .O(gate493inter8));
  nand2 gate934(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate935(.a(s_55), .b(gate493inter3), .O(gate493inter10));
  nor2  gate936(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate937(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate938(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate967(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate968(.a(gate496inter0), .b(s_60), .O(gate496inter1));
  and2  gate969(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate970(.a(s_60), .O(gate496inter3));
  inv1  gate971(.a(s_61), .O(gate496inter4));
  nand2 gate972(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate973(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate974(.a(G1254), .O(gate496inter7));
  inv1  gate975(.a(G1255), .O(gate496inter8));
  nand2 gate976(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate977(.a(s_61), .b(gate496inter3), .O(gate496inter10));
  nor2  gate978(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate979(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate980(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1009(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1010(.a(gate498inter0), .b(s_66), .O(gate498inter1));
  and2  gate1011(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1012(.a(s_66), .O(gate498inter3));
  inv1  gate1013(.a(s_67), .O(gate498inter4));
  nand2 gate1014(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1015(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1016(.a(G1258), .O(gate498inter7));
  inv1  gate1017(.a(G1259), .O(gate498inter8));
  nand2 gate1018(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1019(.a(s_67), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1020(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1021(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1022(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1625(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1626(.a(gate507inter0), .b(s_154), .O(gate507inter1));
  and2  gate1627(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1628(.a(s_154), .O(gate507inter3));
  inv1  gate1629(.a(s_155), .O(gate507inter4));
  nand2 gate1630(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1631(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1632(.a(G1276), .O(gate507inter7));
  inv1  gate1633(.a(G1277), .O(gate507inter8));
  nand2 gate1634(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1635(.a(s_155), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1636(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1637(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1638(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1247(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1248(.a(gate512inter0), .b(s_100), .O(gate512inter1));
  and2  gate1249(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1250(.a(s_100), .O(gate512inter3));
  inv1  gate1251(.a(s_101), .O(gate512inter4));
  nand2 gate1252(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1253(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1254(.a(G1286), .O(gate512inter7));
  inv1  gate1255(.a(G1287), .O(gate512inter8));
  nand2 gate1256(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1257(.a(s_101), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1258(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1259(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1260(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1695(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1696(.a(gate513inter0), .b(s_164), .O(gate513inter1));
  and2  gate1697(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1698(.a(s_164), .O(gate513inter3));
  inv1  gate1699(.a(s_165), .O(gate513inter4));
  nand2 gate1700(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1701(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1702(.a(G1288), .O(gate513inter7));
  inv1  gate1703(.a(G1289), .O(gate513inter8));
  nand2 gate1704(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1705(.a(s_165), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1706(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1707(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1708(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule