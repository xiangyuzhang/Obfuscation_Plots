module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate659(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate660(.a(gate9inter0), .b(s_16), .O(gate9inter1));
  and2  gate661(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate662(.a(s_16), .O(gate9inter3));
  inv1  gate663(.a(s_17), .O(gate9inter4));
  nand2 gate664(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate665(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate666(.a(G1), .O(gate9inter7));
  inv1  gate667(.a(G2), .O(gate9inter8));
  nand2 gate668(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate669(.a(s_17), .b(gate9inter3), .O(gate9inter10));
  nor2  gate670(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate671(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate672(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1065(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1066(.a(gate12inter0), .b(s_74), .O(gate12inter1));
  and2  gate1067(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1068(.a(s_74), .O(gate12inter3));
  inv1  gate1069(.a(s_75), .O(gate12inter4));
  nand2 gate1070(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1071(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1072(.a(G7), .O(gate12inter7));
  inv1  gate1073(.a(G8), .O(gate12inter8));
  nand2 gate1074(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1075(.a(s_75), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1076(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1077(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1078(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate561(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate562(.a(gate13inter0), .b(s_2), .O(gate13inter1));
  and2  gate563(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate564(.a(s_2), .O(gate13inter3));
  inv1  gate565(.a(s_3), .O(gate13inter4));
  nand2 gate566(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate567(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate568(.a(G9), .O(gate13inter7));
  inv1  gate569(.a(G10), .O(gate13inter8));
  nand2 gate570(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate571(.a(s_3), .b(gate13inter3), .O(gate13inter10));
  nor2  gate572(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate573(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate574(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1093(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1094(.a(gate27inter0), .b(s_78), .O(gate27inter1));
  and2  gate1095(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1096(.a(s_78), .O(gate27inter3));
  inv1  gate1097(.a(s_79), .O(gate27inter4));
  nand2 gate1098(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1099(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1100(.a(G2), .O(gate27inter7));
  inv1  gate1101(.a(G6), .O(gate27inter8));
  nand2 gate1102(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1103(.a(s_79), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1104(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1105(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1106(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate855(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate856(.a(gate39inter0), .b(s_44), .O(gate39inter1));
  and2  gate857(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate858(.a(s_44), .O(gate39inter3));
  inv1  gate859(.a(s_45), .O(gate39inter4));
  nand2 gate860(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate861(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate862(.a(G20), .O(gate39inter7));
  inv1  gate863(.a(G24), .O(gate39inter8));
  nand2 gate864(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate865(.a(s_45), .b(gate39inter3), .O(gate39inter10));
  nor2  gate866(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate867(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate868(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate799(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate800(.a(gate42inter0), .b(s_36), .O(gate42inter1));
  and2  gate801(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate802(.a(s_36), .O(gate42inter3));
  inv1  gate803(.a(s_37), .O(gate42inter4));
  nand2 gate804(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate805(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate806(.a(G2), .O(gate42inter7));
  inv1  gate807(.a(G266), .O(gate42inter8));
  nand2 gate808(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate809(.a(s_37), .b(gate42inter3), .O(gate42inter10));
  nor2  gate810(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate811(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate812(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate729(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate730(.a(gate49inter0), .b(s_26), .O(gate49inter1));
  and2  gate731(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate732(.a(s_26), .O(gate49inter3));
  inv1  gate733(.a(s_27), .O(gate49inter4));
  nand2 gate734(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate735(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate736(.a(G9), .O(gate49inter7));
  inv1  gate737(.a(G278), .O(gate49inter8));
  nand2 gate738(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate739(.a(s_27), .b(gate49inter3), .O(gate49inter10));
  nor2  gate740(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate741(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate742(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1219(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1220(.a(gate52inter0), .b(s_96), .O(gate52inter1));
  and2  gate1221(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1222(.a(s_96), .O(gate52inter3));
  inv1  gate1223(.a(s_97), .O(gate52inter4));
  nand2 gate1224(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1225(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1226(.a(G12), .O(gate52inter7));
  inv1  gate1227(.a(G281), .O(gate52inter8));
  nand2 gate1228(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1229(.a(s_97), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1230(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1231(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1232(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1135(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1136(.a(gate53inter0), .b(s_84), .O(gate53inter1));
  and2  gate1137(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1138(.a(s_84), .O(gate53inter3));
  inv1  gate1139(.a(s_85), .O(gate53inter4));
  nand2 gate1140(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1141(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1142(.a(G13), .O(gate53inter7));
  inv1  gate1143(.a(G284), .O(gate53inter8));
  nand2 gate1144(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1145(.a(s_85), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1146(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1147(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1148(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate771(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate772(.a(gate62inter0), .b(s_32), .O(gate62inter1));
  and2  gate773(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate774(.a(s_32), .O(gate62inter3));
  inv1  gate775(.a(s_33), .O(gate62inter4));
  nand2 gate776(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate777(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate778(.a(G22), .O(gate62inter7));
  inv1  gate779(.a(G296), .O(gate62inter8));
  nand2 gate780(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate781(.a(s_33), .b(gate62inter3), .O(gate62inter10));
  nor2  gate782(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate783(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate784(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate603(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate604(.a(gate66inter0), .b(s_8), .O(gate66inter1));
  and2  gate605(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate606(.a(s_8), .O(gate66inter3));
  inv1  gate607(.a(s_9), .O(gate66inter4));
  nand2 gate608(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate609(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate610(.a(G26), .O(gate66inter7));
  inv1  gate611(.a(G302), .O(gate66inter8));
  nand2 gate612(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate613(.a(s_9), .b(gate66inter3), .O(gate66inter10));
  nor2  gate614(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate615(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate616(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate785(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate786(.a(gate70inter0), .b(s_34), .O(gate70inter1));
  and2  gate787(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate788(.a(s_34), .O(gate70inter3));
  inv1  gate789(.a(s_35), .O(gate70inter4));
  nand2 gate790(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate791(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate792(.a(G30), .O(gate70inter7));
  inv1  gate793(.a(G308), .O(gate70inter8));
  nand2 gate794(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate795(.a(s_35), .b(gate70inter3), .O(gate70inter10));
  nor2  gate796(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate797(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate798(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate897(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate898(.a(gate71inter0), .b(s_50), .O(gate71inter1));
  and2  gate899(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate900(.a(s_50), .O(gate71inter3));
  inv1  gate901(.a(s_51), .O(gate71inter4));
  nand2 gate902(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate903(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate904(.a(G31), .O(gate71inter7));
  inv1  gate905(.a(G311), .O(gate71inter8));
  nand2 gate906(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate907(.a(s_51), .b(gate71inter3), .O(gate71inter10));
  nor2  gate908(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate909(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate910(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate939(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate940(.a(gate76inter0), .b(s_56), .O(gate76inter1));
  and2  gate941(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate942(.a(s_56), .O(gate76inter3));
  inv1  gate943(.a(s_57), .O(gate76inter4));
  nand2 gate944(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate945(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate946(.a(G13), .O(gate76inter7));
  inv1  gate947(.a(G317), .O(gate76inter8));
  nand2 gate948(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate949(.a(s_57), .b(gate76inter3), .O(gate76inter10));
  nor2  gate950(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate951(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate952(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate869(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate870(.a(gate80inter0), .b(s_46), .O(gate80inter1));
  and2  gate871(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate872(.a(s_46), .O(gate80inter3));
  inv1  gate873(.a(s_47), .O(gate80inter4));
  nand2 gate874(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate875(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate876(.a(G14), .O(gate80inter7));
  inv1  gate877(.a(G323), .O(gate80inter8));
  nand2 gate878(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate879(.a(s_47), .b(gate80inter3), .O(gate80inter10));
  nor2  gate880(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate881(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate882(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate617(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate618(.a(gate98inter0), .b(s_10), .O(gate98inter1));
  and2  gate619(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate620(.a(s_10), .O(gate98inter3));
  inv1  gate621(.a(s_11), .O(gate98inter4));
  nand2 gate622(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate623(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate624(.a(G23), .O(gate98inter7));
  inv1  gate625(.a(G350), .O(gate98inter8));
  nand2 gate626(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate627(.a(s_11), .b(gate98inter3), .O(gate98inter10));
  nor2  gate628(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate629(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate630(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate911(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate912(.a(gate108inter0), .b(s_52), .O(gate108inter1));
  and2  gate913(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate914(.a(s_52), .O(gate108inter3));
  inv1  gate915(.a(s_53), .O(gate108inter4));
  nand2 gate916(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate917(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate918(.a(G368), .O(gate108inter7));
  inv1  gate919(.a(G369), .O(gate108inter8));
  nand2 gate920(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate921(.a(s_53), .b(gate108inter3), .O(gate108inter10));
  nor2  gate922(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate923(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate924(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1177(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1178(.a(gate110inter0), .b(s_90), .O(gate110inter1));
  and2  gate1179(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1180(.a(s_90), .O(gate110inter3));
  inv1  gate1181(.a(s_91), .O(gate110inter4));
  nand2 gate1182(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1183(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1184(.a(G372), .O(gate110inter7));
  inv1  gate1185(.a(G373), .O(gate110inter8));
  nand2 gate1186(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1187(.a(s_91), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1188(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1189(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1190(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1121(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1122(.a(gate126inter0), .b(s_82), .O(gate126inter1));
  and2  gate1123(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1124(.a(s_82), .O(gate126inter3));
  inv1  gate1125(.a(s_83), .O(gate126inter4));
  nand2 gate1126(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1127(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1128(.a(G404), .O(gate126inter7));
  inv1  gate1129(.a(G405), .O(gate126inter8));
  nand2 gate1130(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1131(.a(s_83), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1132(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1133(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1134(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1247(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1248(.a(gate135inter0), .b(s_100), .O(gate135inter1));
  and2  gate1249(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1250(.a(s_100), .O(gate135inter3));
  inv1  gate1251(.a(s_101), .O(gate135inter4));
  nand2 gate1252(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1253(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1254(.a(G422), .O(gate135inter7));
  inv1  gate1255(.a(G423), .O(gate135inter8));
  nand2 gate1256(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1257(.a(s_101), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1258(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1259(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1260(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate743(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate744(.a(gate144inter0), .b(s_28), .O(gate144inter1));
  and2  gate745(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate746(.a(s_28), .O(gate144inter3));
  inv1  gate747(.a(s_29), .O(gate144inter4));
  nand2 gate748(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate749(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate750(.a(G468), .O(gate144inter7));
  inv1  gate751(.a(G471), .O(gate144inter8));
  nand2 gate752(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate753(.a(s_29), .b(gate144inter3), .O(gate144inter10));
  nor2  gate754(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate755(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate756(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate981(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate982(.a(gate159inter0), .b(s_62), .O(gate159inter1));
  and2  gate983(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate984(.a(s_62), .O(gate159inter3));
  inv1  gate985(.a(s_63), .O(gate159inter4));
  nand2 gate986(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate987(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate988(.a(G444), .O(gate159inter7));
  inv1  gate989(.a(G531), .O(gate159inter8));
  nand2 gate990(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate991(.a(s_63), .b(gate159inter3), .O(gate159inter10));
  nor2  gate992(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate993(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate994(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1205(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1206(.a(gate160inter0), .b(s_94), .O(gate160inter1));
  and2  gate1207(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1208(.a(s_94), .O(gate160inter3));
  inv1  gate1209(.a(s_95), .O(gate160inter4));
  nand2 gate1210(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1211(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1212(.a(G447), .O(gate160inter7));
  inv1  gate1213(.a(G531), .O(gate160inter8));
  nand2 gate1214(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1215(.a(s_95), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1216(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1217(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1218(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate995(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate996(.a(gate166inter0), .b(s_64), .O(gate166inter1));
  and2  gate997(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate998(.a(s_64), .O(gate166inter3));
  inv1  gate999(.a(s_65), .O(gate166inter4));
  nand2 gate1000(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1001(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1002(.a(G465), .O(gate166inter7));
  inv1  gate1003(.a(G540), .O(gate166inter8));
  nand2 gate1004(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1005(.a(s_65), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1006(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1007(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1008(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1023(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1024(.a(gate173inter0), .b(s_68), .O(gate173inter1));
  and2  gate1025(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1026(.a(s_68), .O(gate173inter3));
  inv1  gate1027(.a(s_69), .O(gate173inter4));
  nand2 gate1028(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1029(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1030(.a(G486), .O(gate173inter7));
  inv1  gate1031(.a(G552), .O(gate173inter8));
  nand2 gate1032(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1033(.a(s_69), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1034(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1035(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1036(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate883(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate884(.a(gate189inter0), .b(s_48), .O(gate189inter1));
  and2  gate885(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate886(.a(s_48), .O(gate189inter3));
  inv1  gate887(.a(s_49), .O(gate189inter4));
  nand2 gate888(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate889(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate890(.a(G578), .O(gate189inter7));
  inv1  gate891(.a(G579), .O(gate189inter8));
  nand2 gate892(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate893(.a(s_49), .b(gate189inter3), .O(gate189inter10));
  nor2  gate894(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate895(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate896(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate687(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate688(.a(gate215inter0), .b(s_20), .O(gate215inter1));
  and2  gate689(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate690(.a(s_20), .O(gate215inter3));
  inv1  gate691(.a(s_21), .O(gate215inter4));
  nand2 gate692(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate693(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate694(.a(G607), .O(gate215inter7));
  inv1  gate695(.a(G675), .O(gate215inter8));
  nand2 gate696(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate697(.a(s_21), .b(gate215inter3), .O(gate215inter10));
  nor2  gate698(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate699(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate700(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1037(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1038(.a(gate221inter0), .b(s_70), .O(gate221inter1));
  and2  gate1039(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1040(.a(s_70), .O(gate221inter3));
  inv1  gate1041(.a(s_71), .O(gate221inter4));
  nand2 gate1042(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1043(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1044(.a(G622), .O(gate221inter7));
  inv1  gate1045(.a(G684), .O(gate221inter8));
  nand2 gate1046(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1047(.a(s_71), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1048(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1049(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1050(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate631(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate632(.a(gate228inter0), .b(s_12), .O(gate228inter1));
  and2  gate633(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate634(.a(s_12), .O(gate228inter3));
  inv1  gate635(.a(s_13), .O(gate228inter4));
  nand2 gate636(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate637(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate638(.a(G696), .O(gate228inter7));
  inv1  gate639(.a(G697), .O(gate228inter8));
  nand2 gate640(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate641(.a(s_13), .b(gate228inter3), .O(gate228inter10));
  nor2  gate642(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate643(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate644(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate589(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate590(.a(gate242inter0), .b(s_6), .O(gate242inter1));
  and2  gate591(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate592(.a(s_6), .O(gate242inter3));
  inv1  gate593(.a(s_7), .O(gate242inter4));
  nand2 gate594(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate595(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate596(.a(G718), .O(gate242inter7));
  inv1  gate597(.a(G730), .O(gate242inter8));
  nand2 gate598(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate599(.a(s_7), .b(gate242inter3), .O(gate242inter10));
  nor2  gate600(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate601(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate602(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate715(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate716(.a(gate255inter0), .b(s_24), .O(gate255inter1));
  and2  gate717(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate718(.a(s_24), .O(gate255inter3));
  inv1  gate719(.a(s_25), .O(gate255inter4));
  nand2 gate720(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate721(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate722(.a(G263), .O(gate255inter7));
  inv1  gate723(.a(G751), .O(gate255inter8));
  nand2 gate724(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate725(.a(s_25), .b(gate255inter3), .O(gate255inter10));
  nor2  gate726(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate727(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate728(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate757(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate758(.a(gate258inter0), .b(s_30), .O(gate258inter1));
  and2  gate759(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate760(.a(s_30), .O(gate258inter3));
  inv1  gate761(.a(s_31), .O(gate258inter4));
  nand2 gate762(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate763(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate764(.a(G756), .O(gate258inter7));
  inv1  gate765(.a(G757), .O(gate258inter8));
  nand2 gate766(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate767(.a(s_31), .b(gate258inter3), .O(gate258inter10));
  nor2  gate768(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate769(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate770(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate645(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate646(.a(gate282inter0), .b(s_14), .O(gate282inter1));
  and2  gate647(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate648(.a(s_14), .O(gate282inter3));
  inv1  gate649(.a(s_15), .O(gate282inter4));
  nand2 gate650(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate651(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate652(.a(G782), .O(gate282inter7));
  inv1  gate653(.a(G806), .O(gate282inter8));
  nand2 gate654(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate655(.a(s_15), .b(gate282inter3), .O(gate282inter10));
  nor2  gate656(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate657(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate658(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate701(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate702(.a(gate286inter0), .b(s_22), .O(gate286inter1));
  and2  gate703(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate704(.a(s_22), .O(gate286inter3));
  inv1  gate705(.a(s_23), .O(gate286inter4));
  nand2 gate706(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate707(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate708(.a(G788), .O(gate286inter7));
  inv1  gate709(.a(G812), .O(gate286inter8));
  nand2 gate710(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate711(.a(s_23), .b(gate286inter3), .O(gate286inter10));
  nor2  gate712(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate713(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate714(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1191(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1192(.a(gate290inter0), .b(s_92), .O(gate290inter1));
  and2  gate1193(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1194(.a(s_92), .O(gate290inter3));
  inv1  gate1195(.a(s_93), .O(gate290inter4));
  nand2 gate1196(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1197(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1198(.a(G820), .O(gate290inter7));
  inv1  gate1199(.a(G821), .O(gate290inter8));
  nand2 gate1200(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1201(.a(s_93), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1202(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1203(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1204(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate953(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate954(.a(gate387inter0), .b(s_58), .O(gate387inter1));
  and2  gate955(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate956(.a(s_58), .O(gate387inter3));
  inv1  gate957(.a(s_59), .O(gate387inter4));
  nand2 gate958(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate959(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate960(.a(G1), .O(gate387inter7));
  inv1  gate961(.a(G1036), .O(gate387inter8));
  nand2 gate962(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate963(.a(s_59), .b(gate387inter3), .O(gate387inter10));
  nor2  gate964(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate965(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate966(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1163(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1164(.a(gate393inter0), .b(s_88), .O(gate393inter1));
  and2  gate1165(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1166(.a(s_88), .O(gate393inter3));
  inv1  gate1167(.a(s_89), .O(gate393inter4));
  nand2 gate1168(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1169(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1170(.a(G7), .O(gate393inter7));
  inv1  gate1171(.a(G1054), .O(gate393inter8));
  nand2 gate1172(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1173(.a(s_89), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1174(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1175(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1176(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate827(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate828(.a(gate418inter0), .b(s_40), .O(gate418inter1));
  and2  gate829(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate830(.a(s_40), .O(gate418inter3));
  inv1  gate831(.a(s_41), .O(gate418inter4));
  nand2 gate832(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate833(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate834(.a(G32), .O(gate418inter7));
  inv1  gate835(.a(G1129), .O(gate418inter8));
  nand2 gate836(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate837(.a(s_41), .b(gate418inter3), .O(gate418inter10));
  nor2  gate838(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate839(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate840(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate813(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate814(.a(gate425inter0), .b(s_38), .O(gate425inter1));
  and2  gate815(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate816(.a(s_38), .O(gate425inter3));
  inv1  gate817(.a(s_39), .O(gate425inter4));
  nand2 gate818(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate819(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate820(.a(G4), .O(gate425inter7));
  inv1  gate821(.a(G1141), .O(gate425inter8));
  nand2 gate822(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate823(.a(s_39), .b(gate425inter3), .O(gate425inter10));
  nor2  gate824(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate825(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate826(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1149(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1150(.a(gate426inter0), .b(s_86), .O(gate426inter1));
  and2  gate1151(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1152(.a(s_86), .O(gate426inter3));
  inv1  gate1153(.a(s_87), .O(gate426inter4));
  nand2 gate1154(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1155(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1156(.a(G1045), .O(gate426inter7));
  inv1  gate1157(.a(G1141), .O(gate426inter8));
  nand2 gate1158(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1159(.a(s_87), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1160(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1161(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1162(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate841(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate842(.a(gate433inter0), .b(s_42), .O(gate433inter1));
  and2  gate843(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate844(.a(s_42), .O(gate433inter3));
  inv1  gate845(.a(s_43), .O(gate433inter4));
  nand2 gate846(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate847(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate848(.a(G8), .O(gate433inter7));
  inv1  gate849(.a(G1153), .O(gate433inter8));
  nand2 gate850(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate851(.a(s_43), .b(gate433inter3), .O(gate433inter10));
  nor2  gate852(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate853(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate854(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate925(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate926(.a(gate435inter0), .b(s_54), .O(gate435inter1));
  and2  gate927(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate928(.a(s_54), .O(gate435inter3));
  inv1  gate929(.a(s_55), .O(gate435inter4));
  nand2 gate930(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate931(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate932(.a(G9), .O(gate435inter7));
  inv1  gate933(.a(G1156), .O(gate435inter8));
  nand2 gate934(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate935(.a(s_55), .b(gate435inter3), .O(gate435inter10));
  nor2  gate936(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate937(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate938(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate673(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate674(.a(gate437inter0), .b(s_18), .O(gate437inter1));
  and2  gate675(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate676(.a(s_18), .O(gate437inter3));
  inv1  gate677(.a(s_19), .O(gate437inter4));
  nand2 gate678(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate679(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate680(.a(G10), .O(gate437inter7));
  inv1  gate681(.a(G1159), .O(gate437inter8));
  nand2 gate682(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate683(.a(s_19), .b(gate437inter3), .O(gate437inter10));
  nor2  gate684(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate685(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate686(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1079(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1080(.a(gate450inter0), .b(s_76), .O(gate450inter1));
  and2  gate1081(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1082(.a(s_76), .O(gate450inter3));
  inv1  gate1083(.a(s_77), .O(gate450inter4));
  nand2 gate1084(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1085(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1086(.a(G1081), .O(gate450inter7));
  inv1  gate1087(.a(G1177), .O(gate450inter8));
  nand2 gate1088(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1089(.a(s_77), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1090(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1091(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1092(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1009(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1010(.a(gate470inter0), .b(s_66), .O(gate470inter1));
  and2  gate1011(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1012(.a(s_66), .O(gate470inter3));
  inv1  gate1013(.a(s_67), .O(gate470inter4));
  nand2 gate1014(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1015(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1016(.a(G1111), .O(gate470inter7));
  inv1  gate1017(.a(G1207), .O(gate470inter8));
  nand2 gate1018(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1019(.a(s_67), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1020(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1021(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1022(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1107(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1108(.a(gate475inter0), .b(s_80), .O(gate475inter1));
  and2  gate1109(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1110(.a(s_80), .O(gate475inter3));
  inv1  gate1111(.a(s_81), .O(gate475inter4));
  nand2 gate1112(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1113(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1114(.a(G29), .O(gate475inter7));
  inv1  gate1115(.a(G1216), .O(gate475inter8));
  nand2 gate1116(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1117(.a(s_81), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1118(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1119(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1120(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1051(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1052(.a(gate487inter0), .b(s_72), .O(gate487inter1));
  and2  gate1053(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1054(.a(s_72), .O(gate487inter3));
  inv1  gate1055(.a(s_73), .O(gate487inter4));
  nand2 gate1056(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1057(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1058(.a(G1236), .O(gate487inter7));
  inv1  gate1059(.a(G1237), .O(gate487inter8));
  nand2 gate1060(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1061(.a(s_73), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1062(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1063(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1064(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate547(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate548(.a(gate502inter0), .b(s_0), .O(gate502inter1));
  and2  gate549(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate550(.a(s_0), .O(gate502inter3));
  inv1  gate551(.a(s_1), .O(gate502inter4));
  nand2 gate552(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate553(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate554(.a(G1266), .O(gate502inter7));
  inv1  gate555(.a(G1267), .O(gate502inter8));
  nand2 gate556(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate557(.a(s_1), .b(gate502inter3), .O(gate502inter10));
  nor2  gate558(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate559(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate560(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1233(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1234(.a(gate504inter0), .b(s_98), .O(gate504inter1));
  and2  gate1235(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1236(.a(s_98), .O(gate504inter3));
  inv1  gate1237(.a(s_99), .O(gate504inter4));
  nand2 gate1238(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1239(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1240(.a(G1270), .O(gate504inter7));
  inv1  gate1241(.a(G1271), .O(gate504inter8));
  nand2 gate1242(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1243(.a(s_99), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1244(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1245(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1246(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate967(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate968(.a(gate506inter0), .b(s_60), .O(gate506inter1));
  and2  gate969(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate970(.a(s_60), .O(gate506inter3));
  inv1  gate971(.a(s_61), .O(gate506inter4));
  nand2 gate972(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate973(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate974(.a(G1274), .O(gate506inter7));
  inv1  gate975(.a(G1275), .O(gate506inter8));
  nand2 gate976(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate977(.a(s_61), .b(gate506inter3), .O(gate506inter10));
  nor2  gate978(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate979(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate980(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate575(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate576(.a(gate511inter0), .b(s_4), .O(gate511inter1));
  and2  gate577(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate578(.a(s_4), .O(gate511inter3));
  inv1  gate579(.a(s_5), .O(gate511inter4));
  nand2 gate580(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate581(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate582(.a(G1284), .O(gate511inter7));
  inv1  gate583(.a(G1285), .O(gate511inter8));
  nand2 gate584(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate585(.a(s_5), .b(gate511inter3), .O(gate511inter10));
  nor2  gate586(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate587(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate588(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule