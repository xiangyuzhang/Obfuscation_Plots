module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2451(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2452(.a(gate10inter0), .b(s_272), .O(gate10inter1));
  and2  gate2453(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2454(.a(s_272), .O(gate10inter3));
  inv1  gate2455(.a(s_273), .O(gate10inter4));
  nand2 gate2456(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2457(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2458(.a(G3), .O(gate10inter7));
  inv1  gate2459(.a(G4), .O(gate10inter8));
  nand2 gate2460(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2461(.a(s_273), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2462(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2463(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2464(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2535(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2536(.a(gate13inter0), .b(s_284), .O(gate13inter1));
  and2  gate2537(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2538(.a(s_284), .O(gate13inter3));
  inv1  gate2539(.a(s_285), .O(gate13inter4));
  nand2 gate2540(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2541(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2542(.a(G9), .O(gate13inter7));
  inv1  gate2543(.a(G10), .O(gate13inter8));
  nand2 gate2544(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2545(.a(s_285), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2546(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2547(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2548(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1373(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1374(.a(gate14inter0), .b(s_118), .O(gate14inter1));
  and2  gate1375(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1376(.a(s_118), .O(gate14inter3));
  inv1  gate1377(.a(s_119), .O(gate14inter4));
  nand2 gate1378(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1379(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1380(.a(G11), .O(gate14inter7));
  inv1  gate1381(.a(G12), .O(gate14inter8));
  nand2 gate1382(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1383(.a(s_119), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1384(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1385(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1386(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2521(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2522(.a(gate16inter0), .b(s_282), .O(gate16inter1));
  and2  gate2523(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2524(.a(s_282), .O(gate16inter3));
  inv1  gate2525(.a(s_283), .O(gate16inter4));
  nand2 gate2526(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2527(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2528(.a(G15), .O(gate16inter7));
  inv1  gate2529(.a(G16), .O(gate16inter8));
  nand2 gate2530(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2531(.a(s_283), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2532(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2533(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2534(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2941(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2942(.a(gate20inter0), .b(s_342), .O(gate20inter1));
  and2  gate2943(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2944(.a(s_342), .O(gate20inter3));
  inv1  gate2945(.a(s_343), .O(gate20inter4));
  nand2 gate2946(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2947(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2948(.a(G23), .O(gate20inter7));
  inv1  gate2949(.a(G24), .O(gate20inter8));
  nand2 gate2950(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2951(.a(s_343), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2952(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2953(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2954(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate3039(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate3040(.a(gate21inter0), .b(s_356), .O(gate21inter1));
  and2  gate3041(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate3042(.a(s_356), .O(gate21inter3));
  inv1  gate3043(.a(s_357), .O(gate21inter4));
  nand2 gate3044(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate3045(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate3046(.a(G25), .O(gate21inter7));
  inv1  gate3047(.a(G26), .O(gate21inter8));
  nand2 gate3048(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate3049(.a(s_357), .b(gate21inter3), .O(gate21inter10));
  nor2  gate3050(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate3051(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate3052(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2829(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2830(.a(gate22inter0), .b(s_326), .O(gate22inter1));
  and2  gate2831(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2832(.a(s_326), .O(gate22inter3));
  inv1  gate2833(.a(s_327), .O(gate22inter4));
  nand2 gate2834(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2835(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2836(.a(G27), .O(gate22inter7));
  inv1  gate2837(.a(G28), .O(gate22inter8));
  nand2 gate2838(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2839(.a(s_327), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2840(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2841(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2842(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2773(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2774(.a(gate23inter0), .b(s_318), .O(gate23inter1));
  and2  gate2775(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2776(.a(s_318), .O(gate23inter3));
  inv1  gate2777(.a(s_319), .O(gate23inter4));
  nand2 gate2778(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2779(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2780(.a(G29), .O(gate23inter7));
  inv1  gate2781(.a(G30), .O(gate23inter8));
  nand2 gate2782(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2783(.a(s_319), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2784(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2785(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2786(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1457(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1458(.a(gate27inter0), .b(s_130), .O(gate27inter1));
  and2  gate1459(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1460(.a(s_130), .O(gate27inter3));
  inv1  gate1461(.a(s_131), .O(gate27inter4));
  nand2 gate1462(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1463(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1464(.a(G2), .O(gate27inter7));
  inv1  gate1465(.a(G6), .O(gate27inter8));
  nand2 gate1466(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1467(.a(s_131), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1468(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1469(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1470(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1261(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1262(.a(gate28inter0), .b(s_102), .O(gate28inter1));
  and2  gate1263(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1264(.a(s_102), .O(gate28inter3));
  inv1  gate1265(.a(s_103), .O(gate28inter4));
  nand2 gate1266(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1267(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1268(.a(G10), .O(gate28inter7));
  inv1  gate1269(.a(G14), .O(gate28inter8));
  nand2 gate1270(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1271(.a(s_103), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1272(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1273(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1274(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1009(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1010(.a(gate30inter0), .b(s_66), .O(gate30inter1));
  and2  gate1011(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1012(.a(s_66), .O(gate30inter3));
  inv1  gate1013(.a(s_67), .O(gate30inter4));
  nand2 gate1014(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1015(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1016(.a(G11), .O(gate30inter7));
  inv1  gate1017(.a(G15), .O(gate30inter8));
  nand2 gate1018(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1019(.a(s_67), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1020(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1021(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1022(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1891(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1892(.a(gate31inter0), .b(s_192), .O(gate31inter1));
  and2  gate1893(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1894(.a(s_192), .O(gate31inter3));
  inv1  gate1895(.a(s_193), .O(gate31inter4));
  nand2 gate1896(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1897(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1898(.a(G4), .O(gate31inter7));
  inv1  gate1899(.a(G8), .O(gate31inter8));
  nand2 gate1900(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1901(.a(s_193), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1902(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1903(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1904(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate2297(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2298(.a(gate32inter0), .b(s_250), .O(gate32inter1));
  and2  gate2299(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2300(.a(s_250), .O(gate32inter3));
  inv1  gate2301(.a(s_251), .O(gate32inter4));
  nand2 gate2302(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2303(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2304(.a(G12), .O(gate32inter7));
  inv1  gate2305(.a(G16), .O(gate32inter8));
  nand2 gate2306(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2307(.a(s_251), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2308(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2309(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2310(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1345(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1346(.a(gate33inter0), .b(s_114), .O(gate33inter1));
  and2  gate1347(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1348(.a(s_114), .O(gate33inter3));
  inv1  gate1349(.a(s_115), .O(gate33inter4));
  nand2 gate1350(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1351(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1352(.a(G17), .O(gate33inter7));
  inv1  gate1353(.a(G21), .O(gate33inter8));
  nand2 gate1354(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1355(.a(s_115), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1356(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1357(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1358(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1443(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1444(.a(gate36inter0), .b(s_128), .O(gate36inter1));
  and2  gate1445(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1446(.a(s_128), .O(gate36inter3));
  inv1  gate1447(.a(s_129), .O(gate36inter4));
  nand2 gate1448(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1449(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1450(.a(G26), .O(gate36inter7));
  inv1  gate1451(.a(G30), .O(gate36inter8));
  nand2 gate1452(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1453(.a(s_129), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1454(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1455(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1456(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1961(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1962(.a(gate41inter0), .b(s_202), .O(gate41inter1));
  and2  gate1963(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1964(.a(s_202), .O(gate41inter3));
  inv1  gate1965(.a(s_203), .O(gate41inter4));
  nand2 gate1966(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1967(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1968(.a(G1), .O(gate41inter7));
  inv1  gate1969(.a(G266), .O(gate41inter8));
  nand2 gate1970(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1971(.a(s_203), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1972(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1973(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1974(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1065(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1066(.a(gate47inter0), .b(s_74), .O(gate47inter1));
  and2  gate1067(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1068(.a(s_74), .O(gate47inter3));
  inv1  gate1069(.a(s_75), .O(gate47inter4));
  nand2 gate1070(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1071(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1072(.a(G7), .O(gate47inter7));
  inv1  gate1073(.a(G275), .O(gate47inter8));
  nand2 gate1074(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1075(.a(s_75), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1076(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1077(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1078(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2227(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2228(.a(gate51inter0), .b(s_240), .O(gate51inter1));
  and2  gate2229(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2230(.a(s_240), .O(gate51inter3));
  inv1  gate2231(.a(s_241), .O(gate51inter4));
  nand2 gate2232(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2233(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2234(.a(G11), .O(gate51inter7));
  inv1  gate2235(.a(G281), .O(gate51inter8));
  nand2 gate2236(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2237(.a(s_241), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2238(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2239(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2240(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate3123(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate3124(.a(gate56inter0), .b(s_368), .O(gate56inter1));
  and2  gate3125(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate3126(.a(s_368), .O(gate56inter3));
  inv1  gate3127(.a(s_369), .O(gate56inter4));
  nand2 gate3128(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate3129(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate3130(.a(G16), .O(gate56inter7));
  inv1  gate3131(.a(G287), .O(gate56inter8));
  nand2 gate3132(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate3133(.a(s_369), .b(gate56inter3), .O(gate56inter10));
  nor2  gate3134(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate3135(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate3136(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate841(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate842(.a(gate58inter0), .b(s_42), .O(gate58inter1));
  and2  gate843(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate844(.a(s_42), .O(gate58inter3));
  inv1  gate845(.a(s_43), .O(gate58inter4));
  nand2 gate846(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate847(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate848(.a(G18), .O(gate58inter7));
  inv1  gate849(.a(G290), .O(gate58inter8));
  nand2 gate850(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate851(.a(s_43), .b(gate58inter3), .O(gate58inter10));
  nor2  gate852(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate853(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate854(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1191(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1192(.a(gate62inter0), .b(s_92), .O(gate62inter1));
  and2  gate1193(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1194(.a(s_92), .O(gate62inter3));
  inv1  gate1195(.a(s_93), .O(gate62inter4));
  nand2 gate1196(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1197(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1198(.a(G22), .O(gate62inter7));
  inv1  gate1199(.a(G296), .O(gate62inter8));
  nand2 gate1200(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1201(.a(s_93), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1202(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1203(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1204(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2675(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2676(.a(gate63inter0), .b(s_304), .O(gate63inter1));
  and2  gate2677(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2678(.a(s_304), .O(gate63inter3));
  inv1  gate2679(.a(s_305), .O(gate63inter4));
  nand2 gate2680(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2681(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2682(.a(G23), .O(gate63inter7));
  inv1  gate2683(.a(G299), .O(gate63inter8));
  nand2 gate2684(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2685(.a(s_305), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2686(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2687(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2688(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate2045(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2046(.a(gate65inter0), .b(s_214), .O(gate65inter1));
  and2  gate2047(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2048(.a(s_214), .O(gate65inter3));
  inv1  gate2049(.a(s_215), .O(gate65inter4));
  nand2 gate2050(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2051(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2052(.a(G25), .O(gate65inter7));
  inv1  gate2053(.a(G302), .O(gate65inter8));
  nand2 gate2054(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2055(.a(s_215), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2056(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2057(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2058(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1079(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1080(.a(gate66inter0), .b(s_76), .O(gate66inter1));
  and2  gate1081(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1082(.a(s_76), .O(gate66inter3));
  inv1  gate1083(.a(s_77), .O(gate66inter4));
  nand2 gate1084(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1085(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1086(.a(G26), .O(gate66inter7));
  inv1  gate1087(.a(G302), .O(gate66inter8));
  nand2 gate1088(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1089(.a(s_77), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1090(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1091(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1092(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2101(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2102(.a(gate70inter0), .b(s_222), .O(gate70inter1));
  and2  gate2103(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2104(.a(s_222), .O(gate70inter3));
  inv1  gate2105(.a(s_223), .O(gate70inter4));
  nand2 gate2106(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2107(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2108(.a(G30), .O(gate70inter7));
  inv1  gate2109(.a(G308), .O(gate70inter8));
  nand2 gate2110(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2111(.a(s_223), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2112(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2113(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2114(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1597(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1598(.a(gate71inter0), .b(s_150), .O(gate71inter1));
  and2  gate1599(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1600(.a(s_150), .O(gate71inter3));
  inv1  gate1601(.a(s_151), .O(gate71inter4));
  nand2 gate1602(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1603(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1604(.a(G31), .O(gate71inter7));
  inv1  gate1605(.a(G311), .O(gate71inter8));
  nand2 gate1606(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1607(.a(s_151), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1608(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1609(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1610(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2395(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2396(.a(gate72inter0), .b(s_264), .O(gate72inter1));
  and2  gate2397(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2398(.a(s_264), .O(gate72inter3));
  inv1  gate2399(.a(s_265), .O(gate72inter4));
  nand2 gate2400(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2401(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2402(.a(G32), .O(gate72inter7));
  inv1  gate2403(.a(G311), .O(gate72inter8));
  nand2 gate2404(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2405(.a(s_265), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2406(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2407(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2408(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate883(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate884(.a(gate73inter0), .b(s_48), .O(gate73inter1));
  and2  gate885(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate886(.a(s_48), .O(gate73inter3));
  inv1  gate887(.a(s_49), .O(gate73inter4));
  nand2 gate888(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate889(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate890(.a(G1), .O(gate73inter7));
  inv1  gate891(.a(G314), .O(gate73inter8));
  nand2 gate892(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate893(.a(s_49), .b(gate73inter3), .O(gate73inter10));
  nor2  gate894(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate895(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate896(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2997(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2998(.a(gate78inter0), .b(s_350), .O(gate78inter1));
  and2  gate2999(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate3000(.a(s_350), .O(gate78inter3));
  inv1  gate3001(.a(s_351), .O(gate78inter4));
  nand2 gate3002(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate3003(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate3004(.a(G6), .O(gate78inter7));
  inv1  gate3005(.a(G320), .O(gate78inter8));
  nand2 gate3006(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate3007(.a(s_351), .b(gate78inter3), .O(gate78inter10));
  nor2  gate3008(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate3009(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate3010(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2073(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2074(.a(gate79inter0), .b(s_218), .O(gate79inter1));
  and2  gate2075(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2076(.a(s_218), .O(gate79inter3));
  inv1  gate2077(.a(s_219), .O(gate79inter4));
  nand2 gate2078(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2079(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2080(.a(G10), .O(gate79inter7));
  inv1  gate2081(.a(G323), .O(gate79inter8));
  nand2 gate2082(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2083(.a(s_219), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2084(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2085(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2086(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2605(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2606(.a(gate81inter0), .b(s_294), .O(gate81inter1));
  and2  gate2607(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2608(.a(s_294), .O(gate81inter3));
  inv1  gate2609(.a(s_295), .O(gate81inter4));
  nand2 gate2610(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2611(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2612(.a(G3), .O(gate81inter7));
  inv1  gate2613(.a(G326), .O(gate81inter8));
  nand2 gate2614(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2615(.a(s_295), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2616(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2617(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2618(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate2913(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2914(.a(gate83inter0), .b(s_338), .O(gate83inter1));
  and2  gate2915(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2916(.a(s_338), .O(gate83inter3));
  inv1  gate2917(.a(s_339), .O(gate83inter4));
  nand2 gate2918(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2919(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2920(.a(G11), .O(gate83inter7));
  inv1  gate2921(.a(G329), .O(gate83inter8));
  nand2 gate2922(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2923(.a(s_339), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2924(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2925(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2926(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate911(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate912(.a(gate86inter0), .b(s_52), .O(gate86inter1));
  and2  gate913(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate914(.a(s_52), .O(gate86inter3));
  inv1  gate915(.a(s_53), .O(gate86inter4));
  nand2 gate916(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate917(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate918(.a(G8), .O(gate86inter7));
  inv1  gate919(.a(G332), .O(gate86inter8));
  nand2 gate920(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate921(.a(s_53), .b(gate86inter3), .O(gate86inter10));
  nor2  gate922(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate923(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate924(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2269(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2270(.a(gate87inter0), .b(s_246), .O(gate87inter1));
  and2  gate2271(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2272(.a(s_246), .O(gate87inter3));
  inv1  gate2273(.a(s_247), .O(gate87inter4));
  nand2 gate2274(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2275(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2276(.a(G12), .O(gate87inter7));
  inv1  gate2277(.a(G335), .O(gate87inter8));
  nand2 gate2278(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2279(.a(s_247), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2280(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2281(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2282(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1135(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1136(.a(gate92inter0), .b(s_84), .O(gate92inter1));
  and2  gate1137(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1138(.a(s_84), .O(gate92inter3));
  inv1  gate1139(.a(s_85), .O(gate92inter4));
  nand2 gate1140(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1141(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1142(.a(G29), .O(gate92inter7));
  inv1  gate1143(.a(G341), .O(gate92inter8));
  nand2 gate1144(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1145(.a(s_85), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1146(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1147(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1148(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1849(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1850(.a(gate93inter0), .b(s_186), .O(gate93inter1));
  and2  gate1851(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1852(.a(s_186), .O(gate93inter3));
  inv1  gate1853(.a(s_187), .O(gate93inter4));
  nand2 gate1854(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1855(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1856(.a(G18), .O(gate93inter7));
  inv1  gate1857(.a(G344), .O(gate93inter8));
  nand2 gate1858(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1859(.a(s_187), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1860(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1861(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1862(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate785(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate786(.a(gate95inter0), .b(s_34), .O(gate95inter1));
  and2  gate787(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate788(.a(s_34), .O(gate95inter3));
  inv1  gate789(.a(s_35), .O(gate95inter4));
  nand2 gate790(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate791(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate792(.a(G26), .O(gate95inter7));
  inv1  gate793(.a(G347), .O(gate95inter8));
  nand2 gate794(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate795(.a(s_35), .b(gate95inter3), .O(gate95inter10));
  nor2  gate796(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate797(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate798(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1919(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1920(.a(gate97inter0), .b(s_196), .O(gate97inter1));
  and2  gate1921(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1922(.a(s_196), .O(gate97inter3));
  inv1  gate1923(.a(s_197), .O(gate97inter4));
  nand2 gate1924(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1925(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1926(.a(G19), .O(gate97inter7));
  inv1  gate1927(.a(G350), .O(gate97inter8));
  nand2 gate1928(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1929(.a(s_197), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1930(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1931(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1932(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate547(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate548(.a(gate103inter0), .b(s_0), .O(gate103inter1));
  and2  gate549(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate550(.a(s_0), .O(gate103inter3));
  inv1  gate551(.a(s_1), .O(gate103inter4));
  nand2 gate552(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate553(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate554(.a(G28), .O(gate103inter7));
  inv1  gate555(.a(G359), .O(gate103inter8));
  nand2 gate556(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate557(.a(s_1), .b(gate103inter3), .O(gate103inter10));
  nor2  gate558(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate559(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate560(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate631(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate632(.a(gate107inter0), .b(s_12), .O(gate107inter1));
  and2  gate633(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate634(.a(s_12), .O(gate107inter3));
  inv1  gate635(.a(s_13), .O(gate107inter4));
  nand2 gate636(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate637(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate638(.a(G366), .O(gate107inter7));
  inv1  gate639(.a(G367), .O(gate107inter8));
  nand2 gate640(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate641(.a(s_13), .b(gate107inter3), .O(gate107inter10));
  nor2  gate642(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate643(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate644(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1751(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1752(.a(gate110inter0), .b(s_172), .O(gate110inter1));
  and2  gate1753(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1754(.a(s_172), .O(gate110inter3));
  inv1  gate1755(.a(s_173), .O(gate110inter4));
  nand2 gate1756(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1757(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1758(.a(G372), .O(gate110inter7));
  inv1  gate1759(.a(G373), .O(gate110inter8));
  nand2 gate1760(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1761(.a(s_173), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1762(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1763(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1764(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1569(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1570(.a(gate112inter0), .b(s_146), .O(gate112inter1));
  and2  gate1571(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1572(.a(s_146), .O(gate112inter3));
  inv1  gate1573(.a(s_147), .O(gate112inter4));
  nand2 gate1574(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1575(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1576(.a(G376), .O(gate112inter7));
  inv1  gate1577(.a(G377), .O(gate112inter8));
  nand2 gate1578(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1579(.a(s_147), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1580(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1581(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1582(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate827(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate828(.a(gate113inter0), .b(s_40), .O(gate113inter1));
  and2  gate829(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate830(.a(s_40), .O(gate113inter3));
  inv1  gate831(.a(s_41), .O(gate113inter4));
  nand2 gate832(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate833(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate834(.a(G378), .O(gate113inter7));
  inv1  gate835(.a(G379), .O(gate113inter8));
  nand2 gate836(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate837(.a(s_41), .b(gate113inter3), .O(gate113inter10));
  nor2  gate838(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate839(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate840(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate2815(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2816(.a(gate114inter0), .b(s_324), .O(gate114inter1));
  and2  gate2817(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2818(.a(s_324), .O(gate114inter3));
  inv1  gate2819(.a(s_325), .O(gate114inter4));
  nand2 gate2820(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2821(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2822(.a(G380), .O(gate114inter7));
  inv1  gate2823(.a(G381), .O(gate114inter8));
  nand2 gate2824(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2825(.a(s_325), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2826(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2827(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2828(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1877(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1878(.a(gate116inter0), .b(s_190), .O(gate116inter1));
  and2  gate1879(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1880(.a(s_190), .O(gate116inter3));
  inv1  gate1881(.a(s_191), .O(gate116inter4));
  nand2 gate1882(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1883(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1884(.a(G384), .O(gate116inter7));
  inv1  gate1885(.a(G385), .O(gate116inter8));
  nand2 gate1886(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1887(.a(s_191), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1888(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1889(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1890(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1765(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1766(.a(gate118inter0), .b(s_174), .O(gate118inter1));
  and2  gate1767(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1768(.a(s_174), .O(gate118inter3));
  inv1  gate1769(.a(s_175), .O(gate118inter4));
  nand2 gate1770(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1771(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1772(.a(G388), .O(gate118inter7));
  inv1  gate1773(.a(G389), .O(gate118inter8));
  nand2 gate1774(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1775(.a(s_175), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1776(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1777(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1778(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2885(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2886(.a(gate119inter0), .b(s_334), .O(gate119inter1));
  and2  gate2887(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2888(.a(s_334), .O(gate119inter3));
  inv1  gate2889(.a(s_335), .O(gate119inter4));
  nand2 gate2890(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2891(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2892(.a(G390), .O(gate119inter7));
  inv1  gate2893(.a(G391), .O(gate119inter8));
  nand2 gate2894(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2895(.a(s_335), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2896(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2897(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2898(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate995(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate996(.a(gate120inter0), .b(s_64), .O(gate120inter1));
  and2  gate997(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate998(.a(s_64), .O(gate120inter3));
  inv1  gate999(.a(s_65), .O(gate120inter4));
  nand2 gate1000(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1001(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1002(.a(G392), .O(gate120inter7));
  inv1  gate1003(.a(G393), .O(gate120inter8));
  nand2 gate1004(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1005(.a(s_65), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1006(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1007(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1008(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate2213(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2214(.a(gate121inter0), .b(s_238), .O(gate121inter1));
  and2  gate2215(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2216(.a(s_238), .O(gate121inter3));
  inv1  gate2217(.a(s_239), .O(gate121inter4));
  nand2 gate2218(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2219(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2220(.a(G394), .O(gate121inter7));
  inv1  gate2221(.a(G395), .O(gate121inter8));
  nand2 gate2222(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2223(.a(s_239), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2224(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2225(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2226(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1205(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1206(.a(gate126inter0), .b(s_94), .O(gate126inter1));
  and2  gate1207(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1208(.a(s_94), .O(gate126inter3));
  inv1  gate1209(.a(s_95), .O(gate126inter4));
  nand2 gate1210(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1211(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1212(.a(G404), .O(gate126inter7));
  inv1  gate1213(.a(G405), .O(gate126inter8));
  nand2 gate1214(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1215(.a(s_95), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1216(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1217(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1218(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2437(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2438(.a(gate129inter0), .b(s_270), .O(gate129inter1));
  and2  gate2439(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2440(.a(s_270), .O(gate129inter3));
  inv1  gate2441(.a(s_271), .O(gate129inter4));
  nand2 gate2442(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2443(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2444(.a(G410), .O(gate129inter7));
  inv1  gate2445(.a(G411), .O(gate129inter8));
  nand2 gate2446(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2447(.a(s_271), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2448(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2449(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2450(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate2689(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2690(.a(gate133inter0), .b(s_306), .O(gate133inter1));
  and2  gate2691(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2692(.a(s_306), .O(gate133inter3));
  inv1  gate2693(.a(s_307), .O(gate133inter4));
  nand2 gate2694(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2695(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2696(.a(G418), .O(gate133inter7));
  inv1  gate2697(.a(G419), .O(gate133inter8));
  nand2 gate2698(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2699(.a(s_307), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2700(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2701(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2702(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate869(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate870(.a(gate137inter0), .b(s_46), .O(gate137inter1));
  and2  gate871(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate872(.a(s_46), .O(gate137inter3));
  inv1  gate873(.a(s_47), .O(gate137inter4));
  nand2 gate874(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate875(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate876(.a(G426), .O(gate137inter7));
  inv1  gate877(.a(G429), .O(gate137inter8));
  nand2 gate878(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate879(.a(s_47), .b(gate137inter3), .O(gate137inter10));
  nor2  gate880(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate881(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate882(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate2619(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2620(.a(gate138inter0), .b(s_296), .O(gate138inter1));
  and2  gate2621(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2622(.a(s_296), .O(gate138inter3));
  inv1  gate2623(.a(s_297), .O(gate138inter4));
  nand2 gate2624(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2625(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2626(.a(G432), .O(gate138inter7));
  inv1  gate2627(.a(G435), .O(gate138inter8));
  nand2 gate2628(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2629(.a(s_297), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2630(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2631(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2632(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1821(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1822(.a(gate139inter0), .b(s_182), .O(gate139inter1));
  and2  gate1823(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1824(.a(s_182), .O(gate139inter3));
  inv1  gate1825(.a(s_183), .O(gate139inter4));
  nand2 gate1826(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1827(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1828(.a(G438), .O(gate139inter7));
  inv1  gate1829(.a(G441), .O(gate139inter8));
  nand2 gate1830(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1831(.a(s_183), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1832(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1833(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1834(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2059(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2060(.a(gate140inter0), .b(s_216), .O(gate140inter1));
  and2  gate2061(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2062(.a(s_216), .O(gate140inter3));
  inv1  gate2063(.a(s_217), .O(gate140inter4));
  nand2 gate2064(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2065(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2066(.a(G444), .O(gate140inter7));
  inv1  gate2067(.a(G447), .O(gate140inter8));
  nand2 gate2068(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2069(.a(s_217), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2070(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2071(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2072(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1331(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1332(.a(gate142inter0), .b(s_112), .O(gate142inter1));
  and2  gate1333(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1334(.a(s_112), .O(gate142inter3));
  inv1  gate1335(.a(s_113), .O(gate142inter4));
  nand2 gate1336(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1337(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1338(.a(G456), .O(gate142inter7));
  inv1  gate1339(.a(G459), .O(gate142inter8));
  nand2 gate1340(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1341(.a(s_113), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1342(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1343(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1344(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate3025(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate3026(.a(gate143inter0), .b(s_354), .O(gate143inter1));
  and2  gate3027(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate3028(.a(s_354), .O(gate143inter3));
  inv1  gate3029(.a(s_355), .O(gate143inter4));
  nand2 gate3030(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate3031(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate3032(.a(G462), .O(gate143inter7));
  inv1  gate3033(.a(G465), .O(gate143inter8));
  nand2 gate3034(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate3035(.a(s_355), .b(gate143inter3), .O(gate143inter10));
  nor2  gate3036(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate3037(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate3038(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1975(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1976(.a(gate144inter0), .b(s_204), .O(gate144inter1));
  and2  gate1977(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1978(.a(s_204), .O(gate144inter3));
  inv1  gate1979(.a(s_205), .O(gate144inter4));
  nand2 gate1980(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1981(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1982(.a(G468), .O(gate144inter7));
  inv1  gate1983(.a(G471), .O(gate144inter8));
  nand2 gate1984(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1985(.a(s_205), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1986(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1987(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1988(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1611(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1612(.a(gate146inter0), .b(s_152), .O(gate146inter1));
  and2  gate1613(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1614(.a(s_152), .O(gate146inter3));
  inv1  gate1615(.a(s_153), .O(gate146inter4));
  nand2 gate1616(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1617(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1618(.a(G480), .O(gate146inter7));
  inv1  gate1619(.a(G483), .O(gate146inter8));
  nand2 gate1620(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1621(.a(s_153), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1622(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1623(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1624(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2563(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2564(.a(gate147inter0), .b(s_288), .O(gate147inter1));
  and2  gate2565(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2566(.a(s_288), .O(gate147inter3));
  inv1  gate2567(.a(s_289), .O(gate147inter4));
  nand2 gate2568(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2569(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2570(.a(G486), .O(gate147inter7));
  inv1  gate2571(.a(G489), .O(gate147inter8));
  nand2 gate2572(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2573(.a(s_289), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2574(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2575(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2576(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate673(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate674(.a(gate149inter0), .b(s_18), .O(gate149inter1));
  and2  gate675(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate676(.a(s_18), .O(gate149inter3));
  inv1  gate677(.a(s_19), .O(gate149inter4));
  nand2 gate678(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate679(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate680(.a(G498), .O(gate149inter7));
  inv1  gate681(.a(G501), .O(gate149inter8));
  nand2 gate682(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate683(.a(s_19), .b(gate149inter3), .O(gate149inter10));
  nor2  gate684(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate685(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate686(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2409(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2410(.a(gate150inter0), .b(s_266), .O(gate150inter1));
  and2  gate2411(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2412(.a(s_266), .O(gate150inter3));
  inv1  gate2413(.a(s_267), .O(gate150inter4));
  nand2 gate2414(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2415(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2416(.a(G504), .O(gate150inter7));
  inv1  gate2417(.a(G507), .O(gate150inter8));
  nand2 gate2418(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2419(.a(s_267), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2420(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2421(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2422(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2787(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2788(.a(gate153inter0), .b(s_320), .O(gate153inter1));
  and2  gate2789(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2790(.a(s_320), .O(gate153inter3));
  inv1  gate2791(.a(s_321), .O(gate153inter4));
  nand2 gate2792(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2793(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2794(.a(G426), .O(gate153inter7));
  inv1  gate2795(.a(G522), .O(gate153inter8));
  nand2 gate2796(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2797(.a(s_321), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2798(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2799(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2800(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1149(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1150(.a(gate155inter0), .b(s_86), .O(gate155inter1));
  and2  gate1151(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1152(.a(s_86), .O(gate155inter3));
  inv1  gate1153(.a(s_87), .O(gate155inter4));
  nand2 gate1154(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1155(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1156(.a(G432), .O(gate155inter7));
  inv1  gate1157(.a(G525), .O(gate155inter8));
  nand2 gate1158(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1159(.a(s_87), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1160(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1161(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1162(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate3109(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate3110(.a(gate159inter0), .b(s_366), .O(gate159inter1));
  and2  gate3111(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate3112(.a(s_366), .O(gate159inter3));
  inv1  gate3113(.a(s_367), .O(gate159inter4));
  nand2 gate3114(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate3115(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate3116(.a(G444), .O(gate159inter7));
  inv1  gate3117(.a(G531), .O(gate159inter8));
  nand2 gate3118(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate3119(.a(s_367), .b(gate159inter3), .O(gate159inter10));
  nor2  gate3120(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate3121(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate3122(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1415(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1416(.a(gate160inter0), .b(s_124), .O(gate160inter1));
  and2  gate1417(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1418(.a(s_124), .O(gate160inter3));
  inv1  gate1419(.a(s_125), .O(gate160inter4));
  nand2 gate1420(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1421(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1422(.a(G447), .O(gate160inter7));
  inv1  gate1423(.a(G531), .O(gate160inter8));
  nand2 gate1424(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1425(.a(s_125), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1426(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1427(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1428(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1653(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1654(.a(gate161inter0), .b(s_158), .O(gate161inter1));
  and2  gate1655(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1656(.a(s_158), .O(gate161inter3));
  inv1  gate1657(.a(s_159), .O(gate161inter4));
  nand2 gate1658(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1659(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1660(.a(G450), .O(gate161inter7));
  inv1  gate1661(.a(G534), .O(gate161inter8));
  nand2 gate1662(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1663(.a(s_159), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1664(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1665(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1666(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate3067(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate3068(.a(gate162inter0), .b(s_360), .O(gate162inter1));
  and2  gate3069(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate3070(.a(s_360), .O(gate162inter3));
  inv1  gate3071(.a(s_361), .O(gate162inter4));
  nand2 gate3072(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate3073(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate3074(.a(G453), .O(gate162inter7));
  inv1  gate3075(.a(G534), .O(gate162inter8));
  nand2 gate3076(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate3077(.a(s_361), .b(gate162inter3), .O(gate162inter10));
  nor2  gate3078(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate3079(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate3080(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2717(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2718(.a(gate164inter0), .b(s_310), .O(gate164inter1));
  and2  gate2719(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2720(.a(s_310), .O(gate164inter3));
  inv1  gate2721(.a(s_311), .O(gate164inter4));
  nand2 gate2722(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2723(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2724(.a(G459), .O(gate164inter7));
  inv1  gate2725(.a(G537), .O(gate164inter8));
  nand2 gate2726(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2727(.a(s_311), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2728(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2729(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2730(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1275(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1276(.a(gate166inter0), .b(s_104), .O(gate166inter1));
  and2  gate1277(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1278(.a(s_104), .O(gate166inter3));
  inv1  gate1279(.a(s_105), .O(gate166inter4));
  nand2 gate1280(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1281(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1282(.a(G465), .O(gate166inter7));
  inv1  gate1283(.a(G540), .O(gate166inter8));
  nand2 gate1284(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1285(.a(s_105), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1286(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1287(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1288(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2759(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2760(.a(gate167inter0), .b(s_316), .O(gate167inter1));
  and2  gate2761(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2762(.a(s_316), .O(gate167inter3));
  inv1  gate2763(.a(s_317), .O(gate167inter4));
  nand2 gate2764(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2765(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2766(.a(G468), .O(gate167inter7));
  inv1  gate2767(.a(G543), .O(gate167inter8));
  nand2 gate2768(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2769(.a(s_317), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2770(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2771(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2772(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate575(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate576(.a(gate171inter0), .b(s_4), .O(gate171inter1));
  and2  gate577(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate578(.a(s_4), .O(gate171inter3));
  inv1  gate579(.a(s_5), .O(gate171inter4));
  nand2 gate580(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate581(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate582(.a(G480), .O(gate171inter7));
  inv1  gate583(.a(G549), .O(gate171inter8));
  nand2 gate584(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate585(.a(s_5), .b(gate171inter3), .O(gate171inter10));
  nor2  gate586(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate587(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate588(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate2367(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2368(.a(gate172inter0), .b(s_260), .O(gate172inter1));
  and2  gate2369(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2370(.a(s_260), .O(gate172inter3));
  inv1  gate2371(.a(s_261), .O(gate172inter4));
  nand2 gate2372(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2373(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2374(.a(G483), .O(gate172inter7));
  inv1  gate2375(.a(G549), .O(gate172inter8));
  nand2 gate2376(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2377(.a(s_261), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2378(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2379(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2380(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2955(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2956(.a(gate176inter0), .b(s_344), .O(gate176inter1));
  and2  gate2957(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2958(.a(s_344), .O(gate176inter3));
  inv1  gate2959(.a(s_345), .O(gate176inter4));
  nand2 gate2960(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2961(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2962(.a(G495), .O(gate176inter7));
  inv1  gate2963(.a(G555), .O(gate176inter8));
  nand2 gate2964(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2965(.a(s_345), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2966(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2967(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2968(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1793(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1794(.a(gate180inter0), .b(s_178), .O(gate180inter1));
  and2  gate1795(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1796(.a(s_178), .O(gate180inter3));
  inv1  gate1797(.a(s_179), .O(gate180inter4));
  nand2 gate1798(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1799(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1800(.a(G507), .O(gate180inter7));
  inv1  gate1801(.a(G561), .O(gate180inter8));
  nand2 gate1802(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1803(.a(s_179), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1804(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1805(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1806(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1289(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1290(.a(gate182inter0), .b(s_106), .O(gate182inter1));
  and2  gate1291(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1292(.a(s_106), .O(gate182inter3));
  inv1  gate1293(.a(s_107), .O(gate182inter4));
  nand2 gate1294(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1295(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1296(.a(G513), .O(gate182inter7));
  inv1  gate1297(.a(G564), .O(gate182inter8));
  nand2 gate1298(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1299(.a(s_107), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1300(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1301(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1302(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1737(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1738(.a(gate184inter0), .b(s_170), .O(gate184inter1));
  and2  gate1739(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1740(.a(s_170), .O(gate184inter3));
  inv1  gate1741(.a(s_171), .O(gate184inter4));
  nand2 gate1742(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1743(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1744(.a(G519), .O(gate184inter7));
  inv1  gate1745(.a(G567), .O(gate184inter8));
  nand2 gate1746(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1747(.a(s_171), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1748(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1749(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1750(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1541(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1542(.a(gate187inter0), .b(s_142), .O(gate187inter1));
  and2  gate1543(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1544(.a(s_142), .O(gate187inter3));
  inv1  gate1545(.a(s_143), .O(gate187inter4));
  nand2 gate1546(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1547(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1548(.a(G574), .O(gate187inter7));
  inv1  gate1549(.a(G575), .O(gate187inter8));
  nand2 gate1550(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1551(.a(s_143), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1552(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1553(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1554(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1401(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1402(.a(gate188inter0), .b(s_122), .O(gate188inter1));
  and2  gate1403(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1404(.a(s_122), .O(gate188inter3));
  inv1  gate1405(.a(s_123), .O(gate188inter4));
  nand2 gate1406(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1407(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1408(.a(G576), .O(gate188inter7));
  inv1  gate1409(.a(G577), .O(gate188inter8));
  nand2 gate1410(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1411(.a(s_123), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1412(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1413(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1414(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2353(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2354(.a(gate189inter0), .b(s_258), .O(gate189inter1));
  and2  gate2355(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2356(.a(s_258), .O(gate189inter3));
  inv1  gate2357(.a(s_259), .O(gate189inter4));
  nand2 gate2358(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2359(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2360(.a(G578), .O(gate189inter7));
  inv1  gate2361(.a(G579), .O(gate189inter8));
  nand2 gate2362(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2363(.a(s_259), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2364(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2365(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2366(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate855(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate856(.a(gate190inter0), .b(s_44), .O(gate190inter1));
  and2  gate857(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate858(.a(s_44), .O(gate190inter3));
  inv1  gate859(.a(s_45), .O(gate190inter4));
  nand2 gate860(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate861(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate862(.a(G580), .O(gate190inter7));
  inv1  gate863(.a(G581), .O(gate190inter8));
  nand2 gate864(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate865(.a(s_45), .b(gate190inter3), .O(gate190inter10));
  nor2  gate866(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate867(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate868(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate2311(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2312(.a(gate194inter0), .b(s_252), .O(gate194inter1));
  and2  gate2313(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2314(.a(s_252), .O(gate194inter3));
  inv1  gate2315(.a(s_253), .O(gate194inter4));
  nand2 gate2316(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2317(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2318(.a(G588), .O(gate194inter7));
  inv1  gate2319(.a(G589), .O(gate194inter8));
  nand2 gate2320(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2321(.a(s_253), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2322(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2323(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2324(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1527(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1528(.a(gate195inter0), .b(s_140), .O(gate195inter1));
  and2  gate1529(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1530(.a(s_140), .O(gate195inter3));
  inv1  gate1531(.a(s_141), .O(gate195inter4));
  nand2 gate1532(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1533(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1534(.a(G590), .O(gate195inter7));
  inv1  gate1535(.a(G591), .O(gate195inter8));
  nand2 gate1536(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1537(.a(s_141), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1538(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1539(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1540(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2983(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2984(.a(gate198inter0), .b(s_348), .O(gate198inter1));
  and2  gate2985(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2986(.a(s_348), .O(gate198inter3));
  inv1  gate2987(.a(s_349), .O(gate198inter4));
  nand2 gate2988(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2989(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2990(.a(G596), .O(gate198inter7));
  inv1  gate2991(.a(G597), .O(gate198inter8));
  nand2 gate2992(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2993(.a(s_349), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2994(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2995(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2996(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2171(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2172(.a(gate205inter0), .b(s_232), .O(gate205inter1));
  and2  gate2173(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2174(.a(s_232), .O(gate205inter3));
  inv1  gate2175(.a(s_233), .O(gate205inter4));
  nand2 gate2176(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2177(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2178(.a(G622), .O(gate205inter7));
  inv1  gate2179(.a(G627), .O(gate205inter8));
  nand2 gate2180(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2181(.a(s_233), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2182(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2183(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2184(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1499(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1500(.a(gate206inter0), .b(s_136), .O(gate206inter1));
  and2  gate1501(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1502(.a(s_136), .O(gate206inter3));
  inv1  gate1503(.a(s_137), .O(gate206inter4));
  nand2 gate1504(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1505(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1506(.a(G632), .O(gate206inter7));
  inv1  gate1507(.a(G637), .O(gate206inter8));
  nand2 gate1508(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1509(.a(s_137), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1510(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1511(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1512(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1639(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1640(.a(gate207inter0), .b(s_156), .O(gate207inter1));
  and2  gate1641(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1642(.a(s_156), .O(gate207inter3));
  inv1  gate1643(.a(s_157), .O(gate207inter4));
  nand2 gate1644(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1645(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1646(.a(G622), .O(gate207inter7));
  inv1  gate1647(.a(G632), .O(gate207inter8));
  nand2 gate1648(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1649(.a(s_157), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1650(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1651(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1652(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1359(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1360(.a(gate208inter0), .b(s_116), .O(gate208inter1));
  and2  gate1361(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1362(.a(s_116), .O(gate208inter3));
  inv1  gate1363(.a(s_117), .O(gate208inter4));
  nand2 gate1364(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1365(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1366(.a(G627), .O(gate208inter7));
  inv1  gate1367(.a(G637), .O(gate208inter8));
  nand2 gate1368(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1369(.a(s_117), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1370(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1371(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1372(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate687(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate688(.a(gate210inter0), .b(s_20), .O(gate210inter1));
  and2  gate689(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate690(.a(s_20), .O(gate210inter3));
  inv1  gate691(.a(s_21), .O(gate210inter4));
  nand2 gate692(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate693(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate694(.a(G607), .O(gate210inter7));
  inv1  gate695(.a(G666), .O(gate210inter8));
  nand2 gate696(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate697(.a(s_21), .b(gate210inter3), .O(gate210inter10));
  nor2  gate698(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate699(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate700(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate3011(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate3012(.a(gate212inter0), .b(s_352), .O(gate212inter1));
  and2  gate3013(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate3014(.a(s_352), .O(gate212inter3));
  inv1  gate3015(.a(s_353), .O(gate212inter4));
  nand2 gate3016(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate3017(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate3018(.a(G617), .O(gate212inter7));
  inv1  gate3019(.a(G669), .O(gate212inter8));
  nand2 gate3020(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate3021(.a(s_353), .b(gate212inter3), .O(gate212inter10));
  nor2  gate3022(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate3023(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate3024(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate2115(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2116(.a(gate213inter0), .b(s_224), .O(gate213inter1));
  and2  gate2117(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2118(.a(s_224), .O(gate213inter3));
  inv1  gate2119(.a(s_225), .O(gate213inter4));
  nand2 gate2120(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2121(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2122(.a(G602), .O(gate213inter7));
  inv1  gate2123(.a(G672), .O(gate213inter8));
  nand2 gate2124(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2125(.a(s_225), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2126(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2127(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2128(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1947(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1948(.a(gate215inter0), .b(s_200), .O(gate215inter1));
  and2  gate1949(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1950(.a(s_200), .O(gate215inter3));
  inv1  gate1951(.a(s_201), .O(gate215inter4));
  nand2 gate1952(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1953(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1954(.a(G607), .O(gate215inter7));
  inv1  gate1955(.a(G675), .O(gate215inter8));
  nand2 gate1956(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1957(.a(s_201), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1958(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1959(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1960(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1555(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1556(.a(gate219inter0), .b(s_144), .O(gate219inter1));
  and2  gate1557(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1558(.a(s_144), .O(gate219inter3));
  inv1  gate1559(.a(s_145), .O(gate219inter4));
  nand2 gate1560(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1561(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1562(.a(G632), .O(gate219inter7));
  inv1  gate1563(.a(G681), .O(gate219inter8));
  nand2 gate1564(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1565(.a(s_145), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1566(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1567(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1568(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2927(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2928(.a(gate220inter0), .b(s_340), .O(gate220inter1));
  and2  gate2929(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2930(.a(s_340), .O(gate220inter3));
  inv1  gate2931(.a(s_341), .O(gate220inter4));
  nand2 gate2932(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2933(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2934(.a(G637), .O(gate220inter7));
  inv1  gate2935(.a(G681), .O(gate220inter8));
  nand2 gate2936(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2937(.a(s_341), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2938(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2939(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2940(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate2325(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2326(.a(gate221inter0), .b(s_254), .O(gate221inter1));
  and2  gate2327(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2328(.a(s_254), .O(gate221inter3));
  inv1  gate2329(.a(s_255), .O(gate221inter4));
  nand2 gate2330(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2331(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2332(.a(G622), .O(gate221inter7));
  inv1  gate2333(.a(G684), .O(gate221inter8));
  nand2 gate2334(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2335(.a(s_255), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2336(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2337(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2338(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate2465(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2466(.a(gate222inter0), .b(s_274), .O(gate222inter1));
  and2  gate2467(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2468(.a(s_274), .O(gate222inter3));
  inv1  gate2469(.a(s_275), .O(gate222inter4));
  nand2 gate2470(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2471(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2472(.a(G632), .O(gate222inter7));
  inv1  gate2473(.a(G684), .O(gate222inter8));
  nand2 gate2474(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2475(.a(s_275), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2476(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2477(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2478(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1247(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1248(.a(gate225inter0), .b(s_100), .O(gate225inter1));
  and2  gate1249(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1250(.a(s_100), .O(gate225inter3));
  inv1  gate1251(.a(s_101), .O(gate225inter4));
  nand2 gate1252(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1253(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1254(.a(G690), .O(gate225inter7));
  inv1  gate1255(.a(G691), .O(gate225inter8));
  nand2 gate1256(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1257(.a(s_101), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1258(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1259(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1260(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1933(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1934(.a(gate226inter0), .b(s_198), .O(gate226inter1));
  and2  gate1935(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1936(.a(s_198), .O(gate226inter3));
  inv1  gate1937(.a(s_199), .O(gate226inter4));
  nand2 gate1938(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1939(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1940(.a(G692), .O(gate226inter7));
  inv1  gate1941(.a(G693), .O(gate226inter8));
  nand2 gate1942(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1943(.a(s_199), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1944(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1945(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1946(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate967(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate968(.a(gate227inter0), .b(s_60), .O(gate227inter1));
  and2  gate969(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate970(.a(s_60), .O(gate227inter3));
  inv1  gate971(.a(s_61), .O(gate227inter4));
  nand2 gate972(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate973(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate974(.a(G694), .O(gate227inter7));
  inv1  gate975(.a(G695), .O(gate227inter8));
  nand2 gate976(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate977(.a(s_61), .b(gate227inter3), .O(gate227inter10));
  nor2  gate978(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate979(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate980(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1863(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1864(.a(gate229inter0), .b(s_188), .O(gate229inter1));
  and2  gate1865(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1866(.a(s_188), .O(gate229inter3));
  inv1  gate1867(.a(s_189), .O(gate229inter4));
  nand2 gate1868(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1869(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1870(.a(G698), .O(gate229inter7));
  inv1  gate1871(.a(G699), .O(gate229inter8));
  nand2 gate1872(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1873(.a(s_189), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1874(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1875(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1876(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate715(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate716(.a(gate230inter0), .b(s_24), .O(gate230inter1));
  and2  gate717(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate718(.a(s_24), .O(gate230inter3));
  inv1  gate719(.a(s_25), .O(gate230inter4));
  nand2 gate720(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate721(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate722(.a(G700), .O(gate230inter7));
  inv1  gate723(.a(G701), .O(gate230inter8));
  nand2 gate724(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate725(.a(s_25), .b(gate230inter3), .O(gate230inter10));
  nor2  gate726(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate727(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate728(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1485(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1486(.a(gate231inter0), .b(s_134), .O(gate231inter1));
  and2  gate1487(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1488(.a(s_134), .O(gate231inter3));
  inv1  gate1489(.a(s_135), .O(gate231inter4));
  nand2 gate1490(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1491(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1492(.a(G702), .O(gate231inter7));
  inv1  gate1493(.a(G703), .O(gate231inter8));
  nand2 gate1494(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1495(.a(s_135), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1496(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1497(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1498(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1163(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1164(.a(gate245inter0), .b(s_88), .O(gate245inter1));
  and2  gate1165(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1166(.a(s_88), .O(gate245inter3));
  inv1  gate1167(.a(s_89), .O(gate245inter4));
  nand2 gate1168(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1169(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1170(.a(G248), .O(gate245inter7));
  inv1  gate1171(.a(G736), .O(gate245inter8));
  nand2 gate1172(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1173(.a(s_89), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1174(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1175(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1176(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1471(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1472(.a(gate246inter0), .b(s_132), .O(gate246inter1));
  and2  gate1473(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1474(.a(s_132), .O(gate246inter3));
  inv1  gate1475(.a(s_133), .O(gate246inter4));
  nand2 gate1476(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1477(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1478(.a(G724), .O(gate246inter7));
  inv1  gate1479(.a(G736), .O(gate246inter8));
  nand2 gate1480(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1481(.a(s_133), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1482(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1483(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1484(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate561(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate562(.a(gate248inter0), .b(s_2), .O(gate248inter1));
  and2  gate563(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate564(.a(s_2), .O(gate248inter3));
  inv1  gate565(.a(s_3), .O(gate248inter4));
  nand2 gate566(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate567(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate568(.a(G727), .O(gate248inter7));
  inv1  gate569(.a(G739), .O(gate248inter8));
  nand2 gate570(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate571(.a(s_3), .b(gate248inter3), .O(gate248inter10));
  nor2  gate572(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate573(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate574(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate813(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate814(.a(gate254inter0), .b(s_38), .O(gate254inter1));
  and2  gate815(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate816(.a(s_38), .O(gate254inter3));
  inv1  gate817(.a(s_39), .O(gate254inter4));
  nand2 gate818(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate819(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate820(.a(G712), .O(gate254inter7));
  inv1  gate821(.a(G748), .O(gate254inter8));
  nand2 gate822(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate823(.a(s_39), .b(gate254inter3), .O(gate254inter10));
  nor2  gate824(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate825(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate826(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate925(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate926(.a(gate256inter0), .b(s_54), .O(gate256inter1));
  and2  gate927(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate928(.a(s_54), .O(gate256inter3));
  inv1  gate929(.a(s_55), .O(gate256inter4));
  nand2 gate930(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate931(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate932(.a(G715), .O(gate256inter7));
  inv1  gate933(.a(G751), .O(gate256inter8));
  nand2 gate934(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate935(.a(s_55), .b(gate256inter3), .O(gate256inter10));
  nor2  gate936(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate937(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate938(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate2185(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2186(.a(gate257inter0), .b(s_234), .O(gate257inter1));
  and2  gate2187(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2188(.a(s_234), .O(gate257inter3));
  inv1  gate2189(.a(s_235), .O(gate257inter4));
  nand2 gate2190(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2191(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2192(.a(G754), .O(gate257inter7));
  inv1  gate2193(.a(G755), .O(gate257inter8));
  nand2 gate2194(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2195(.a(s_235), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2196(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2197(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2198(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2899(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2900(.a(gate261inter0), .b(s_336), .O(gate261inter1));
  and2  gate2901(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2902(.a(s_336), .O(gate261inter3));
  inv1  gate2903(.a(s_337), .O(gate261inter4));
  nand2 gate2904(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2905(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2906(.a(G762), .O(gate261inter7));
  inv1  gate2907(.a(G763), .O(gate261inter8));
  nand2 gate2908(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2909(.a(s_337), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2910(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2911(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2912(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1023(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1024(.a(gate262inter0), .b(s_68), .O(gate262inter1));
  and2  gate1025(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1026(.a(s_68), .O(gate262inter3));
  inv1  gate1027(.a(s_69), .O(gate262inter4));
  nand2 gate1028(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1029(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1030(.a(G764), .O(gate262inter7));
  inv1  gate1031(.a(G765), .O(gate262inter8));
  nand2 gate1032(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1033(.a(s_69), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1034(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1035(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1036(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2493(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2494(.a(gate264inter0), .b(s_278), .O(gate264inter1));
  and2  gate2495(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2496(.a(s_278), .O(gate264inter3));
  inv1  gate2497(.a(s_279), .O(gate264inter4));
  nand2 gate2498(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2499(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2500(.a(G768), .O(gate264inter7));
  inv1  gate2501(.a(G769), .O(gate264inter8));
  nand2 gate2502(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2503(.a(s_279), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2504(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2505(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2506(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1989(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1990(.a(gate265inter0), .b(s_206), .O(gate265inter1));
  and2  gate1991(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1992(.a(s_206), .O(gate265inter3));
  inv1  gate1993(.a(s_207), .O(gate265inter4));
  nand2 gate1994(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1995(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1996(.a(G642), .O(gate265inter7));
  inv1  gate1997(.a(G770), .O(gate265inter8));
  nand2 gate1998(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1999(.a(s_207), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2000(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2001(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2002(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1121(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1122(.a(gate269inter0), .b(s_82), .O(gate269inter1));
  and2  gate1123(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1124(.a(s_82), .O(gate269inter3));
  inv1  gate1125(.a(s_83), .O(gate269inter4));
  nand2 gate1126(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1127(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1128(.a(G654), .O(gate269inter7));
  inv1  gate1129(.a(G782), .O(gate269inter8));
  nand2 gate1130(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1131(.a(s_83), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1132(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1133(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1134(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1905(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1906(.a(gate271inter0), .b(s_194), .O(gate271inter1));
  and2  gate1907(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1908(.a(s_194), .O(gate271inter3));
  inv1  gate1909(.a(s_195), .O(gate271inter4));
  nand2 gate1910(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1911(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1912(.a(G660), .O(gate271inter7));
  inv1  gate1913(.a(G788), .O(gate271inter8));
  nand2 gate1914(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1915(.a(s_195), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1916(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1917(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1918(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2969(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2970(.a(gate272inter0), .b(s_346), .O(gate272inter1));
  and2  gate2971(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2972(.a(s_346), .O(gate272inter3));
  inv1  gate2973(.a(s_347), .O(gate272inter4));
  nand2 gate2974(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2975(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2976(.a(G663), .O(gate272inter7));
  inv1  gate2977(.a(G791), .O(gate272inter8));
  nand2 gate2978(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2979(.a(s_347), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2980(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2981(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2982(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2647(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2648(.a(gate274inter0), .b(s_300), .O(gate274inter1));
  and2  gate2649(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2650(.a(s_300), .O(gate274inter3));
  inv1  gate2651(.a(s_301), .O(gate274inter4));
  nand2 gate2652(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2653(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2654(.a(G770), .O(gate274inter7));
  inv1  gate2655(.a(G794), .O(gate274inter8));
  nand2 gate2656(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2657(.a(s_301), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2658(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2659(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2660(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate743(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate744(.a(gate277inter0), .b(s_28), .O(gate277inter1));
  and2  gate745(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate746(.a(s_28), .O(gate277inter3));
  inv1  gate747(.a(s_29), .O(gate277inter4));
  nand2 gate748(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate749(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate750(.a(G648), .O(gate277inter7));
  inv1  gate751(.a(G800), .O(gate277inter8));
  nand2 gate752(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate753(.a(s_29), .b(gate277inter3), .O(gate277inter10));
  nor2  gate754(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate755(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate756(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate3081(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate3082(.a(gate282inter0), .b(s_362), .O(gate282inter1));
  and2  gate3083(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate3084(.a(s_362), .O(gate282inter3));
  inv1  gate3085(.a(s_363), .O(gate282inter4));
  nand2 gate3086(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate3087(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate3088(.a(G782), .O(gate282inter7));
  inv1  gate3089(.a(G806), .O(gate282inter8));
  nand2 gate3090(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate3091(.a(s_363), .b(gate282inter3), .O(gate282inter10));
  nor2  gate3092(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate3093(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate3094(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1303(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1304(.a(gate284inter0), .b(s_108), .O(gate284inter1));
  and2  gate1305(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1306(.a(s_108), .O(gate284inter3));
  inv1  gate1307(.a(s_109), .O(gate284inter4));
  nand2 gate1308(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1309(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1310(.a(G785), .O(gate284inter7));
  inv1  gate1311(.a(G809), .O(gate284inter8));
  nand2 gate1312(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1313(.a(s_109), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1314(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1315(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1316(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1219(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1220(.a(gate291inter0), .b(s_96), .O(gate291inter1));
  and2  gate1221(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1222(.a(s_96), .O(gate291inter3));
  inv1  gate1223(.a(s_97), .O(gate291inter4));
  nand2 gate1224(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1225(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1226(.a(G822), .O(gate291inter7));
  inv1  gate1227(.a(G823), .O(gate291inter8));
  nand2 gate1228(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1229(.a(s_97), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1230(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1231(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1232(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate589(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate590(.a(gate295inter0), .b(s_6), .O(gate295inter1));
  and2  gate591(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate592(.a(s_6), .O(gate295inter3));
  inv1  gate593(.a(s_7), .O(gate295inter4));
  nand2 gate594(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate595(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate596(.a(G830), .O(gate295inter7));
  inv1  gate597(.a(G831), .O(gate295inter8));
  nand2 gate598(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate599(.a(s_7), .b(gate295inter3), .O(gate295inter10));
  nor2  gate600(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate601(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate602(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1429(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1430(.a(gate296inter0), .b(s_126), .O(gate296inter1));
  and2  gate1431(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1432(.a(s_126), .O(gate296inter3));
  inv1  gate1433(.a(s_127), .O(gate296inter4));
  nand2 gate1434(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1435(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1436(.a(G826), .O(gate296inter7));
  inv1  gate1437(.a(G827), .O(gate296inter8));
  nand2 gate1438(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1439(.a(s_127), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1440(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1441(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1442(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2731(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2732(.a(gate387inter0), .b(s_312), .O(gate387inter1));
  and2  gate2733(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2734(.a(s_312), .O(gate387inter3));
  inv1  gate2735(.a(s_313), .O(gate387inter4));
  nand2 gate2736(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2737(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2738(.a(G1), .O(gate387inter7));
  inv1  gate2739(.a(G1036), .O(gate387inter8));
  nand2 gate2740(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2741(.a(s_313), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2742(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2743(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2744(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate701(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate702(.a(gate388inter0), .b(s_22), .O(gate388inter1));
  and2  gate703(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate704(.a(s_22), .O(gate388inter3));
  inv1  gate705(.a(s_23), .O(gate388inter4));
  nand2 gate706(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate707(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate708(.a(G2), .O(gate388inter7));
  inv1  gate709(.a(G1039), .O(gate388inter8));
  nand2 gate710(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate711(.a(s_23), .b(gate388inter3), .O(gate388inter10));
  nor2  gate712(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate713(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate714(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2507(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2508(.a(gate389inter0), .b(s_280), .O(gate389inter1));
  and2  gate2509(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2510(.a(s_280), .O(gate389inter3));
  inv1  gate2511(.a(s_281), .O(gate389inter4));
  nand2 gate2512(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2513(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2514(.a(G3), .O(gate389inter7));
  inv1  gate2515(.a(G1042), .O(gate389inter8));
  nand2 gate2516(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2517(.a(s_281), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2518(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2519(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2520(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate617(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate618(.a(gate391inter0), .b(s_10), .O(gate391inter1));
  and2  gate619(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate620(.a(s_10), .O(gate391inter3));
  inv1  gate621(.a(s_11), .O(gate391inter4));
  nand2 gate622(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate623(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate624(.a(G5), .O(gate391inter7));
  inv1  gate625(.a(G1048), .O(gate391inter8));
  nand2 gate626(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate627(.a(s_11), .b(gate391inter3), .O(gate391inter10));
  nor2  gate628(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate629(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate630(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2423(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2424(.a(gate393inter0), .b(s_268), .O(gate393inter1));
  and2  gate2425(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2426(.a(s_268), .O(gate393inter3));
  inv1  gate2427(.a(s_269), .O(gate393inter4));
  nand2 gate2428(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2429(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2430(.a(G7), .O(gate393inter7));
  inv1  gate2431(.a(G1054), .O(gate393inter8));
  nand2 gate2432(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2433(.a(s_269), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2434(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2435(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2436(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1317(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1318(.a(gate395inter0), .b(s_110), .O(gate395inter1));
  and2  gate1319(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1320(.a(s_110), .O(gate395inter3));
  inv1  gate1321(.a(s_111), .O(gate395inter4));
  nand2 gate1322(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1323(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1324(.a(G9), .O(gate395inter7));
  inv1  gate1325(.a(G1060), .O(gate395inter8));
  nand2 gate1326(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1327(.a(s_111), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1328(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1329(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1330(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1093(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1094(.a(gate397inter0), .b(s_78), .O(gate397inter1));
  and2  gate1095(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1096(.a(s_78), .O(gate397inter3));
  inv1  gate1097(.a(s_79), .O(gate397inter4));
  nand2 gate1098(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1099(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1100(.a(G11), .O(gate397inter7));
  inv1  gate1101(.a(G1066), .O(gate397inter8));
  nand2 gate1102(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1103(.a(s_79), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1104(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1105(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1106(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2031(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2032(.a(gate398inter0), .b(s_212), .O(gate398inter1));
  and2  gate2033(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2034(.a(s_212), .O(gate398inter3));
  inv1  gate2035(.a(s_213), .O(gate398inter4));
  nand2 gate2036(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2037(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2038(.a(G12), .O(gate398inter7));
  inv1  gate2039(.a(G1069), .O(gate398inter8));
  nand2 gate2040(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2041(.a(s_213), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2042(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2043(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2044(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2087(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2088(.a(gate400inter0), .b(s_220), .O(gate400inter1));
  and2  gate2089(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2090(.a(s_220), .O(gate400inter3));
  inv1  gate2091(.a(s_221), .O(gate400inter4));
  nand2 gate2092(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2093(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2094(.a(G14), .O(gate400inter7));
  inv1  gate2095(.a(G1075), .O(gate400inter8));
  nand2 gate2096(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2097(.a(s_221), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2098(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2099(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2100(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate3095(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate3096(.a(gate402inter0), .b(s_364), .O(gate402inter1));
  and2  gate3097(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate3098(.a(s_364), .O(gate402inter3));
  inv1  gate3099(.a(s_365), .O(gate402inter4));
  nand2 gate3100(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate3101(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate3102(.a(G16), .O(gate402inter7));
  inv1  gate3103(.a(G1081), .O(gate402inter8));
  nand2 gate3104(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate3105(.a(s_365), .b(gate402inter3), .O(gate402inter10));
  nor2  gate3106(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate3107(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate3108(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate981(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate982(.a(gate405inter0), .b(s_62), .O(gate405inter1));
  and2  gate983(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate984(.a(s_62), .O(gate405inter3));
  inv1  gate985(.a(s_63), .O(gate405inter4));
  nand2 gate986(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate987(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate988(.a(G19), .O(gate405inter7));
  inv1  gate989(.a(G1090), .O(gate405inter8));
  nand2 gate990(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate991(.a(s_63), .b(gate405inter3), .O(gate405inter10));
  nor2  gate992(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate993(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate994(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1051(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1052(.a(gate410inter0), .b(s_72), .O(gate410inter1));
  and2  gate1053(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1054(.a(s_72), .O(gate410inter3));
  inv1  gate1055(.a(s_73), .O(gate410inter4));
  nand2 gate1056(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1057(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1058(.a(G24), .O(gate410inter7));
  inv1  gate1059(.a(G1105), .O(gate410inter8));
  nand2 gate1060(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1061(.a(s_73), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1062(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1063(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1064(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1835(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1836(.a(gate411inter0), .b(s_184), .O(gate411inter1));
  and2  gate1837(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1838(.a(s_184), .O(gate411inter3));
  inv1  gate1839(.a(s_185), .O(gate411inter4));
  nand2 gate1840(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1841(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1842(.a(G25), .O(gate411inter7));
  inv1  gate1843(.a(G1108), .O(gate411inter8));
  nand2 gate1844(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1845(.a(s_185), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1846(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1847(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1848(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2199(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2200(.a(gate414inter0), .b(s_236), .O(gate414inter1));
  and2  gate2201(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2202(.a(s_236), .O(gate414inter3));
  inv1  gate2203(.a(s_237), .O(gate414inter4));
  nand2 gate2204(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2205(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2206(.a(G28), .O(gate414inter7));
  inv1  gate2207(.a(G1117), .O(gate414inter8));
  nand2 gate2208(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2209(.a(s_237), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2210(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2211(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2212(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate757(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate758(.a(gate417inter0), .b(s_30), .O(gate417inter1));
  and2  gate759(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate760(.a(s_30), .O(gate417inter3));
  inv1  gate761(.a(s_31), .O(gate417inter4));
  nand2 gate762(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate763(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate764(.a(G31), .O(gate417inter7));
  inv1  gate765(.a(G1126), .O(gate417inter8));
  nand2 gate766(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate767(.a(s_31), .b(gate417inter3), .O(gate417inter10));
  nor2  gate768(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate769(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate770(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate771(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate772(.a(gate419inter0), .b(s_32), .O(gate419inter1));
  and2  gate773(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate774(.a(s_32), .O(gate419inter3));
  inv1  gate775(.a(s_33), .O(gate419inter4));
  nand2 gate776(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate777(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate778(.a(G1), .O(gate419inter7));
  inv1  gate779(.a(G1132), .O(gate419inter8));
  nand2 gate780(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate781(.a(s_33), .b(gate419inter3), .O(gate419inter10));
  nor2  gate782(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate783(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate784(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2577(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2578(.a(gate428inter0), .b(s_290), .O(gate428inter1));
  and2  gate2579(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2580(.a(s_290), .O(gate428inter3));
  inv1  gate2581(.a(s_291), .O(gate428inter4));
  nand2 gate2582(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2583(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2584(.a(G1048), .O(gate428inter7));
  inv1  gate2585(.a(G1144), .O(gate428inter8));
  nand2 gate2586(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2587(.a(s_291), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2588(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2589(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2590(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2843(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2844(.a(gate431inter0), .b(s_328), .O(gate431inter1));
  and2  gate2845(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2846(.a(s_328), .O(gate431inter3));
  inv1  gate2847(.a(s_329), .O(gate431inter4));
  nand2 gate2848(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2849(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2850(.a(G7), .O(gate431inter7));
  inv1  gate2851(.a(G1150), .O(gate431inter8));
  nand2 gate2852(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2853(.a(s_329), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2854(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2855(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2856(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2857(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2858(.a(gate432inter0), .b(s_330), .O(gate432inter1));
  and2  gate2859(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2860(.a(s_330), .O(gate432inter3));
  inv1  gate2861(.a(s_331), .O(gate432inter4));
  nand2 gate2862(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2863(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2864(.a(G1054), .O(gate432inter7));
  inv1  gate2865(.a(G1150), .O(gate432inter8));
  nand2 gate2866(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2867(.a(s_331), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2868(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2869(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2870(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1723(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1724(.a(gate435inter0), .b(s_168), .O(gate435inter1));
  and2  gate1725(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1726(.a(s_168), .O(gate435inter3));
  inv1  gate1727(.a(s_169), .O(gate435inter4));
  nand2 gate1728(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1729(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1730(.a(G9), .O(gate435inter7));
  inv1  gate1731(.a(G1156), .O(gate435inter8));
  nand2 gate1732(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1733(.a(s_169), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1734(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1735(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1736(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2703(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2704(.a(gate438inter0), .b(s_308), .O(gate438inter1));
  and2  gate2705(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2706(.a(s_308), .O(gate438inter3));
  inv1  gate2707(.a(s_309), .O(gate438inter4));
  nand2 gate2708(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2709(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2710(.a(G1063), .O(gate438inter7));
  inv1  gate2711(.a(G1159), .O(gate438inter8));
  nand2 gate2712(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2713(.a(s_309), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2714(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2715(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2716(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate603(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate604(.a(gate439inter0), .b(s_8), .O(gate439inter1));
  and2  gate605(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate606(.a(s_8), .O(gate439inter3));
  inv1  gate607(.a(s_9), .O(gate439inter4));
  nand2 gate608(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate609(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate610(.a(G11), .O(gate439inter7));
  inv1  gate611(.a(G1162), .O(gate439inter8));
  nand2 gate612(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate613(.a(s_9), .b(gate439inter3), .O(gate439inter10));
  nor2  gate614(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate615(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate616(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2479(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2480(.a(gate441inter0), .b(s_276), .O(gate441inter1));
  and2  gate2481(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2482(.a(s_276), .O(gate441inter3));
  inv1  gate2483(.a(s_277), .O(gate441inter4));
  nand2 gate2484(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2485(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2486(.a(G12), .O(gate441inter7));
  inv1  gate2487(.a(G1165), .O(gate441inter8));
  nand2 gate2488(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2489(.a(s_277), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2490(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2491(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2492(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2157(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2158(.a(gate443inter0), .b(s_230), .O(gate443inter1));
  and2  gate2159(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2160(.a(s_230), .O(gate443inter3));
  inv1  gate2161(.a(s_231), .O(gate443inter4));
  nand2 gate2162(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2163(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2164(.a(G13), .O(gate443inter7));
  inv1  gate2165(.a(G1168), .O(gate443inter8));
  nand2 gate2166(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2167(.a(s_231), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2168(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2169(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2170(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate2143(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2144(.a(gate447inter0), .b(s_228), .O(gate447inter1));
  and2  gate2145(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2146(.a(s_228), .O(gate447inter3));
  inv1  gate2147(.a(s_229), .O(gate447inter4));
  nand2 gate2148(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2149(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2150(.a(G15), .O(gate447inter7));
  inv1  gate2151(.a(G1174), .O(gate447inter8));
  nand2 gate2152(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2153(.a(s_229), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2154(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2155(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2156(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1107(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1108(.a(gate448inter0), .b(s_80), .O(gate448inter1));
  and2  gate1109(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1110(.a(s_80), .O(gate448inter3));
  inv1  gate1111(.a(s_81), .O(gate448inter4));
  nand2 gate1112(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1113(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1114(.a(G1078), .O(gate448inter7));
  inv1  gate1115(.a(G1174), .O(gate448inter8));
  nand2 gate1116(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1117(.a(s_81), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1118(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1119(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1120(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1233(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1234(.a(gate449inter0), .b(s_98), .O(gate449inter1));
  and2  gate1235(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1236(.a(s_98), .O(gate449inter3));
  inv1  gate1237(.a(s_99), .O(gate449inter4));
  nand2 gate1238(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1239(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1240(.a(G16), .O(gate449inter7));
  inv1  gate1241(.a(G1177), .O(gate449inter8));
  nand2 gate1242(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1243(.a(s_99), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1244(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1245(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1246(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate2549(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2550(.a(gate450inter0), .b(s_286), .O(gate450inter1));
  and2  gate2551(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2552(.a(s_286), .O(gate450inter3));
  inv1  gate2553(.a(s_287), .O(gate450inter4));
  nand2 gate2554(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2555(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2556(.a(G1081), .O(gate450inter7));
  inv1  gate2557(.a(G1177), .O(gate450inter8));
  nand2 gate2558(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2559(.a(s_287), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2560(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2561(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2562(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2633(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2634(.a(gate454inter0), .b(s_298), .O(gate454inter1));
  and2  gate2635(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2636(.a(s_298), .O(gate454inter3));
  inv1  gate2637(.a(s_299), .O(gate454inter4));
  nand2 gate2638(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2639(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2640(.a(G1087), .O(gate454inter7));
  inv1  gate2641(.a(G1183), .O(gate454inter8));
  nand2 gate2642(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2643(.a(s_299), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2644(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2645(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2646(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1513(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1514(.a(gate456inter0), .b(s_138), .O(gate456inter1));
  and2  gate1515(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1516(.a(s_138), .O(gate456inter3));
  inv1  gate1517(.a(s_139), .O(gate456inter4));
  nand2 gate1518(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1519(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1520(.a(G1090), .O(gate456inter7));
  inv1  gate1521(.a(G1186), .O(gate456inter8));
  nand2 gate1522(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1523(.a(s_139), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1524(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1525(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1526(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1583(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1584(.a(gate458inter0), .b(s_148), .O(gate458inter1));
  and2  gate1585(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1586(.a(s_148), .O(gate458inter3));
  inv1  gate1587(.a(s_149), .O(gate458inter4));
  nand2 gate1588(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1589(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1590(.a(G1093), .O(gate458inter7));
  inv1  gate1591(.a(G1189), .O(gate458inter8));
  nand2 gate1592(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1593(.a(s_149), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1594(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1595(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1596(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1807(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1808(.a(gate459inter0), .b(s_180), .O(gate459inter1));
  and2  gate1809(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1810(.a(s_180), .O(gate459inter3));
  inv1  gate1811(.a(s_181), .O(gate459inter4));
  nand2 gate1812(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1813(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1814(.a(G21), .O(gate459inter7));
  inv1  gate1815(.a(G1192), .O(gate459inter8));
  nand2 gate1816(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1817(.a(s_181), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1818(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1819(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1820(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2801(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2802(.a(gate461inter0), .b(s_322), .O(gate461inter1));
  and2  gate2803(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2804(.a(s_322), .O(gate461inter3));
  inv1  gate2805(.a(s_323), .O(gate461inter4));
  nand2 gate2806(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2807(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2808(.a(G22), .O(gate461inter7));
  inv1  gate2809(.a(G1195), .O(gate461inter8));
  nand2 gate2810(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2811(.a(s_323), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2812(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2813(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2814(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate659(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate660(.a(gate462inter0), .b(s_16), .O(gate462inter1));
  and2  gate661(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate662(.a(s_16), .O(gate462inter3));
  inv1  gate663(.a(s_17), .O(gate462inter4));
  nand2 gate664(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate665(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate666(.a(G1099), .O(gate462inter7));
  inv1  gate667(.a(G1195), .O(gate462inter8));
  nand2 gate668(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate669(.a(s_17), .b(gate462inter3), .O(gate462inter10));
  nor2  gate670(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate671(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate672(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2241(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2242(.a(gate463inter0), .b(s_242), .O(gate463inter1));
  and2  gate2243(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2244(.a(s_242), .O(gate463inter3));
  inv1  gate2245(.a(s_243), .O(gate463inter4));
  nand2 gate2246(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2247(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2248(.a(G23), .O(gate463inter7));
  inv1  gate2249(.a(G1198), .O(gate463inter8));
  nand2 gate2250(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2251(.a(s_243), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2252(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2253(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2254(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2745(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2746(.a(gate465inter0), .b(s_314), .O(gate465inter1));
  and2  gate2747(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2748(.a(s_314), .O(gate465inter3));
  inv1  gate2749(.a(s_315), .O(gate465inter4));
  nand2 gate2750(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2751(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2752(.a(G24), .O(gate465inter7));
  inv1  gate2753(.a(G1201), .O(gate465inter8));
  nand2 gate2754(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2755(.a(s_315), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2756(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2757(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2758(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2661(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2662(.a(gate469inter0), .b(s_302), .O(gate469inter1));
  and2  gate2663(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2664(.a(s_302), .O(gate469inter3));
  inv1  gate2665(.a(s_303), .O(gate469inter4));
  nand2 gate2666(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2667(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2668(.a(G26), .O(gate469inter7));
  inv1  gate2669(.a(G1207), .O(gate469inter8));
  nand2 gate2670(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2671(.a(s_303), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2672(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2673(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2674(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1177(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1178(.a(gate471inter0), .b(s_90), .O(gate471inter1));
  and2  gate1179(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1180(.a(s_90), .O(gate471inter3));
  inv1  gate1181(.a(s_91), .O(gate471inter4));
  nand2 gate1182(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1183(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1184(.a(G27), .O(gate471inter7));
  inv1  gate1185(.a(G1210), .O(gate471inter8));
  nand2 gate1186(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1187(.a(s_91), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1188(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1189(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1190(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate3137(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate3138(.a(gate472inter0), .b(s_370), .O(gate472inter1));
  and2  gate3139(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate3140(.a(s_370), .O(gate472inter3));
  inv1  gate3141(.a(s_371), .O(gate472inter4));
  nand2 gate3142(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate3143(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate3144(.a(G1114), .O(gate472inter7));
  inv1  gate3145(.a(G1210), .O(gate472inter8));
  nand2 gate3146(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate3147(.a(s_371), .b(gate472inter3), .O(gate472inter10));
  nor2  gate3148(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate3149(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate3150(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate2283(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2284(.a(gate473inter0), .b(s_248), .O(gate473inter1));
  and2  gate2285(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2286(.a(s_248), .O(gate473inter3));
  inv1  gate2287(.a(s_249), .O(gate473inter4));
  nand2 gate2288(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2289(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2290(.a(G28), .O(gate473inter7));
  inv1  gate2291(.a(G1213), .O(gate473inter8));
  nand2 gate2292(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2293(.a(s_249), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2294(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2295(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2296(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2871(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2872(.a(gate474inter0), .b(s_332), .O(gate474inter1));
  and2  gate2873(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2874(.a(s_332), .O(gate474inter3));
  inv1  gate2875(.a(s_333), .O(gate474inter4));
  nand2 gate2876(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2877(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2878(.a(G1117), .O(gate474inter7));
  inv1  gate2879(.a(G1213), .O(gate474inter8));
  nand2 gate2880(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2881(.a(s_333), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2882(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2883(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2884(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate939(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate940(.a(gate476inter0), .b(s_56), .O(gate476inter1));
  and2  gate941(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate942(.a(s_56), .O(gate476inter3));
  inv1  gate943(.a(s_57), .O(gate476inter4));
  nand2 gate944(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate945(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate946(.a(G1120), .O(gate476inter7));
  inv1  gate947(.a(G1216), .O(gate476inter8));
  nand2 gate948(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate949(.a(s_57), .b(gate476inter3), .O(gate476inter10));
  nor2  gate950(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate951(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate952(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate2003(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2004(.a(gate477inter0), .b(s_208), .O(gate477inter1));
  and2  gate2005(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2006(.a(s_208), .O(gate477inter3));
  inv1  gate2007(.a(s_209), .O(gate477inter4));
  nand2 gate2008(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2009(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2010(.a(G30), .O(gate477inter7));
  inv1  gate2011(.a(G1219), .O(gate477inter8));
  nand2 gate2012(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2013(.a(s_209), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2014(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2015(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2016(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2591(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2592(.a(gate478inter0), .b(s_292), .O(gate478inter1));
  and2  gate2593(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2594(.a(s_292), .O(gate478inter3));
  inv1  gate2595(.a(s_293), .O(gate478inter4));
  nand2 gate2596(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2597(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2598(.a(G1123), .O(gate478inter7));
  inv1  gate2599(.a(G1219), .O(gate478inter8));
  nand2 gate2600(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2601(.a(s_293), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2602(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2603(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2604(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate645(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate646(.a(gate479inter0), .b(s_14), .O(gate479inter1));
  and2  gate647(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate648(.a(s_14), .O(gate479inter3));
  inv1  gate649(.a(s_15), .O(gate479inter4));
  nand2 gate650(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate651(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate652(.a(G31), .O(gate479inter7));
  inv1  gate653(.a(G1222), .O(gate479inter8));
  nand2 gate654(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate655(.a(s_15), .b(gate479inter3), .O(gate479inter10));
  nor2  gate656(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate657(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate658(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1625(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1626(.a(gate480inter0), .b(s_154), .O(gate480inter1));
  and2  gate1627(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1628(.a(s_154), .O(gate480inter3));
  inv1  gate1629(.a(s_155), .O(gate480inter4));
  nand2 gate1630(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1631(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1632(.a(G1126), .O(gate480inter7));
  inv1  gate1633(.a(G1222), .O(gate480inter8));
  nand2 gate1634(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1635(.a(s_155), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1636(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1637(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1638(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate3053(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate3054(.a(gate482inter0), .b(s_358), .O(gate482inter1));
  and2  gate3055(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate3056(.a(s_358), .O(gate482inter3));
  inv1  gate3057(.a(s_359), .O(gate482inter4));
  nand2 gate3058(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate3059(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate3060(.a(G1129), .O(gate482inter7));
  inv1  gate3061(.a(G1225), .O(gate482inter8));
  nand2 gate3062(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate3063(.a(s_359), .b(gate482inter3), .O(gate482inter10));
  nor2  gate3064(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate3065(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate3066(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1779(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1780(.a(gate483inter0), .b(s_176), .O(gate483inter1));
  and2  gate1781(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1782(.a(s_176), .O(gate483inter3));
  inv1  gate1783(.a(s_177), .O(gate483inter4));
  nand2 gate1784(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1785(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1786(.a(G1228), .O(gate483inter7));
  inv1  gate1787(.a(G1229), .O(gate483inter8));
  nand2 gate1788(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1789(.a(s_177), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1790(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1791(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1792(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1681(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1682(.a(gate485inter0), .b(s_162), .O(gate485inter1));
  and2  gate1683(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1684(.a(s_162), .O(gate485inter3));
  inv1  gate1685(.a(s_163), .O(gate485inter4));
  nand2 gate1686(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1687(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1688(.a(G1232), .O(gate485inter7));
  inv1  gate1689(.a(G1233), .O(gate485inter8));
  nand2 gate1690(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1691(.a(s_163), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1692(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1693(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1694(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1709(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1710(.a(gate486inter0), .b(s_166), .O(gate486inter1));
  and2  gate1711(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1712(.a(s_166), .O(gate486inter3));
  inv1  gate1713(.a(s_167), .O(gate486inter4));
  nand2 gate1714(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1715(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1716(.a(G1234), .O(gate486inter7));
  inv1  gate1717(.a(G1235), .O(gate486inter8));
  nand2 gate1718(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1719(.a(s_167), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1720(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1721(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1722(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1667(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1668(.a(gate488inter0), .b(s_160), .O(gate488inter1));
  and2  gate1669(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1670(.a(s_160), .O(gate488inter3));
  inv1  gate1671(.a(s_161), .O(gate488inter4));
  nand2 gate1672(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1673(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1674(.a(G1238), .O(gate488inter7));
  inv1  gate1675(.a(G1239), .O(gate488inter8));
  nand2 gate1676(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1677(.a(s_161), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1678(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1679(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1680(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate2255(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2256(.a(gate489inter0), .b(s_244), .O(gate489inter1));
  and2  gate2257(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2258(.a(s_244), .O(gate489inter3));
  inv1  gate2259(.a(s_245), .O(gate489inter4));
  nand2 gate2260(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2261(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2262(.a(G1240), .O(gate489inter7));
  inv1  gate2263(.a(G1241), .O(gate489inter8));
  nand2 gate2264(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2265(.a(s_245), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2266(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2267(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2268(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate2339(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2340(.a(gate490inter0), .b(s_256), .O(gate490inter1));
  and2  gate2341(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2342(.a(s_256), .O(gate490inter3));
  inv1  gate2343(.a(s_257), .O(gate490inter4));
  nand2 gate2344(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2345(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2346(.a(G1242), .O(gate490inter7));
  inv1  gate2347(.a(G1243), .O(gate490inter8));
  nand2 gate2348(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2349(.a(s_257), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2350(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2351(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2352(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate799(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate800(.a(gate494inter0), .b(s_36), .O(gate494inter1));
  and2  gate801(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate802(.a(s_36), .O(gate494inter3));
  inv1  gate803(.a(s_37), .O(gate494inter4));
  nand2 gate804(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate805(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate806(.a(G1250), .O(gate494inter7));
  inv1  gate807(.a(G1251), .O(gate494inter8));
  nand2 gate808(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate809(.a(s_37), .b(gate494inter3), .O(gate494inter10));
  nor2  gate810(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate811(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate812(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate729(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate730(.a(gate495inter0), .b(s_26), .O(gate495inter1));
  and2  gate731(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate732(.a(s_26), .O(gate495inter3));
  inv1  gate733(.a(s_27), .O(gate495inter4));
  nand2 gate734(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate735(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate736(.a(G1252), .O(gate495inter7));
  inv1  gate737(.a(G1253), .O(gate495inter8));
  nand2 gate738(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate739(.a(s_27), .b(gate495inter3), .O(gate495inter10));
  nor2  gate740(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate741(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate742(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2381(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2382(.a(gate497inter0), .b(s_262), .O(gate497inter1));
  and2  gate2383(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2384(.a(s_262), .O(gate497inter3));
  inv1  gate2385(.a(s_263), .O(gate497inter4));
  nand2 gate2386(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2387(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2388(.a(G1256), .O(gate497inter7));
  inv1  gate2389(.a(G1257), .O(gate497inter8));
  nand2 gate2390(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2391(.a(s_263), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2392(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2393(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2394(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate2129(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2130(.a(gate498inter0), .b(s_226), .O(gate498inter1));
  and2  gate2131(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2132(.a(s_226), .O(gate498inter3));
  inv1  gate2133(.a(s_227), .O(gate498inter4));
  nand2 gate2134(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2135(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2136(.a(G1258), .O(gate498inter7));
  inv1  gate2137(.a(G1259), .O(gate498inter8));
  nand2 gate2138(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2139(.a(s_227), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2140(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2141(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2142(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate897(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate898(.a(gate499inter0), .b(s_50), .O(gate499inter1));
  and2  gate899(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate900(.a(s_50), .O(gate499inter3));
  inv1  gate901(.a(s_51), .O(gate499inter4));
  nand2 gate902(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate903(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate904(.a(G1260), .O(gate499inter7));
  inv1  gate905(.a(G1261), .O(gate499inter8));
  nand2 gate906(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate907(.a(s_51), .b(gate499inter3), .O(gate499inter10));
  nor2  gate908(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate909(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate910(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1387(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1388(.a(gate502inter0), .b(s_120), .O(gate502inter1));
  and2  gate1389(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1390(.a(s_120), .O(gate502inter3));
  inv1  gate1391(.a(s_121), .O(gate502inter4));
  nand2 gate1392(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1393(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1394(.a(G1266), .O(gate502inter7));
  inv1  gate1395(.a(G1267), .O(gate502inter8));
  nand2 gate1396(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1397(.a(s_121), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1398(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1399(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1400(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2017(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2018(.a(gate503inter0), .b(s_210), .O(gate503inter1));
  and2  gate2019(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2020(.a(s_210), .O(gate503inter3));
  inv1  gate2021(.a(s_211), .O(gate503inter4));
  nand2 gate2022(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2023(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2024(.a(G1268), .O(gate503inter7));
  inv1  gate2025(.a(G1269), .O(gate503inter8));
  nand2 gate2026(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2027(.a(s_211), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2028(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2029(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2030(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1037(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1038(.a(gate505inter0), .b(s_70), .O(gate505inter1));
  and2  gate1039(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1040(.a(s_70), .O(gate505inter3));
  inv1  gate1041(.a(s_71), .O(gate505inter4));
  nand2 gate1042(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1043(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1044(.a(G1272), .O(gate505inter7));
  inv1  gate1045(.a(G1273), .O(gate505inter8));
  nand2 gate1046(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1047(.a(s_71), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1048(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1049(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1050(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1695(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1696(.a(gate507inter0), .b(s_164), .O(gate507inter1));
  and2  gate1697(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1698(.a(s_164), .O(gate507inter3));
  inv1  gate1699(.a(s_165), .O(gate507inter4));
  nand2 gate1700(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1701(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1702(.a(G1276), .O(gate507inter7));
  inv1  gate1703(.a(G1277), .O(gate507inter8));
  nand2 gate1704(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1705(.a(s_165), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1706(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1707(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1708(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate953(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate954(.a(gate514inter0), .b(s_58), .O(gate514inter1));
  and2  gate955(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate956(.a(s_58), .O(gate514inter3));
  inv1  gate957(.a(s_59), .O(gate514inter4));
  nand2 gate958(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate959(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate960(.a(G1290), .O(gate514inter7));
  inv1  gate961(.a(G1291), .O(gate514inter8));
  nand2 gate962(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate963(.a(s_59), .b(gate514inter3), .O(gate514inter10));
  nor2  gate964(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate965(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate966(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule