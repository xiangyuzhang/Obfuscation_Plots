module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate609(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate610(.a(gate3inter0), .b(s_58), .O(gate3inter1));
  and2  gate611(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate612(.a(s_58), .O(gate3inter3));
  inv1  gate613(.a(s_59), .O(gate3inter4));
  nand2 gate614(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate615(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate616(.a(N17), .O(gate3inter7));
  inv1  gate617(.a(N21), .O(gate3inter8));
  nand2 gate618(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate619(.a(s_59), .b(gate3inter3), .O(gate3inter10));
  nor2  gate620(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate621(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate622(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );

  xor2  gate413(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate414(.a(gate11inter0), .b(s_30), .O(gate11inter1));
  and2  gate415(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate416(.a(s_30), .O(gate11inter3));
  inv1  gate417(.a(s_31), .O(gate11inter4));
  nand2 gate418(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate419(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate420(.a(N81), .O(gate11inter7));
  inv1  gate421(.a(N85), .O(gate11inter8));
  nand2 gate422(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate423(.a(s_31), .b(gate11inter3), .O(gate11inter10));
  nor2  gate424(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate425(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate426(.a(gate11inter12), .b(gate11inter1), .O(N260));
xor2 gate12( .a(N89), .b(N93), .O(N261) );

  xor2  gate511(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate512(.a(gate13inter0), .b(s_44), .O(gate13inter1));
  and2  gate513(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate514(.a(s_44), .O(gate13inter3));
  inv1  gate515(.a(s_45), .O(gate13inter4));
  nand2 gate516(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate517(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate518(.a(N97), .O(gate13inter7));
  inv1  gate519(.a(N101), .O(gate13inter8));
  nand2 gate520(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate521(.a(s_45), .b(gate13inter3), .O(gate13inter10));
  nor2  gate522(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate523(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate524(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate595(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate596(.a(gate25inter0), .b(s_56), .O(gate25inter1));
  and2  gate597(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate598(.a(s_56), .O(gate25inter3));
  inv1  gate599(.a(s_57), .O(gate25inter4));
  nand2 gate600(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate601(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate602(.a(N1), .O(gate25inter7));
  inv1  gate603(.a(N17), .O(gate25inter8));
  nand2 gate604(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate605(.a(s_57), .b(gate25inter3), .O(gate25inter10));
  nor2  gate606(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate607(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate608(.a(gate25inter12), .b(gate25inter1), .O(N274));
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );

  xor2  gate469(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate470(.a(gate29inter0), .b(s_38), .O(gate29inter1));
  and2  gate471(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate472(.a(s_38), .O(gate29inter3));
  inv1  gate473(.a(s_39), .O(gate29inter4));
  nand2 gate474(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate475(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate476(.a(N9), .O(gate29inter7));
  inv1  gate477(.a(N25), .O(gate29inter8));
  nand2 gate478(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate479(.a(s_39), .b(gate29inter3), .O(gate29inter10));
  nor2  gate480(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate481(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate482(.a(gate29inter12), .b(gate29inter1), .O(N278));
xor2 gate30( .a(N41), .b(N57), .O(N279) );

  xor2  gate357(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate358(.a(gate31inter0), .b(s_22), .O(gate31inter1));
  and2  gate359(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate360(.a(s_22), .O(gate31inter3));
  inv1  gate361(.a(s_23), .O(gate31inter4));
  nand2 gate362(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate363(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate364(.a(N13), .O(gate31inter7));
  inv1  gate365(.a(N29), .O(gate31inter8));
  nand2 gate366(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate367(.a(s_23), .b(gate31inter3), .O(gate31inter10));
  nor2  gate368(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate369(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate370(.a(gate31inter12), .b(gate31inter1), .O(N280));

  xor2  gate567(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate568(.a(gate32inter0), .b(s_52), .O(gate32inter1));
  and2  gate569(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate570(.a(s_52), .O(gate32inter3));
  inv1  gate571(.a(s_53), .O(gate32inter4));
  nand2 gate572(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate573(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate574(.a(N45), .O(gate32inter7));
  inv1  gate575(.a(N61), .O(gate32inter8));
  nand2 gate576(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate577(.a(s_53), .b(gate32inter3), .O(gate32inter10));
  nor2  gate578(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate579(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate580(.a(gate32inter12), .b(gate32inter1), .O(N281));
xor2 gate33( .a(N65), .b(N81), .O(N282) );

  xor2  gate315(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate316(.a(gate34inter0), .b(s_16), .O(gate34inter1));
  and2  gate317(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate318(.a(s_16), .O(gate34inter3));
  inv1  gate319(.a(s_17), .O(gate34inter4));
  nand2 gate320(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate321(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate322(.a(N97), .O(gate34inter7));
  inv1  gate323(.a(N113), .O(gate34inter8));
  nand2 gate324(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate325(.a(s_17), .b(gate34inter3), .O(gate34inter10));
  nor2  gate326(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate327(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate328(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );

  xor2  gate455(.a(N251), .b(N250), .O(gate41inter0));
  nand2 gate456(.a(gate41inter0), .b(s_36), .O(gate41inter1));
  and2  gate457(.a(N251), .b(N250), .O(gate41inter2));
  inv1  gate458(.a(s_36), .O(gate41inter3));
  inv1  gate459(.a(s_37), .O(gate41inter4));
  nand2 gate460(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate461(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate462(.a(N250), .O(gate41inter7));
  inv1  gate463(.a(N251), .O(gate41inter8));
  nand2 gate464(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate465(.a(s_37), .b(gate41inter3), .O(gate41inter10));
  nor2  gate466(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate467(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate468(.a(gate41inter12), .b(gate41inter1), .O(N290));
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );

  xor2  gate245(.a(N257), .b(N256), .O(gate44inter0));
  nand2 gate246(.a(gate44inter0), .b(s_6), .O(gate44inter1));
  and2  gate247(.a(N257), .b(N256), .O(gate44inter2));
  inv1  gate248(.a(s_6), .O(gate44inter3));
  inv1  gate249(.a(s_7), .O(gate44inter4));
  nand2 gate250(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate251(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate252(.a(N256), .O(gate44inter7));
  inv1  gate253(.a(N257), .O(gate44inter8));
  nand2 gate254(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate255(.a(s_7), .b(gate44inter3), .O(gate44inter10));
  nor2  gate256(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate257(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate258(.a(gate44inter12), .b(gate44inter1), .O(N299));

  xor2  gate637(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate638(.a(gate45inter0), .b(s_62), .O(gate45inter1));
  and2  gate639(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate640(.a(s_62), .O(gate45inter3));
  inv1  gate641(.a(s_63), .O(gate45inter4));
  nand2 gate642(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate643(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate644(.a(N258), .O(gate45inter7));
  inv1  gate645(.a(N259), .O(gate45inter8));
  nand2 gate646(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate647(.a(s_63), .b(gate45inter3), .O(gate45inter10));
  nor2  gate648(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate649(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate650(.a(gate45inter12), .b(gate45inter1), .O(N302));

  xor2  gate385(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate386(.a(gate46inter0), .b(s_26), .O(gate46inter1));
  and2  gate387(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate388(.a(s_26), .O(gate46inter3));
  inv1  gate389(.a(s_27), .O(gate46inter4));
  nand2 gate390(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate391(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate392(.a(N260), .O(gate46inter7));
  inv1  gate393(.a(N261), .O(gate46inter8));
  nand2 gate394(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate395(.a(s_27), .b(gate46inter3), .O(gate46inter10));
  nor2  gate396(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate397(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate398(.a(gate46inter12), .b(gate46inter1), .O(N305));
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate203(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate204(.a(gate50inter0), .b(s_0), .O(gate50inter1));
  and2  gate205(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate206(.a(s_0), .O(gate50inter3));
  inv1  gate207(.a(s_1), .O(gate50inter4));
  nand2 gate208(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate209(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate210(.a(N276), .O(gate50inter7));
  inv1  gate211(.a(N277), .O(gate50inter8));
  nand2 gate212(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate213(.a(s_1), .b(gate50inter3), .O(gate50inter10));
  nor2  gate214(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate215(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate216(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );

  xor2  gate371(.a(N281), .b(N280), .O(gate52inter0));
  nand2 gate372(.a(gate52inter0), .b(s_24), .O(gate52inter1));
  and2  gate373(.a(N281), .b(N280), .O(gate52inter2));
  inv1  gate374(.a(s_24), .O(gate52inter3));
  inv1  gate375(.a(s_25), .O(gate52inter4));
  nand2 gate376(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate377(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate378(.a(N280), .O(gate52inter7));
  inv1  gate379(.a(N281), .O(gate52inter8));
  nand2 gate380(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate381(.a(s_25), .b(gate52inter3), .O(gate52inter10));
  nor2  gate382(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate383(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate384(.a(gate52inter12), .b(gate52inter1), .O(N317));
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );

  xor2  gate483(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate484(.a(gate58inter0), .b(s_40), .O(gate58inter1));
  and2  gate485(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate486(.a(s_40), .O(gate58inter3));
  inv1  gate487(.a(s_41), .O(gate58inter4));
  nand2 gate488(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate489(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate490(.a(N296), .O(gate58inter7));
  inv1  gate491(.a(N299), .O(gate58inter8));
  nand2 gate492(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate493(.a(s_41), .b(gate58inter3), .O(gate58inter10));
  nor2  gate494(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate495(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate496(.a(gate58inter12), .b(gate58inter1), .O(N339));
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate623(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate624(.a(gate62inter0), .b(s_60), .O(gate62inter1));
  and2  gate625(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate626(.a(s_60), .O(gate62inter3));
  inv1  gate627(.a(s_61), .O(gate62inter4));
  nand2 gate628(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate629(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate630(.a(N308), .O(gate62inter7));
  inv1  gate631(.a(N311), .O(gate62inter8));
  nand2 gate632(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate633(.a(s_61), .b(gate62inter3), .O(gate62inter10));
  nor2  gate634(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate635(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate636(.a(gate62inter12), .b(gate62inter1), .O(N343));

  xor2  gate651(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate652(.a(gate63inter0), .b(s_64), .O(gate63inter1));
  and2  gate653(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate654(.a(s_64), .O(gate63inter3));
  inv1  gate655(.a(s_65), .O(gate63inter4));
  nand2 gate656(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate657(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate658(.a(N302), .O(gate63inter7));
  inv1  gate659(.a(N308), .O(gate63inter8));
  nand2 gate660(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate661(.a(s_65), .b(gate63inter3), .O(gate63inter10));
  nor2  gate662(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate663(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate664(.a(gate63inter12), .b(gate63inter1), .O(N344));
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate329(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate330(.a(gate65inter0), .b(s_18), .O(gate65inter1));
  and2  gate331(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate332(.a(s_18), .O(gate65inter3));
  inv1  gate333(.a(s_19), .O(gate65inter4));
  nand2 gate334(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate335(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate336(.a(N266), .O(gate65inter7));
  inv1  gate337(.a(N342), .O(gate65inter8));
  nand2 gate338(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate339(.a(s_19), .b(gate65inter3), .O(gate65inter10));
  nor2  gate340(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate341(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate342(.a(gate65inter12), .b(gate65inter1), .O(N346));

  xor2  gate665(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate666(.a(gate66inter0), .b(s_66), .O(gate66inter1));
  and2  gate667(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate668(.a(s_66), .O(gate66inter3));
  inv1  gate669(.a(s_67), .O(gate66inter4));
  nand2 gate670(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate671(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate672(.a(N267), .O(gate66inter7));
  inv1  gate673(.a(N343), .O(gate66inter8));
  nand2 gate674(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate675(.a(s_67), .b(gate66inter3), .O(gate66inter10));
  nor2  gate676(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate677(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate678(.a(gate66inter12), .b(gate66inter1), .O(N347));
xor2 gate67( .a(N268), .b(N344), .O(N348) );

  xor2  gate273(.a(N345), .b(N269), .O(gate68inter0));
  nand2 gate274(.a(gate68inter0), .b(s_10), .O(gate68inter1));
  and2  gate275(.a(N345), .b(N269), .O(gate68inter2));
  inv1  gate276(.a(s_10), .O(gate68inter3));
  inv1  gate277(.a(s_11), .O(gate68inter4));
  nand2 gate278(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate279(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate280(.a(N269), .O(gate68inter7));
  inv1  gate281(.a(N345), .O(gate68inter8));
  nand2 gate282(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate283(.a(s_11), .b(gate68inter3), .O(gate68inter10));
  nor2  gate284(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate285(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate286(.a(gate68inter12), .b(gate68inter1), .O(N349));
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate679(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate680(.a(gate70inter0), .b(s_68), .O(gate70inter1));
  and2  gate681(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate682(.a(s_68), .O(gate70inter3));
  inv1  gate683(.a(s_69), .O(gate70inter4));
  nand2 gate684(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate685(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate686(.a(N271), .O(gate70inter7));
  inv1  gate687(.a(N339), .O(gate70inter8));
  nand2 gate688(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate689(.a(s_69), .b(gate70inter3), .O(gate70inter10));
  nor2  gate690(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate691(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate692(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );

  xor2  gate259(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate260(.a(gate74inter0), .b(s_8), .O(gate74inter1));
  and2  gate261(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate262(.a(s_8), .O(gate74inter3));
  inv1  gate263(.a(s_9), .O(gate74inter4));
  nand2 gate264(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate265(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate266(.a(N315), .O(gate74inter7));
  inv1  gate267(.a(N347), .O(gate74inter8));
  nand2 gate268(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate269(.a(s_9), .b(gate74inter3), .O(gate74inter10));
  nor2  gate270(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate271(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate272(.a(gate74inter12), .b(gate74inter1), .O(N367));

  xor2  gate301(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate302(.a(gate75inter0), .b(s_14), .O(gate75inter1));
  and2  gate303(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate304(.a(s_14), .O(gate75inter3));
  inv1  gate305(.a(s_15), .O(gate75inter4));
  nand2 gate306(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate307(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate308(.a(N316), .O(gate75inter7));
  inv1  gate309(.a(N348), .O(gate75inter8));
  nand2 gate310(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate311(.a(s_15), .b(gate75inter3), .O(gate75inter10));
  nor2  gate312(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate313(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate314(.a(gate75inter12), .b(gate75inter1), .O(N380));

  xor2  gate693(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate694(.a(gate76inter0), .b(s_70), .O(gate76inter1));
  and2  gate695(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate696(.a(s_70), .O(gate76inter3));
  inv1  gate697(.a(s_71), .O(gate76inter4));
  nand2 gate698(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate699(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate700(.a(N317), .O(gate76inter7));
  inv1  gate701(.a(N349), .O(gate76inter8));
  nand2 gate702(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate703(.a(s_71), .b(gate76inter3), .O(gate76inter10));
  nor2  gate704(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate705(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate706(.a(gate76inter12), .b(gate76inter1), .O(N393));
xor2 gate77( .a(N318), .b(N350), .O(N406) );

  xor2  gate581(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate582(.a(gate78inter0), .b(s_54), .O(gate78inter1));
  and2  gate583(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate584(.a(s_54), .O(gate78inter3));
  inv1  gate585(.a(s_55), .O(gate78inter4));
  nand2 gate586(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate587(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate588(.a(N319), .O(gate78inter7));
  inv1  gate589(.a(N351), .O(gate78inter8));
  nand2 gate590(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate591(.a(s_55), .b(gate78inter3), .O(gate78inter10));
  nor2  gate592(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate593(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate594(.a(gate78inter12), .b(gate78inter1), .O(N419));

  xor2  gate553(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate554(.a(gate79inter0), .b(s_50), .O(gate79inter1));
  and2  gate555(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate556(.a(s_50), .O(gate79inter3));
  inv1  gate557(.a(s_51), .O(gate79inter4));
  nand2 gate558(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate559(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate560(.a(N320), .O(gate79inter7));
  inv1  gate561(.a(N352), .O(gate79inter8));
  nand2 gate562(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate563(.a(s_51), .b(gate79inter3), .O(gate79inter10));
  nor2  gate564(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate565(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate566(.a(gate79inter12), .b(gate79inter1), .O(N432));
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate217(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate218(.a(gate172inter0), .b(s_2), .O(gate172inter1));
  and2  gate219(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate220(.a(s_2), .O(gate172inter3));
  inv1  gate221(.a(s_3), .O(gate172inter4));
  nand2 gate222(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate223(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate224(.a(N5), .O(gate172inter7));
  inv1  gate225(.a(N693), .O(gate172inter8));
  nand2 gate226(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate227(.a(s_3), .b(gate172inter3), .O(gate172inter10));
  nor2  gate228(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate229(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate230(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate287(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate288(.a(gate177inter0), .b(s_12), .O(gate177inter1));
  and2  gate289(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate290(.a(s_12), .O(gate177inter3));
  inv1  gate291(.a(s_13), .O(gate177inter4));
  nand2 gate292(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate293(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate294(.a(N25), .O(gate177inter7));
  inv1  gate295(.a(N698), .O(gate177inter8));
  nand2 gate296(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate297(.a(s_13), .b(gate177inter3), .O(gate177inter10));
  nor2  gate298(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate299(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate300(.a(gate177inter12), .b(gate177inter1), .O(N730));
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );

  xor2  gate427(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate428(.a(gate183inter0), .b(s_32), .O(gate183inter1));
  and2  gate429(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate430(.a(s_32), .O(gate183inter3));
  inv1  gate431(.a(s_33), .O(gate183inter4));
  nand2 gate432(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate433(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate434(.a(N49), .O(gate183inter7));
  inv1  gate435(.a(N704), .O(gate183inter8));
  nand2 gate436(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate437(.a(s_33), .b(gate183inter3), .O(gate183inter10));
  nor2  gate438(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate439(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate440(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );

  xor2  gate497(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate498(.a(gate188inter0), .b(s_42), .O(gate188inter1));
  and2  gate499(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate500(.a(s_42), .O(gate188inter3));
  inv1  gate501(.a(s_43), .O(gate188inter4));
  nand2 gate502(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate503(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate504(.a(N69), .O(gate188inter7));
  inv1  gate505(.a(N709), .O(gate188inter8));
  nand2 gate506(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate507(.a(s_43), .b(gate188inter3), .O(gate188inter10));
  nor2  gate508(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate509(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate510(.a(gate188inter12), .b(gate188inter1), .O(N741));

  xor2  gate441(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate442(.a(gate189inter0), .b(s_34), .O(gate189inter1));
  and2  gate443(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate444(.a(s_34), .O(gate189inter3));
  inv1  gate445(.a(s_35), .O(gate189inter4));
  nand2 gate446(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate447(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate448(.a(N73), .O(gate189inter7));
  inv1  gate449(.a(N710), .O(gate189inter8));
  nand2 gate450(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate451(.a(s_35), .b(gate189inter3), .O(gate189inter10));
  nor2  gate452(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate453(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate454(.a(gate189inter12), .b(gate189inter1), .O(N742));
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );

  xor2  gate539(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate540(.a(gate192inter0), .b(s_48), .O(gate192inter1));
  and2  gate541(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate542(.a(s_48), .O(gate192inter3));
  inv1  gate543(.a(s_49), .O(gate192inter4));
  nand2 gate544(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate545(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate546(.a(N85), .O(gate192inter7));
  inv1  gate547(.a(N713), .O(gate192inter8));
  nand2 gate548(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate549(.a(s_49), .b(gate192inter3), .O(gate192inter10));
  nor2  gate550(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate551(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate552(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );

  xor2  gate343(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate344(.a(gate194inter0), .b(s_20), .O(gate194inter1));
  and2  gate345(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate346(.a(s_20), .O(gate194inter3));
  inv1  gate347(.a(s_21), .O(gate194inter4));
  nand2 gate348(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate349(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate350(.a(N93), .O(gate194inter7));
  inv1  gate351(.a(N715), .O(gate194inter8));
  nand2 gate352(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate353(.a(s_21), .b(gate194inter3), .O(gate194inter10));
  nor2  gate354(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate355(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate356(.a(gate194inter12), .b(gate194inter1), .O(N747));

  xor2  gate231(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate232(.a(gate195inter0), .b(s_4), .O(gate195inter1));
  and2  gate233(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate234(.a(s_4), .O(gate195inter3));
  inv1  gate235(.a(s_5), .O(gate195inter4));
  nand2 gate236(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate237(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate238(.a(N97), .O(gate195inter7));
  inv1  gate239(.a(N716), .O(gate195inter8));
  nand2 gate240(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate241(.a(s_5), .b(gate195inter3), .O(gate195inter10));
  nor2  gate242(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate243(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate244(.a(gate195inter12), .b(gate195inter1), .O(N748));
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate525(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate526(.a(gate201inter0), .b(s_46), .O(gate201inter1));
  and2  gate527(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate528(.a(s_46), .O(gate201inter3));
  inv1  gate529(.a(s_47), .O(gate201inter4));
  nand2 gate530(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate531(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate532(.a(N121), .O(gate201inter7));
  inv1  gate533(.a(N722), .O(gate201inter8));
  nand2 gate534(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate535(.a(s_47), .b(gate201inter3), .O(gate201inter10));
  nor2  gate536(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate537(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate538(.a(gate201inter12), .b(gate201inter1), .O(N754));

  xor2  gate399(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate400(.a(gate202inter0), .b(s_28), .O(gate202inter1));
  and2  gate401(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate402(.a(s_28), .O(gate202inter3));
  inv1  gate403(.a(s_29), .O(gate202inter4));
  nand2 gate404(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate405(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate406(.a(N125), .O(gate202inter7));
  inv1  gate407(.a(N723), .O(gate202inter8));
  nand2 gate408(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate409(.a(s_29), .b(gate202inter3), .O(gate202inter10));
  nor2  gate410(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate411(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate412(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule