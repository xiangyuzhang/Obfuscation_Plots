module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1415(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1416(.a(gate10inter0), .b(s_124), .O(gate10inter1));
  and2  gate1417(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1418(.a(s_124), .O(gate10inter3));
  inv1  gate1419(.a(s_125), .O(gate10inter4));
  nand2 gate1420(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1421(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1422(.a(G3), .O(gate10inter7));
  inv1  gate1423(.a(G4), .O(gate10inter8));
  nand2 gate1424(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1425(.a(s_125), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1426(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1427(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1428(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1373(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1374(.a(gate13inter0), .b(s_118), .O(gate13inter1));
  and2  gate1375(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1376(.a(s_118), .O(gate13inter3));
  inv1  gate1377(.a(s_119), .O(gate13inter4));
  nand2 gate1378(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1379(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1380(.a(G9), .O(gate13inter7));
  inv1  gate1381(.a(G10), .O(gate13inter8));
  nand2 gate1382(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1383(.a(s_119), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1384(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1385(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1386(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1457(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1458(.a(gate15inter0), .b(s_130), .O(gate15inter1));
  and2  gate1459(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1460(.a(s_130), .O(gate15inter3));
  inv1  gate1461(.a(s_131), .O(gate15inter4));
  nand2 gate1462(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1463(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1464(.a(G13), .O(gate15inter7));
  inv1  gate1465(.a(G14), .O(gate15inter8));
  nand2 gate1466(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1467(.a(s_131), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1468(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1469(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1470(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1835(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1836(.a(gate18inter0), .b(s_184), .O(gate18inter1));
  and2  gate1837(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1838(.a(s_184), .O(gate18inter3));
  inv1  gate1839(.a(s_185), .O(gate18inter4));
  nand2 gate1840(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1841(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1842(.a(G19), .O(gate18inter7));
  inv1  gate1843(.a(G20), .O(gate18inter8));
  nand2 gate1844(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1845(.a(s_185), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1846(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1847(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1848(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate869(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate870(.a(gate19inter0), .b(s_46), .O(gate19inter1));
  and2  gate871(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate872(.a(s_46), .O(gate19inter3));
  inv1  gate873(.a(s_47), .O(gate19inter4));
  nand2 gate874(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate875(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate876(.a(G21), .O(gate19inter7));
  inv1  gate877(.a(G22), .O(gate19inter8));
  nand2 gate878(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate879(.a(s_47), .b(gate19inter3), .O(gate19inter10));
  nor2  gate880(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate881(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate882(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1919(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1920(.a(gate35inter0), .b(s_196), .O(gate35inter1));
  and2  gate1921(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1922(.a(s_196), .O(gate35inter3));
  inv1  gate1923(.a(s_197), .O(gate35inter4));
  nand2 gate1924(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1925(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1926(.a(G18), .O(gate35inter7));
  inv1  gate1927(.a(G22), .O(gate35inter8));
  nand2 gate1928(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1929(.a(s_197), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1930(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1931(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1932(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate827(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate828(.a(gate37inter0), .b(s_40), .O(gate37inter1));
  and2  gate829(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate830(.a(s_40), .O(gate37inter3));
  inv1  gate831(.a(s_41), .O(gate37inter4));
  nand2 gate832(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate833(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate834(.a(G19), .O(gate37inter7));
  inv1  gate835(.a(G23), .O(gate37inter8));
  nand2 gate836(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate837(.a(s_41), .b(gate37inter3), .O(gate37inter10));
  nor2  gate838(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate839(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate840(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1317(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1318(.a(gate38inter0), .b(s_110), .O(gate38inter1));
  and2  gate1319(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1320(.a(s_110), .O(gate38inter3));
  inv1  gate1321(.a(s_111), .O(gate38inter4));
  nand2 gate1322(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1323(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1324(.a(G27), .O(gate38inter7));
  inv1  gate1325(.a(G31), .O(gate38inter8));
  nand2 gate1326(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1327(.a(s_111), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1328(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1329(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1330(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1023(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1024(.a(gate42inter0), .b(s_68), .O(gate42inter1));
  and2  gate1025(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1026(.a(s_68), .O(gate42inter3));
  inv1  gate1027(.a(s_69), .O(gate42inter4));
  nand2 gate1028(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1029(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1030(.a(G2), .O(gate42inter7));
  inv1  gate1031(.a(G266), .O(gate42inter8));
  nand2 gate1032(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1033(.a(s_69), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1034(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1035(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1036(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1639(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1640(.a(gate46inter0), .b(s_156), .O(gate46inter1));
  and2  gate1641(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1642(.a(s_156), .O(gate46inter3));
  inv1  gate1643(.a(s_157), .O(gate46inter4));
  nand2 gate1644(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1645(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1646(.a(G6), .O(gate46inter7));
  inv1  gate1647(.a(G272), .O(gate46inter8));
  nand2 gate1648(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1649(.a(s_157), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1650(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1651(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1652(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1331(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1332(.a(gate47inter0), .b(s_112), .O(gate47inter1));
  and2  gate1333(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1334(.a(s_112), .O(gate47inter3));
  inv1  gate1335(.a(s_113), .O(gate47inter4));
  nand2 gate1336(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1337(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1338(.a(G7), .O(gate47inter7));
  inv1  gate1339(.a(G275), .O(gate47inter8));
  nand2 gate1340(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1341(.a(s_113), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1342(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1343(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1344(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2157(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2158(.a(gate48inter0), .b(s_230), .O(gate48inter1));
  and2  gate2159(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2160(.a(s_230), .O(gate48inter3));
  inv1  gate2161(.a(s_231), .O(gate48inter4));
  nand2 gate2162(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2163(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2164(.a(G8), .O(gate48inter7));
  inv1  gate2165(.a(G275), .O(gate48inter8));
  nand2 gate2166(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2167(.a(s_231), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2168(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2169(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2170(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1569(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1570(.a(gate61inter0), .b(s_146), .O(gate61inter1));
  and2  gate1571(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1572(.a(s_146), .O(gate61inter3));
  inv1  gate1573(.a(s_147), .O(gate61inter4));
  nand2 gate1574(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1575(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1576(.a(G21), .O(gate61inter7));
  inv1  gate1577(.a(G296), .O(gate61inter8));
  nand2 gate1578(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1579(.a(s_147), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1580(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1581(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1582(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1961(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1962(.a(gate71inter0), .b(s_202), .O(gate71inter1));
  and2  gate1963(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1964(.a(s_202), .O(gate71inter3));
  inv1  gate1965(.a(s_203), .O(gate71inter4));
  nand2 gate1966(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1967(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1968(.a(G31), .O(gate71inter7));
  inv1  gate1969(.a(G311), .O(gate71inter8));
  nand2 gate1970(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1971(.a(s_203), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1972(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1973(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1974(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1513(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1514(.a(gate73inter0), .b(s_138), .O(gate73inter1));
  and2  gate1515(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1516(.a(s_138), .O(gate73inter3));
  inv1  gate1517(.a(s_139), .O(gate73inter4));
  nand2 gate1518(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1519(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1520(.a(G1), .O(gate73inter7));
  inv1  gate1521(.a(G314), .O(gate73inter8));
  nand2 gate1522(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1523(.a(s_139), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1524(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1525(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1526(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1037(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1038(.a(gate82inter0), .b(s_70), .O(gate82inter1));
  and2  gate1039(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1040(.a(s_70), .O(gate82inter3));
  inv1  gate1041(.a(s_71), .O(gate82inter4));
  nand2 gate1042(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1043(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1044(.a(G7), .O(gate82inter7));
  inv1  gate1045(.a(G326), .O(gate82inter8));
  nand2 gate1046(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1047(.a(s_71), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1048(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1049(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1050(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1583(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1584(.a(gate83inter0), .b(s_148), .O(gate83inter1));
  and2  gate1585(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1586(.a(s_148), .O(gate83inter3));
  inv1  gate1587(.a(s_149), .O(gate83inter4));
  nand2 gate1588(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1589(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1590(.a(G11), .O(gate83inter7));
  inv1  gate1591(.a(G329), .O(gate83inter8));
  nand2 gate1592(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1593(.a(s_149), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1594(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1595(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1596(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate1891(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1892(.a(gate84inter0), .b(s_192), .O(gate84inter1));
  and2  gate1893(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1894(.a(s_192), .O(gate84inter3));
  inv1  gate1895(.a(s_193), .O(gate84inter4));
  nand2 gate1896(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1897(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1898(.a(G15), .O(gate84inter7));
  inv1  gate1899(.a(G329), .O(gate84inter8));
  nand2 gate1900(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1901(.a(s_193), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1902(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1903(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1904(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate561(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate562(.a(gate88inter0), .b(s_2), .O(gate88inter1));
  and2  gate563(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate564(.a(s_2), .O(gate88inter3));
  inv1  gate565(.a(s_3), .O(gate88inter4));
  nand2 gate566(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate567(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate568(.a(G16), .O(gate88inter7));
  inv1  gate569(.a(G335), .O(gate88inter8));
  nand2 gate570(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate571(.a(s_3), .b(gate88inter3), .O(gate88inter10));
  nor2  gate572(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate573(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate574(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1751(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1752(.a(gate93inter0), .b(s_172), .O(gate93inter1));
  and2  gate1753(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1754(.a(s_172), .O(gate93inter3));
  inv1  gate1755(.a(s_173), .O(gate93inter4));
  nand2 gate1756(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1757(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1758(.a(G18), .O(gate93inter7));
  inv1  gate1759(.a(G344), .O(gate93inter8));
  nand2 gate1760(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1761(.a(s_173), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1762(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1763(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1764(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2115(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2116(.a(gate95inter0), .b(s_224), .O(gate95inter1));
  and2  gate2117(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2118(.a(s_224), .O(gate95inter3));
  inv1  gate2119(.a(s_225), .O(gate95inter4));
  nand2 gate2120(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2121(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2122(.a(G26), .O(gate95inter7));
  inv1  gate2123(.a(G347), .O(gate95inter8));
  nand2 gate2124(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2125(.a(s_225), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2126(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2127(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2128(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate883(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate884(.a(gate96inter0), .b(s_48), .O(gate96inter1));
  and2  gate885(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate886(.a(s_48), .O(gate96inter3));
  inv1  gate887(.a(s_49), .O(gate96inter4));
  nand2 gate888(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate889(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate890(.a(G30), .O(gate96inter7));
  inv1  gate891(.a(G347), .O(gate96inter8));
  nand2 gate892(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate893(.a(s_49), .b(gate96inter3), .O(gate96inter10));
  nor2  gate894(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate895(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate896(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1989(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1990(.a(gate97inter0), .b(s_206), .O(gate97inter1));
  and2  gate1991(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1992(.a(s_206), .O(gate97inter3));
  inv1  gate1993(.a(s_207), .O(gate97inter4));
  nand2 gate1994(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1995(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1996(.a(G19), .O(gate97inter7));
  inv1  gate1997(.a(G350), .O(gate97inter8));
  nand2 gate1998(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1999(.a(s_207), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2000(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2001(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2002(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1709(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1710(.a(gate100inter0), .b(s_166), .O(gate100inter1));
  and2  gate1711(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1712(.a(s_166), .O(gate100inter3));
  inv1  gate1713(.a(s_167), .O(gate100inter4));
  nand2 gate1714(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1715(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1716(.a(G31), .O(gate100inter7));
  inv1  gate1717(.a(G353), .O(gate100inter8));
  nand2 gate1718(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1719(.a(s_167), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1720(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1721(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1722(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2283(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2284(.a(gate102inter0), .b(s_248), .O(gate102inter1));
  and2  gate2285(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2286(.a(s_248), .O(gate102inter3));
  inv1  gate2287(.a(s_249), .O(gate102inter4));
  nand2 gate2288(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2289(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2290(.a(G24), .O(gate102inter7));
  inv1  gate2291(.a(G356), .O(gate102inter8));
  nand2 gate2292(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2293(.a(s_249), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2294(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2295(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2296(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate2227(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2228(.a(gate103inter0), .b(s_240), .O(gate103inter1));
  and2  gate2229(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2230(.a(s_240), .O(gate103inter3));
  inv1  gate2231(.a(s_241), .O(gate103inter4));
  nand2 gate2232(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2233(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2234(.a(G28), .O(gate103inter7));
  inv1  gate2235(.a(G359), .O(gate103inter8));
  nand2 gate2236(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2237(.a(s_241), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2238(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2239(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2240(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate687(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate688(.a(gate104inter0), .b(s_20), .O(gate104inter1));
  and2  gate689(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate690(.a(s_20), .O(gate104inter3));
  inv1  gate691(.a(s_21), .O(gate104inter4));
  nand2 gate692(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate693(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate694(.a(G32), .O(gate104inter7));
  inv1  gate695(.a(G359), .O(gate104inter8));
  nand2 gate696(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate697(.a(s_21), .b(gate104inter3), .O(gate104inter10));
  nor2  gate698(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate699(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate700(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate757(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate758(.a(gate105inter0), .b(s_30), .O(gate105inter1));
  and2  gate759(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate760(.a(s_30), .O(gate105inter3));
  inv1  gate761(.a(s_31), .O(gate105inter4));
  nand2 gate762(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate763(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate764(.a(G362), .O(gate105inter7));
  inv1  gate765(.a(G363), .O(gate105inter8));
  nand2 gate766(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate767(.a(s_31), .b(gate105inter3), .O(gate105inter10));
  nor2  gate768(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate769(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate770(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate673(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate674(.a(gate106inter0), .b(s_18), .O(gate106inter1));
  and2  gate675(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate676(.a(s_18), .O(gate106inter3));
  inv1  gate677(.a(s_19), .O(gate106inter4));
  nand2 gate678(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate679(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate680(.a(G364), .O(gate106inter7));
  inv1  gate681(.a(G365), .O(gate106inter8));
  nand2 gate682(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate683(.a(s_19), .b(gate106inter3), .O(gate106inter10));
  nor2  gate684(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate685(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate686(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate575(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate576(.a(gate109inter0), .b(s_4), .O(gate109inter1));
  and2  gate577(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate578(.a(s_4), .O(gate109inter3));
  inv1  gate579(.a(s_5), .O(gate109inter4));
  nand2 gate580(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate581(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate582(.a(G370), .O(gate109inter7));
  inv1  gate583(.a(G371), .O(gate109inter8));
  nand2 gate584(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate585(.a(s_5), .b(gate109inter3), .O(gate109inter10));
  nor2  gate586(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate587(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate588(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1653(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1654(.a(gate110inter0), .b(s_158), .O(gate110inter1));
  and2  gate1655(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1656(.a(s_158), .O(gate110inter3));
  inv1  gate1657(.a(s_159), .O(gate110inter4));
  nand2 gate1658(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1659(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1660(.a(G372), .O(gate110inter7));
  inv1  gate1661(.a(G373), .O(gate110inter8));
  nand2 gate1662(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1663(.a(s_159), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1664(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1665(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1666(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1527(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1528(.a(gate114inter0), .b(s_140), .O(gate114inter1));
  and2  gate1529(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1530(.a(s_140), .O(gate114inter3));
  inv1  gate1531(.a(s_141), .O(gate114inter4));
  nand2 gate1532(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1533(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1534(.a(G380), .O(gate114inter7));
  inv1  gate1535(.a(G381), .O(gate114inter8));
  nand2 gate1536(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1537(.a(s_141), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1538(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1539(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1540(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate2045(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2046(.a(gate115inter0), .b(s_214), .O(gate115inter1));
  and2  gate2047(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2048(.a(s_214), .O(gate115inter3));
  inv1  gate2049(.a(s_215), .O(gate115inter4));
  nand2 gate2050(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2051(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2052(.a(G382), .O(gate115inter7));
  inv1  gate2053(.a(G383), .O(gate115inter8));
  nand2 gate2054(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2055(.a(s_215), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2056(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2057(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2058(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1359(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1360(.a(gate116inter0), .b(s_116), .O(gate116inter1));
  and2  gate1361(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1362(.a(s_116), .O(gate116inter3));
  inv1  gate1363(.a(s_117), .O(gate116inter4));
  nand2 gate1364(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1365(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1366(.a(G384), .O(gate116inter7));
  inv1  gate1367(.a(G385), .O(gate116inter8));
  nand2 gate1368(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1369(.a(s_117), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1370(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1371(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1372(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate701(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate702(.a(gate118inter0), .b(s_22), .O(gate118inter1));
  and2  gate703(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate704(.a(s_22), .O(gate118inter3));
  inv1  gate705(.a(s_23), .O(gate118inter4));
  nand2 gate706(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate707(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate708(.a(G388), .O(gate118inter7));
  inv1  gate709(.a(G389), .O(gate118inter8));
  nand2 gate710(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate711(.a(s_23), .b(gate118inter3), .O(gate118inter10));
  nor2  gate712(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate713(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate714(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1387(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1388(.a(gate119inter0), .b(s_120), .O(gate119inter1));
  and2  gate1389(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1390(.a(s_120), .O(gate119inter3));
  inv1  gate1391(.a(s_121), .O(gate119inter4));
  nand2 gate1392(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1393(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1394(.a(G390), .O(gate119inter7));
  inv1  gate1395(.a(G391), .O(gate119inter8));
  nand2 gate1396(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1397(.a(s_121), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1398(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1399(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1400(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1863(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1864(.a(gate120inter0), .b(s_188), .O(gate120inter1));
  and2  gate1865(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1866(.a(s_188), .O(gate120inter3));
  inv1  gate1867(.a(s_189), .O(gate120inter4));
  nand2 gate1868(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1869(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1870(.a(G392), .O(gate120inter7));
  inv1  gate1871(.a(G393), .O(gate120inter8));
  nand2 gate1872(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1873(.a(s_189), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1874(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1875(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1876(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1849(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1850(.a(gate127inter0), .b(s_186), .O(gate127inter1));
  and2  gate1851(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1852(.a(s_186), .O(gate127inter3));
  inv1  gate1853(.a(s_187), .O(gate127inter4));
  nand2 gate1854(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1855(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1856(.a(G406), .O(gate127inter7));
  inv1  gate1857(.a(G407), .O(gate127inter8));
  nand2 gate1858(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1859(.a(s_187), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1860(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1861(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1862(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate729(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate730(.a(gate131inter0), .b(s_26), .O(gate131inter1));
  and2  gate731(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate732(.a(s_26), .O(gate131inter3));
  inv1  gate733(.a(s_27), .O(gate131inter4));
  nand2 gate734(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate735(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate736(.a(G414), .O(gate131inter7));
  inv1  gate737(.a(G415), .O(gate131inter8));
  nand2 gate738(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate739(.a(s_27), .b(gate131inter3), .O(gate131inter10));
  nor2  gate740(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate741(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate742(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate659(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate660(.a(gate134inter0), .b(s_16), .O(gate134inter1));
  and2  gate661(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate662(.a(s_16), .O(gate134inter3));
  inv1  gate663(.a(s_17), .O(gate134inter4));
  nand2 gate664(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate665(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate666(.a(G420), .O(gate134inter7));
  inv1  gate667(.a(G421), .O(gate134inter8));
  nand2 gate668(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate669(.a(s_17), .b(gate134inter3), .O(gate134inter10));
  nor2  gate670(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate671(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate672(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1681(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1682(.a(gate136inter0), .b(s_162), .O(gate136inter1));
  and2  gate1683(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1684(.a(s_162), .O(gate136inter3));
  inv1  gate1685(.a(s_163), .O(gate136inter4));
  nand2 gate1686(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1687(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1688(.a(G424), .O(gate136inter7));
  inv1  gate1689(.a(G425), .O(gate136inter8));
  nand2 gate1690(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1691(.a(s_163), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1692(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1693(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1694(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2255(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2256(.a(gate137inter0), .b(s_244), .O(gate137inter1));
  and2  gate2257(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2258(.a(s_244), .O(gate137inter3));
  inv1  gate2259(.a(s_245), .O(gate137inter4));
  nand2 gate2260(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2261(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2262(.a(G426), .O(gate137inter7));
  inv1  gate2263(.a(G429), .O(gate137inter8));
  nand2 gate2264(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2265(.a(s_245), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2266(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2267(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2268(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1345(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1346(.a(gate140inter0), .b(s_114), .O(gate140inter1));
  and2  gate1347(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1348(.a(s_114), .O(gate140inter3));
  inv1  gate1349(.a(s_115), .O(gate140inter4));
  nand2 gate1350(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1351(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1352(.a(G444), .O(gate140inter7));
  inv1  gate1353(.a(G447), .O(gate140inter8));
  nand2 gate1354(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1355(.a(s_115), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1356(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1357(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1358(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1471(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1472(.a(gate141inter0), .b(s_132), .O(gate141inter1));
  and2  gate1473(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1474(.a(s_132), .O(gate141inter3));
  inv1  gate1475(.a(s_133), .O(gate141inter4));
  nand2 gate1476(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1477(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1478(.a(G450), .O(gate141inter7));
  inv1  gate1479(.a(G453), .O(gate141inter8));
  nand2 gate1480(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1481(.a(s_133), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1482(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1483(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1484(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate855(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate856(.a(gate145inter0), .b(s_44), .O(gate145inter1));
  and2  gate857(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate858(.a(s_44), .O(gate145inter3));
  inv1  gate859(.a(s_45), .O(gate145inter4));
  nand2 gate860(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate861(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate862(.a(G474), .O(gate145inter7));
  inv1  gate863(.a(G477), .O(gate145inter8));
  nand2 gate864(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate865(.a(s_45), .b(gate145inter3), .O(gate145inter10));
  nor2  gate866(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate867(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate868(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1541(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1542(.a(gate147inter0), .b(s_142), .O(gate147inter1));
  and2  gate1543(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1544(.a(s_142), .O(gate147inter3));
  inv1  gate1545(.a(s_143), .O(gate147inter4));
  nand2 gate1546(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1547(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1548(.a(G486), .O(gate147inter7));
  inv1  gate1549(.a(G489), .O(gate147inter8));
  nand2 gate1550(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1551(.a(s_143), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1552(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1553(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1554(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1975(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1976(.a(gate152inter0), .b(s_204), .O(gate152inter1));
  and2  gate1977(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1978(.a(s_204), .O(gate152inter3));
  inv1  gate1979(.a(s_205), .O(gate152inter4));
  nand2 gate1980(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1981(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1982(.a(G516), .O(gate152inter7));
  inv1  gate1983(.a(G519), .O(gate152inter8));
  nand2 gate1984(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1985(.a(s_205), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1986(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1987(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1988(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2129(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2130(.a(gate154inter0), .b(s_226), .O(gate154inter1));
  and2  gate2131(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2132(.a(s_226), .O(gate154inter3));
  inv1  gate2133(.a(s_227), .O(gate154inter4));
  nand2 gate2134(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2135(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2136(.a(G429), .O(gate154inter7));
  inv1  gate2137(.a(G522), .O(gate154inter8));
  nand2 gate2138(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2139(.a(s_227), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2140(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2141(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2142(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1807(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1808(.a(gate156inter0), .b(s_180), .O(gate156inter1));
  and2  gate1809(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1810(.a(s_180), .O(gate156inter3));
  inv1  gate1811(.a(s_181), .O(gate156inter4));
  nand2 gate1812(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1813(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1814(.a(G435), .O(gate156inter7));
  inv1  gate1815(.a(G525), .O(gate156inter8));
  nand2 gate1816(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1817(.a(s_181), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1818(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1819(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1820(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2143(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2144(.a(gate157inter0), .b(s_228), .O(gate157inter1));
  and2  gate2145(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2146(.a(s_228), .O(gate157inter3));
  inv1  gate2147(.a(s_229), .O(gate157inter4));
  nand2 gate2148(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2149(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2150(.a(G438), .O(gate157inter7));
  inv1  gate2151(.a(G528), .O(gate157inter8));
  nand2 gate2152(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2153(.a(s_229), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2154(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2155(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2156(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate771(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate772(.a(gate159inter0), .b(s_32), .O(gate159inter1));
  and2  gate773(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate774(.a(s_32), .O(gate159inter3));
  inv1  gate775(.a(s_33), .O(gate159inter4));
  nand2 gate776(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate777(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate778(.a(G444), .O(gate159inter7));
  inv1  gate779(.a(G531), .O(gate159inter8));
  nand2 gate780(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate781(.a(s_33), .b(gate159inter3), .O(gate159inter10));
  nor2  gate782(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate783(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate784(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1163(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1164(.a(gate162inter0), .b(s_88), .O(gate162inter1));
  and2  gate1165(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1166(.a(s_88), .O(gate162inter3));
  inv1  gate1167(.a(s_89), .O(gate162inter4));
  nand2 gate1168(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1169(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1170(.a(G453), .O(gate162inter7));
  inv1  gate1171(.a(G534), .O(gate162inter8));
  nand2 gate1172(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1173(.a(s_89), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1174(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1175(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1176(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1107(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1108(.a(gate167inter0), .b(s_80), .O(gate167inter1));
  and2  gate1109(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1110(.a(s_80), .O(gate167inter3));
  inv1  gate1111(.a(s_81), .O(gate167inter4));
  nand2 gate1112(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1113(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1114(.a(G468), .O(gate167inter7));
  inv1  gate1115(.a(G543), .O(gate167inter8));
  nand2 gate1116(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1117(.a(s_81), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1118(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1119(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1120(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate743(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate744(.a(gate168inter0), .b(s_28), .O(gate168inter1));
  and2  gate745(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate746(.a(s_28), .O(gate168inter3));
  inv1  gate747(.a(s_29), .O(gate168inter4));
  nand2 gate748(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate749(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate750(.a(G471), .O(gate168inter7));
  inv1  gate751(.a(G543), .O(gate168inter8));
  nand2 gate752(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate753(.a(s_29), .b(gate168inter3), .O(gate168inter10));
  nor2  gate754(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate755(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate756(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1191(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1192(.a(gate170inter0), .b(s_92), .O(gate170inter1));
  and2  gate1193(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1194(.a(s_92), .O(gate170inter3));
  inv1  gate1195(.a(s_93), .O(gate170inter4));
  nand2 gate1196(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1197(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1198(.a(G477), .O(gate170inter7));
  inv1  gate1199(.a(G546), .O(gate170inter8));
  nand2 gate1200(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1201(.a(s_93), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1202(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1203(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1204(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2087(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2088(.a(gate181inter0), .b(s_220), .O(gate181inter1));
  and2  gate2089(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2090(.a(s_220), .O(gate181inter3));
  inv1  gate2091(.a(s_221), .O(gate181inter4));
  nand2 gate2092(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2093(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2094(.a(G510), .O(gate181inter7));
  inv1  gate2095(.a(G564), .O(gate181inter8));
  nand2 gate2096(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2097(.a(s_221), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2098(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2099(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2100(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2269(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2270(.a(gate183inter0), .b(s_246), .O(gate183inter1));
  and2  gate2271(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2272(.a(s_246), .O(gate183inter3));
  inv1  gate2273(.a(s_247), .O(gate183inter4));
  nand2 gate2274(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2275(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2276(.a(G516), .O(gate183inter7));
  inv1  gate2277(.a(G567), .O(gate183inter8));
  nand2 gate2278(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2279(.a(s_247), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2280(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2281(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2282(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2101(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2102(.a(gate185inter0), .b(s_222), .O(gate185inter1));
  and2  gate2103(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2104(.a(s_222), .O(gate185inter3));
  inv1  gate2105(.a(s_223), .O(gate185inter4));
  nand2 gate2106(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2107(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2108(.a(G570), .O(gate185inter7));
  inv1  gate2109(.a(G571), .O(gate185inter8));
  nand2 gate2110(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2111(.a(s_223), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2112(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2113(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2114(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate925(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate926(.a(gate188inter0), .b(s_54), .O(gate188inter1));
  and2  gate927(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate928(.a(s_54), .O(gate188inter3));
  inv1  gate929(.a(s_55), .O(gate188inter4));
  nand2 gate930(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate931(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate932(.a(G576), .O(gate188inter7));
  inv1  gate933(.a(G577), .O(gate188inter8));
  nand2 gate934(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate935(.a(s_55), .b(gate188inter3), .O(gate188inter10));
  nor2  gate936(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate937(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate938(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1737(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1738(.a(gate190inter0), .b(s_170), .O(gate190inter1));
  and2  gate1739(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1740(.a(s_170), .O(gate190inter3));
  inv1  gate1741(.a(s_171), .O(gate190inter4));
  nand2 gate1742(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1743(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1744(.a(G580), .O(gate190inter7));
  inv1  gate1745(.a(G581), .O(gate190inter8));
  nand2 gate1746(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1747(.a(s_171), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1748(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1749(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1750(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate939(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate940(.a(gate195inter0), .b(s_56), .O(gate195inter1));
  and2  gate941(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate942(.a(s_56), .O(gate195inter3));
  inv1  gate943(.a(s_57), .O(gate195inter4));
  nand2 gate944(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate945(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate946(.a(G590), .O(gate195inter7));
  inv1  gate947(.a(G591), .O(gate195inter8));
  nand2 gate948(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate949(.a(s_57), .b(gate195inter3), .O(gate195inter10));
  nor2  gate950(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate951(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate952(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate953(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate954(.a(gate197inter0), .b(s_58), .O(gate197inter1));
  and2  gate955(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate956(.a(s_58), .O(gate197inter3));
  inv1  gate957(.a(s_59), .O(gate197inter4));
  nand2 gate958(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate959(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate960(.a(G594), .O(gate197inter7));
  inv1  gate961(.a(G595), .O(gate197inter8));
  nand2 gate962(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate963(.a(s_59), .b(gate197inter3), .O(gate197inter10));
  nor2  gate964(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate965(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate966(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1219(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1220(.a(gate199inter0), .b(s_96), .O(gate199inter1));
  and2  gate1221(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1222(.a(s_96), .O(gate199inter3));
  inv1  gate1223(.a(s_97), .O(gate199inter4));
  nand2 gate1224(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1225(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1226(.a(G598), .O(gate199inter7));
  inv1  gate1227(.a(G599), .O(gate199inter8));
  nand2 gate1228(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1229(.a(s_97), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1230(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1231(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1232(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate785(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate786(.a(gate201inter0), .b(s_34), .O(gate201inter1));
  and2  gate787(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate788(.a(s_34), .O(gate201inter3));
  inv1  gate789(.a(s_35), .O(gate201inter4));
  nand2 gate790(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate791(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate792(.a(G602), .O(gate201inter7));
  inv1  gate793(.a(G607), .O(gate201inter8));
  nand2 gate794(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate795(.a(s_35), .b(gate201inter3), .O(gate201inter10));
  nor2  gate796(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate797(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate798(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1093(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1094(.a(gate202inter0), .b(s_78), .O(gate202inter1));
  and2  gate1095(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1096(.a(s_78), .O(gate202inter3));
  inv1  gate1097(.a(s_79), .O(gate202inter4));
  nand2 gate1098(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1099(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1100(.a(G612), .O(gate202inter7));
  inv1  gate1101(.a(G617), .O(gate202inter8));
  nand2 gate1102(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1103(.a(s_79), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1104(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1105(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1106(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate617(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate618(.a(gate207inter0), .b(s_10), .O(gate207inter1));
  and2  gate619(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate620(.a(s_10), .O(gate207inter3));
  inv1  gate621(.a(s_11), .O(gate207inter4));
  nand2 gate622(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate623(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate624(.a(G622), .O(gate207inter7));
  inv1  gate625(.a(G632), .O(gate207inter8));
  nand2 gate626(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate627(.a(s_11), .b(gate207inter3), .O(gate207inter10));
  nor2  gate628(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate629(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate630(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1905(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1906(.a(gate211inter0), .b(s_194), .O(gate211inter1));
  and2  gate1907(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1908(.a(s_194), .O(gate211inter3));
  inv1  gate1909(.a(s_195), .O(gate211inter4));
  nand2 gate1910(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1911(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1912(.a(G612), .O(gate211inter7));
  inv1  gate1913(.a(G669), .O(gate211inter8));
  nand2 gate1914(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1915(.a(s_195), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1916(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1917(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1918(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2171(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2172(.a(gate212inter0), .b(s_232), .O(gate212inter1));
  and2  gate2173(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2174(.a(s_232), .O(gate212inter3));
  inv1  gate2175(.a(s_233), .O(gate212inter4));
  nand2 gate2176(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2177(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2178(.a(G617), .O(gate212inter7));
  inv1  gate2179(.a(G669), .O(gate212inter8));
  nand2 gate2180(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2181(.a(s_233), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2182(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2183(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2184(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate841(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate842(.a(gate215inter0), .b(s_42), .O(gate215inter1));
  and2  gate843(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate844(.a(s_42), .O(gate215inter3));
  inv1  gate845(.a(s_43), .O(gate215inter4));
  nand2 gate846(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate847(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate848(.a(G607), .O(gate215inter7));
  inv1  gate849(.a(G675), .O(gate215inter8));
  nand2 gate850(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate851(.a(s_43), .b(gate215inter3), .O(gate215inter10));
  nor2  gate852(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate853(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate854(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1933(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1934(.a(gate216inter0), .b(s_198), .O(gate216inter1));
  and2  gate1935(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1936(.a(s_198), .O(gate216inter3));
  inv1  gate1937(.a(s_199), .O(gate216inter4));
  nand2 gate1938(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1939(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1940(.a(G617), .O(gate216inter7));
  inv1  gate1941(.a(G675), .O(gate216inter8));
  nand2 gate1942(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1943(.a(s_199), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1944(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1945(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1946(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1247(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1248(.a(gate221inter0), .b(s_100), .O(gate221inter1));
  and2  gate1249(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1250(.a(s_100), .O(gate221inter3));
  inv1  gate1251(.a(s_101), .O(gate221inter4));
  nand2 gate1252(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1253(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1254(.a(G622), .O(gate221inter7));
  inv1  gate1255(.a(G684), .O(gate221inter8));
  nand2 gate1256(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1257(.a(s_101), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1258(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1259(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1260(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1009(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1010(.a(gate222inter0), .b(s_66), .O(gate222inter1));
  and2  gate1011(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1012(.a(s_66), .O(gate222inter3));
  inv1  gate1013(.a(s_67), .O(gate222inter4));
  nand2 gate1014(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1015(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1016(.a(G632), .O(gate222inter7));
  inv1  gate1017(.a(G684), .O(gate222inter8));
  nand2 gate1018(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1019(.a(s_67), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1020(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1021(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1022(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1177(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1178(.a(gate225inter0), .b(s_90), .O(gate225inter1));
  and2  gate1179(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1180(.a(s_90), .O(gate225inter3));
  inv1  gate1181(.a(s_91), .O(gate225inter4));
  nand2 gate1182(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1183(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1184(.a(G690), .O(gate225inter7));
  inv1  gate1185(.a(G691), .O(gate225inter8));
  nand2 gate1186(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1187(.a(s_91), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1188(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1189(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1190(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2059(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2060(.a(gate229inter0), .b(s_216), .O(gate229inter1));
  and2  gate2061(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2062(.a(s_216), .O(gate229inter3));
  inv1  gate2063(.a(s_217), .O(gate229inter4));
  nand2 gate2064(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2065(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2066(.a(G698), .O(gate229inter7));
  inv1  gate2067(.a(G699), .O(gate229inter8));
  nand2 gate2068(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2069(.a(s_217), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2070(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2071(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2072(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate897(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate898(.a(gate235inter0), .b(s_50), .O(gate235inter1));
  and2  gate899(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate900(.a(s_50), .O(gate235inter3));
  inv1  gate901(.a(s_51), .O(gate235inter4));
  nand2 gate902(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate903(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate904(.a(G248), .O(gate235inter7));
  inv1  gate905(.a(G724), .O(gate235inter8));
  nand2 gate906(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate907(.a(s_51), .b(gate235inter3), .O(gate235inter10));
  nor2  gate908(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate909(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate910(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate799(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate800(.a(gate238inter0), .b(s_36), .O(gate238inter1));
  and2  gate801(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate802(.a(s_36), .O(gate238inter3));
  inv1  gate803(.a(s_37), .O(gate238inter4));
  nand2 gate804(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate805(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate806(.a(G257), .O(gate238inter7));
  inv1  gate807(.a(G709), .O(gate238inter8));
  nand2 gate808(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate809(.a(s_37), .b(gate238inter3), .O(gate238inter10));
  nor2  gate810(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate811(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate812(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate589(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate590(.a(gate240inter0), .b(s_6), .O(gate240inter1));
  and2  gate591(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate592(.a(s_6), .O(gate240inter3));
  inv1  gate593(.a(s_7), .O(gate240inter4));
  nand2 gate594(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate595(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate596(.a(G263), .O(gate240inter7));
  inv1  gate597(.a(G715), .O(gate240inter8));
  nand2 gate598(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate599(.a(s_7), .b(gate240inter3), .O(gate240inter10));
  nor2  gate600(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate601(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate602(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1611(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1612(.a(gate242inter0), .b(s_152), .O(gate242inter1));
  and2  gate1613(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1614(.a(s_152), .O(gate242inter3));
  inv1  gate1615(.a(s_153), .O(gate242inter4));
  nand2 gate1616(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1617(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1618(.a(G718), .O(gate242inter7));
  inv1  gate1619(.a(G730), .O(gate242inter8));
  nand2 gate1620(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1621(.a(s_153), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1622(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1623(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1624(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate967(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate968(.a(gate243inter0), .b(s_60), .O(gate243inter1));
  and2  gate969(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate970(.a(s_60), .O(gate243inter3));
  inv1  gate971(.a(s_61), .O(gate243inter4));
  nand2 gate972(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate973(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate974(.a(G245), .O(gate243inter7));
  inv1  gate975(.a(G733), .O(gate243inter8));
  nand2 gate976(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate977(.a(s_61), .b(gate243inter3), .O(gate243inter10));
  nor2  gate978(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate979(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate980(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1429(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1430(.a(gate245inter0), .b(s_126), .O(gate245inter1));
  and2  gate1431(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1432(.a(s_126), .O(gate245inter3));
  inv1  gate1433(.a(s_127), .O(gate245inter4));
  nand2 gate1434(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1435(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1436(.a(G248), .O(gate245inter7));
  inv1  gate1437(.a(G736), .O(gate245inter8));
  nand2 gate1438(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1439(.a(s_127), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1440(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1441(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1442(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate981(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate982(.a(gate246inter0), .b(s_62), .O(gate246inter1));
  and2  gate983(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate984(.a(s_62), .O(gate246inter3));
  inv1  gate985(.a(s_63), .O(gate246inter4));
  nand2 gate986(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate987(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate988(.a(G724), .O(gate246inter7));
  inv1  gate989(.a(G736), .O(gate246inter8));
  nand2 gate990(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate991(.a(s_63), .b(gate246inter3), .O(gate246inter10));
  nor2  gate992(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate993(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate994(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1065(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1066(.a(gate254inter0), .b(s_74), .O(gate254inter1));
  and2  gate1067(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1068(.a(s_74), .O(gate254inter3));
  inv1  gate1069(.a(s_75), .O(gate254inter4));
  nand2 gate1070(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1071(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1072(.a(G712), .O(gate254inter7));
  inv1  gate1073(.a(G748), .O(gate254inter8));
  nand2 gate1074(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1075(.a(s_75), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1076(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1077(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1078(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1135(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1136(.a(gate258inter0), .b(s_84), .O(gate258inter1));
  and2  gate1137(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1138(.a(s_84), .O(gate258inter3));
  inv1  gate1139(.a(s_85), .O(gate258inter4));
  nand2 gate1140(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1141(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1142(.a(G756), .O(gate258inter7));
  inv1  gate1143(.a(G757), .O(gate258inter8));
  nand2 gate1144(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1145(.a(s_85), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1146(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1147(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1148(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate631(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate632(.a(gate259inter0), .b(s_12), .O(gate259inter1));
  and2  gate633(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate634(.a(s_12), .O(gate259inter3));
  inv1  gate635(.a(s_13), .O(gate259inter4));
  nand2 gate636(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate637(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate638(.a(G758), .O(gate259inter7));
  inv1  gate639(.a(G759), .O(gate259inter8));
  nand2 gate640(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate641(.a(s_13), .b(gate259inter3), .O(gate259inter10));
  nor2  gate642(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate643(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate644(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate911(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate912(.a(gate267inter0), .b(s_52), .O(gate267inter1));
  and2  gate913(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate914(.a(s_52), .O(gate267inter3));
  inv1  gate915(.a(s_53), .O(gate267inter4));
  nand2 gate916(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate917(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate918(.a(G648), .O(gate267inter7));
  inv1  gate919(.a(G776), .O(gate267inter8));
  nand2 gate920(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate921(.a(s_53), .b(gate267inter3), .O(gate267inter10));
  nor2  gate922(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate923(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate924(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2073(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2074(.a(gate268inter0), .b(s_218), .O(gate268inter1));
  and2  gate2075(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2076(.a(s_218), .O(gate268inter3));
  inv1  gate2077(.a(s_219), .O(gate268inter4));
  nand2 gate2078(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2079(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2080(.a(G651), .O(gate268inter7));
  inv1  gate2081(.a(G779), .O(gate268inter8));
  nand2 gate2082(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2083(.a(s_219), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2084(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2085(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2086(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate715(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate716(.a(gate269inter0), .b(s_24), .O(gate269inter1));
  and2  gate717(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate718(.a(s_24), .O(gate269inter3));
  inv1  gate719(.a(s_25), .O(gate269inter4));
  nand2 gate720(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate721(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate722(.a(G654), .O(gate269inter7));
  inv1  gate723(.a(G782), .O(gate269inter8));
  nand2 gate724(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate725(.a(s_25), .b(gate269inter3), .O(gate269inter10));
  nor2  gate726(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate727(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate728(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1443(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1444(.a(gate272inter0), .b(s_128), .O(gate272inter1));
  and2  gate1445(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1446(.a(s_128), .O(gate272inter3));
  inv1  gate1447(.a(s_129), .O(gate272inter4));
  nand2 gate1448(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1449(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1450(.a(G663), .O(gate272inter7));
  inv1  gate1451(.a(G791), .O(gate272inter8));
  nand2 gate1452(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1453(.a(s_129), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1454(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1455(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1456(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2017(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2018(.a(gate275inter0), .b(s_210), .O(gate275inter1));
  and2  gate2019(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2020(.a(s_210), .O(gate275inter3));
  inv1  gate2021(.a(s_211), .O(gate275inter4));
  nand2 gate2022(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2023(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2024(.a(G645), .O(gate275inter7));
  inv1  gate2025(.a(G797), .O(gate275inter8));
  nand2 gate2026(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2027(.a(s_211), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2028(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2029(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2030(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1499(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1500(.a(gate284inter0), .b(s_136), .O(gate284inter1));
  and2  gate1501(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1502(.a(s_136), .O(gate284inter3));
  inv1  gate1503(.a(s_137), .O(gate284inter4));
  nand2 gate1504(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1505(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1506(.a(G785), .O(gate284inter7));
  inv1  gate1507(.a(G809), .O(gate284inter8));
  nand2 gate1508(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1509(.a(s_137), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1510(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1511(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1512(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1261(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1262(.a(gate285inter0), .b(s_102), .O(gate285inter1));
  and2  gate1263(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1264(.a(s_102), .O(gate285inter3));
  inv1  gate1265(.a(s_103), .O(gate285inter4));
  nand2 gate1266(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1267(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1268(.a(G660), .O(gate285inter7));
  inv1  gate1269(.a(G812), .O(gate285inter8));
  nand2 gate1270(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1271(.a(s_103), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1272(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1273(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1274(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1821(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1822(.a(gate287inter0), .b(s_182), .O(gate287inter1));
  and2  gate1823(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1824(.a(s_182), .O(gate287inter3));
  inv1  gate1825(.a(s_183), .O(gate287inter4));
  nand2 gate1826(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1827(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1828(.a(G663), .O(gate287inter7));
  inv1  gate1829(.a(G815), .O(gate287inter8));
  nand2 gate1830(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1831(.a(s_183), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1832(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1833(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1834(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1079(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1080(.a(gate295inter0), .b(s_76), .O(gate295inter1));
  and2  gate1081(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1082(.a(s_76), .O(gate295inter3));
  inv1  gate1083(.a(s_77), .O(gate295inter4));
  nand2 gate1084(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1085(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1086(.a(G830), .O(gate295inter7));
  inv1  gate1087(.a(G831), .O(gate295inter8));
  nand2 gate1088(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1089(.a(s_77), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1090(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1091(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1092(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2031(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2032(.a(gate387inter0), .b(s_212), .O(gate387inter1));
  and2  gate2033(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2034(.a(s_212), .O(gate387inter3));
  inv1  gate2035(.a(s_213), .O(gate387inter4));
  nand2 gate2036(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2037(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2038(.a(G1), .O(gate387inter7));
  inv1  gate2039(.a(G1036), .O(gate387inter8));
  nand2 gate2040(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2041(.a(s_213), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2042(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2043(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2044(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1667(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1668(.a(gate388inter0), .b(s_160), .O(gate388inter1));
  and2  gate1669(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1670(.a(s_160), .O(gate388inter3));
  inv1  gate1671(.a(s_161), .O(gate388inter4));
  nand2 gate1672(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1673(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1674(.a(G2), .O(gate388inter7));
  inv1  gate1675(.a(G1039), .O(gate388inter8));
  nand2 gate1676(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1677(.a(s_161), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1678(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1679(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1680(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1121(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1122(.a(gate389inter0), .b(s_82), .O(gate389inter1));
  and2  gate1123(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1124(.a(s_82), .O(gate389inter3));
  inv1  gate1125(.a(s_83), .O(gate389inter4));
  nand2 gate1126(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1127(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1128(.a(G3), .O(gate389inter7));
  inv1  gate1129(.a(G1042), .O(gate389inter8));
  nand2 gate1130(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1131(.a(s_83), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1132(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1133(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1134(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1625(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1626(.a(gate390inter0), .b(s_154), .O(gate390inter1));
  and2  gate1627(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1628(.a(s_154), .O(gate390inter3));
  inv1  gate1629(.a(s_155), .O(gate390inter4));
  nand2 gate1630(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1631(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1632(.a(G4), .O(gate390inter7));
  inv1  gate1633(.a(G1045), .O(gate390inter8));
  nand2 gate1634(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1635(.a(s_155), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1636(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1637(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1638(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1401(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1402(.a(gate397inter0), .b(s_122), .O(gate397inter1));
  and2  gate1403(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1404(.a(s_122), .O(gate397inter3));
  inv1  gate1405(.a(s_123), .O(gate397inter4));
  nand2 gate1406(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1407(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1408(.a(G11), .O(gate397inter7));
  inv1  gate1409(.a(G1066), .O(gate397inter8));
  nand2 gate1410(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1411(.a(s_123), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1412(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1413(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1414(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1877(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1878(.a(gate399inter0), .b(s_190), .O(gate399inter1));
  and2  gate1879(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1880(.a(s_190), .O(gate399inter3));
  inv1  gate1881(.a(s_191), .O(gate399inter4));
  nand2 gate1882(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1883(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1884(.a(G13), .O(gate399inter7));
  inv1  gate1885(.a(G1072), .O(gate399inter8));
  nand2 gate1886(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1887(.a(s_191), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1888(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1889(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1890(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1149(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1150(.a(gate402inter0), .b(s_86), .O(gate402inter1));
  and2  gate1151(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1152(.a(s_86), .O(gate402inter3));
  inv1  gate1153(.a(s_87), .O(gate402inter4));
  nand2 gate1154(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1155(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1156(.a(G16), .O(gate402inter7));
  inv1  gate1157(.a(G1081), .O(gate402inter8));
  nand2 gate1158(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1159(.a(s_87), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1160(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1161(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1162(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate603(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate604(.a(gate403inter0), .b(s_8), .O(gate403inter1));
  and2  gate605(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate606(.a(s_8), .O(gate403inter3));
  inv1  gate607(.a(s_9), .O(gate403inter4));
  nand2 gate608(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate609(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate610(.a(G17), .O(gate403inter7));
  inv1  gate611(.a(G1084), .O(gate403inter8));
  nand2 gate612(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate613(.a(s_9), .b(gate403inter3), .O(gate403inter10));
  nor2  gate614(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate615(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate616(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1303(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1304(.a(gate404inter0), .b(s_108), .O(gate404inter1));
  and2  gate1305(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1306(.a(s_108), .O(gate404inter3));
  inv1  gate1307(.a(s_109), .O(gate404inter4));
  nand2 gate1308(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1309(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1310(.a(G18), .O(gate404inter7));
  inv1  gate1311(.a(G1087), .O(gate404inter8));
  nand2 gate1312(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1313(.a(s_109), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1314(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1315(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1316(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1723(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1724(.a(gate406inter0), .b(s_168), .O(gate406inter1));
  and2  gate1725(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1726(.a(s_168), .O(gate406inter3));
  inv1  gate1727(.a(s_169), .O(gate406inter4));
  nand2 gate1728(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1729(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1730(.a(G20), .O(gate406inter7));
  inv1  gate1731(.a(G1093), .O(gate406inter8));
  nand2 gate1732(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1733(.a(s_169), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1734(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1735(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1736(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2199(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2200(.a(gate409inter0), .b(s_236), .O(gate409inter1));
  and2  gate2201(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2202(.a(s_236), .O(gate409inter3));
  inv1  gate2203(.a(s_237), .O(gate409inter4));
  nand2 gate2204(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2205(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2206(.a(G23), .O(gate409inter7));
  inv1  gate2207(.a(G1102), .O(gate409inter8));
  nand2 gate2208(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2209(.a(s_237), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2210(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2211(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2212(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1947(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1948(.a(gate410inter0), .b(s_200), .O(gate410inter1));
  and2  gate1949(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1950(.a(s_200), .O(gate410inter3));
  inv1  gate1951(.a(s_201), .O(gate410inter4));
  nand2 gate1952(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1953(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1954(.a(G24), .O(gate410inter7));
  inv1  gate1955(.a(G1105), .O(gate410inter8));
  nand2 gate1956(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1957(.a(s_201), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1958(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1959(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1960(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1205(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1206(.a(gate413inter0), .b(s_94), .O(gate413inter1));
  and2  gate1207(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1208(.a(s_94), .O(gate413inter3));
  inv1  gate1209(.a(s_95), .O(gate413inter4));
  nand2 gate1210(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1211(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1212(.a(G27), .O(gate413inter7));
  inv1  gate1213(.a(G1114), .O(gate413inter8));
  nand2 gate1214(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1215(.a(s_95), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1216(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1217(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1218(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2213(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2214(.a(gate425inter0), .b(s_238), .O(gate425inter1));
  and2  gate2215(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2216(.a(s_238), .O(gate425inter3));
  inv1  gate2217(.a(s_239), .O(gate425inter4));
  nand2 gate2218(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2219(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2220(.a(G4), .O(gate425inter7));
  inv1  gate2221(.a(G1141), .O(gate425inter8));
  nand2 gate2222(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2223(.a(s_239), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2224(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2225(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2226(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1793(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1794(.a(gate427inter0), .b(s_178), .O(gate427inter1));
  and2  gate1795(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1796(.a(s_178), .O(gate427inter3));
  inv1  gate1797(.a(s_179), .O(gate427inter4));
  nand2 gate1798(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1799(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1800(.a(G5), .O(gate427inter7));
  inv1  gate1801(.a(G1144), .O(gate427inter8));
  nand2 gate1802(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1803(.a(s_179), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1804(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1805(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1806(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate995(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate996(.a(gate431inter0), .b(s_64), .O(gate431inter1));
  and2  gate997(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate998(.a(s_64), .O(gate431inter3));
  inv1  gate999(.a(s_65), .O(gate431inter4));
  nand2 gate1000(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1001(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1002(.a(G7), .O(gate431inter7));
  inv1  gate1003(.a(G1150), .O(gate431inter8));
  nand2 gate1004(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1005(.a(s_65), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1006(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1007(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1008(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2241(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2242(.a(gate435inter0), .b(s_242), .O(gate435inter1));
  and2  gate2243(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2244(.a(s_242), .O(gate435inter3));
  inv1  gate2245(.a(s_243), .O(gate435inter4));
  nand2 gate2246(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2247(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2248(.a(G9), .O(gate435inter7));
  inv1  gate2249(.a(G1156), .O(gate435inter8));
  nand2 gate2250(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2251(.a(s_243), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2252(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2253(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2254(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate547(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate548(.a(gate436inter0), .b(s_0), .O(gate436inter1));
  and2  gate549(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate550(.a(s_0), .O(gate436inter3));
  inv1  gate551(.a(s_1), .O(gate436inter4));
  nand2 gate552(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate553(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate554(.a(G1060), .O(gate436inter7));
  inv1  gate555(.a(G1156), .O(gate436inter8));
  nand2 gate556(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate557(.a(s_1), .b(gate436inter3), .O(gate436inter10));
  nor2  gate558(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate559(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate560(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2297(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2298(.a(gate442inter0), .b(s_250), .O(gate442inter1));
  and2  gate2299(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2300(.a(s_250), .O(gate442inter3));
  inv1  gate2301(.a(s_251), .O(gate442inter4));
  nand2 gate2302(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2303(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2304(.a(G1069), .O(gate442inter7));
  inv1  gate2305(.a(G1165), .O(gate442inter8));
  nand2 gate2306(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2307(.a(s_251), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2308(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2309(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2310(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1779(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1780(.a(gate458inter0), .b(s_176), .O(gate458inter1));
  and2  gate1781(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1782(.a(s_176), .O(gate458inter3));
  inv1  gate1783(.a(s_177), .O(gate458inter4));
  nand2 gate1784(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1785(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1786(.a(G1093), .O(gate458inter7));
  inv1  gate1787(.a(G1189), .O(gate458inter8));
  nand2 gate1788(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1789(.a(s_177), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1790(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1791(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1792(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1233(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1234(.a(gate462inter0), .b(s_98), .O(gate462inter1));
  and2  gate1235(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1236(.a(s_98), .O(gate462inter3));
  inv1  gate1237(.a(s_99), .O(gate462inter4));
  nand2 gate1238(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1239(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1240(.a(G1099), .O(gate462inter7));
  inv1  gate1241(.a(G1195), .O(gate462inter8));
  nand2 gate1242(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1243(.a(s_99), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1244(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1245(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1246(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate813(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate814(.a(gate470inter0), .b(s_38), .O(gate470inter1));
  and2  gate815(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate816(.a(s_38), .O(gate470inter3));
  inv1  gate817(.a(s_39), .O(gate470inter4));
  nand2 gate818(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate819(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate820(.a(G1111), .O(gate470inter7));
  inv1  gate821(.a(G1207), .O(gate470inter8));
  nand2 gate822(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate823(.a(s_39), .b(gate470inter3), .O(gate470inter10));
  nor2  gate824(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate825(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate826(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1051(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1052(.a(gate471inter0), .b(s_72), .O(gate471inter1));
  and2  gate1053(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1054(.a(s_72), .O(gate471inter3));
  inv1  gate1055(.a(s_73), .O(gate471inter4));
  nand2 gate1056(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1057(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1058(.a(G27), .O(gate471inter7));
  inv1  gate1059(.a(G1210), .O(gate471inter8));
  nand2 gate1060(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1061(.a(s_73), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1062(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1063(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1064(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2003(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2004(.a(gate475inter0), .b(s_208), .O(gate475inter1));
  and2  gate2005(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2006(.a(s_208), .O(gate475inter3));
  inv1  gate2007(.a(s_209), .O(gate475inter4));
  nand2 gate2008(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2009(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2010(.a(G29), .O(gate475inter7));
  inv1  gate2011(.a(G1216), .O(gate475inter8));
  nand2 gate2012(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2013(.a(s_209), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2014(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2015(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2016(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2185(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2186(.a(gate476inter0), .b(s_234), .O(gate476inter1));
  and2  gate2187(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2188(.a(s_234), .O(gate476inter3));
  inv1  gate2189(.a(s_235), .O(gate476inter4));
  nand2 gate2190(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2191(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2192(.a(G1120), .O(gate476inter7));
  inv1  gate2193(.a(G1216), .O(gate476inter8));
  nand2 gate2194(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2195(.a(s_235), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2196(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2197(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2198(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1695(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1696(.a(gate479inter0), .b(s_164), .O(gate479inter1));
  and2  gate1697(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1698(.a(s_164), .O(gate479inter3));
  inv1  gate1699(.a(s_165), .O(gate479inter4));
  nand2 gate1700(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1701(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1702(.a(G31), .O(gate479inter7));
  inv1  gate1703(.a(G1222), .O(gate479inter8));
  nand2 gate1704(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1705(.a(s_165), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1706(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1707(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1708(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1289(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1290(.a(gate482inter0), .b(s_106), .O(gate482inter1));
  and2  gate1291(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1292(.a(s_106), .O(gate482inter3));
  inv1  gate1293(.a(s_107), .O(gate482inter4));
  nand2 gate1294(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1295(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1296(.a(G1129), .O(gate482inter7));
  inv1  gate1297(.a(G1225), .O(gate482inter8));
  nand2 gate1298(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1299(.a(s_107), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1300(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1301(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1302(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1597(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1598(.a(gate485inter0), .b(s_150), .O(gate485inter1));
  and2  gate1599(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1600(.a(s_150), .O(gate485inter3));
  inv1  gate1601(.a(s_151), .O(gate485inter4));
  nand2 gate1602(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1603(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1604(.a(G1232), .O(gate485inter7));
  inv1  gate1605(.a(G1233), .O(gate485inter8));
  nand2 gate1606(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1607(.a(s_151), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1608(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1609(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1610(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1485(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1486(.a(gate488inter0), .b(s_134), .O(gate488inter1));
  and2  gate1487(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1488(.a(s_134), .O(gate488inter3));
  inv1  gate1489(.a(s_135), .O(gate488inter4));
  nand2 gate1490(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1491(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1492(.a(G1238), .O(gate488inter7));
  inv1  gate1493(.a(G1239), .O(gate488inter8));
  nand2 gate1494(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1495(.a(s_135), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1496(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1497(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1498(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1555(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1556(.a(gate490inter0), .b(s_144), .O(gate490inter1));
  and2  gate1557(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1558(.a(s_144), .O(gate490inter3));
  inv1  gate1559(.a(s_145), .O(gate490inter4));
  nand2 gate1560(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1561(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1562(.a(G1242), .O(gate490inter7));
  inv1  gate1563(.a(G1243), .O(gate490inter8));
  nand2 gate1564(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1565(.a(s_145), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1566(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1567(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1568(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate645(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate646(.a(gate492inter0), .b(s_14), .O(gate492inter1));
  and2  gate647(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate648(.a(s_14), .O(gate492inter3));
  inv1  gate649(.a(s_15), .O(gate492inter4));
  nand2 gate650(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate651(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate652(.a(G1246), .O(gate492inter7));
  inv1  gate653(.a(G1247), .O(gate492inter8));
  nand2 gate654(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate655(.a(s_15), .b(gate492inter3), .O(gate492inter10));
  nor2  gate656(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate657(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate658(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1765(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1766(.a(gate494inter0), .b(s_174), .O(gate494inter1));
  and2  gate1767(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1768(.a(s_174), .O(gate494inter3));
  inv1  gate1769(.a(s_175), .O(gate494inter4));
  nand2 gate1770(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1771(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1772(.a(G1250), .O(gate494inter7));
  inv1  gate1773(.a(G1251), .O(gate494inter8));
  nand2 gate1774(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1775(.a(s_175), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1776(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1777(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1778(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1275(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1276(.a(gate505inter0), .b(s_104), .O(gate505inter1));
  and2  gate1277(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1278(.a(s_104), .O(gate505inter3));
  inv1  gate1279(.a(s_105), .O(gate505inter4));
  nand2 gate1280(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1281(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1282(.a(G1272), .O(gate505inter7));
  inv1  gate1283(.a(G1273), .O(gate505inter8));
  nand2 gate1284(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1285(.a(s_105), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1286(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1287(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1288(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule