module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate637(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate638(.a(gate19inter0), .b(s_68), .O(gate19inter1));
  and2  gate639(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate640(.a(s_68), .O(gate19inter3));
  inv1  gate641(.a(s_69), .O(gate19inter4));
  nand2 gate642(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate643(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate644(.a(N118), .O(gate19inter7));
  inv1  gate645(.a(N4), .O(gate19inter8));
  nand2 gate646(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate647(.a(s_69), .b(gate19inter3), .O(gate19inter10));
  nor2  gate648(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate649(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate650(.a(gate19inter12), .b(gate19inter1), .O(N154));
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate189(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate190(.a(gate22inter0), .b(s_4), .O(gate22inter1));
  and2  gate191(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate192(.a(s_4), .O(gate22inter3));
  inv1  gate193(.a(s_5), .O(gate22inter4));
  nand2 gate194(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate195(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate196(.a(N122), .O(gate22inter7));
  inv1  gate197(.a(N17), .O(gate22inter8));
  nand2 gate198(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate199(.a(s_5), .b(gate22inter3), .O(gate22inter10));
  nor2  gate200(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate201(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate202(.a(gate22inter12), .b(gate22inter1), .O(N159));

  xor2  gate427(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate428(.a(gate23inter0), .b(s_38), .O(gate23inter1));
  and2  gate429(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate430(.a(s_38), .O(gate23inter3));
  inv1  gate431(.a(s_39), .O(gate23inter4));
  nand2 gate432(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate433(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate434(.a(N126), .O(gate23inter7));
  inv1  gate435(.a(N30), .O(gate23inter8));
  nand2 gate436(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate437(.a(s_39), .b(gate23inter3), .O(gate23inter10));
  nor2  gate438(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate439(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate440(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate203(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate204(.a(gate27inter0), .b(s_6), .O(gate27inter1));
  and2  gate205(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate206(.a(s_6), .O(gate27inter3));
  inv1  gate207(.a(s_7), .O(gate27inter4));
  nand2 gate208(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate209(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate210(.a(N142), .O(gate27inter7));
  inv1  gate211(.a(N82), .O(gate27inter8));
  nand2 gate212(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate213(.a(s_7), .b(gate27inter3), .O(gate27inter10));
  nor2  gate214(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate215(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate216(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate329(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate330(.a(gate29inter0), .b(s_24), .O(gate29inter1));
  and2  gate331(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate332(.a(s_24), .O(gate29inter3));
  inv1  gate333(.a(s_25), .O(gate29inter4));
  nand2 gate334(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate335(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate336(.a(N150), .O(gate29inter7));
  inv1  gate337(.a(N108), .O(gate29inter8));
  nand2 gate338(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate339(.a(s_25), .b(gate29inter3), .O(gate29inter10));
  nor2  gate340(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate341(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate342(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );

  xor2  gate175(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate176(.a(gate31inter0), .b(s_2), .O(gate31inter1));
  and2  gate177(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate178(.a(s_2), .O(gate31inter3));
  inv1  gate179(.a(s_3), .O(gate31inter4));
  nand2 gate180(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate181(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate182(.a(N27), .O(gate31inter7));
  inv1  gate183(.a(N123), .O(gate31inter8));
  nand2 gate184(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate185(.a(s_3), .b(gate31inter3), .O(gate31inter10));
  nor2  gate186(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate187(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate188(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );

  xor2  gate273(.a(N127), .b(N40), .O(gate33inter0));
  nand2 gate274(.a(gate33inter0), .b(s_16), .O(gate33inter1));
  and2  gate275(.a(N127), .b(N40), .O(gate33inter2));
  inv1  gate276(.a(s_16), .O(gate33inter3));
  inv1  gate277(.a(s_17), .O(gate33inter4));
  nand2 gate278(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate279(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate280(.a(N40), .O(gate33inter7));
  inv1  gate281(.a(N127), .O(gate33inter8));
  nand2 gate282(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate283(.a(s_17), .b(gate33inter3), .O(gate33inter10));
  nor2  gate284(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate285(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate286(.a(gate33inter12), .b(gate33inter1), .O(N186));

  xor2  gate483(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate484(.a(gate34inter0), .b(s_46), .O(gate34inter1));
  and2  gate485(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate486(.a(s_46), .O(gate34inter3));
  inv1  gate487(.a(s_47), .O(gate34inter4));
  nand2 gate488(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate489(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate490(.a(N47), .O(gate34inter7));
  inv1  gate491(.a(N131), .O(gate34inter8));
  nand2 gate492(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate493(.a(s_47), .b(gate34inter3), .O(gate34inter10));
  nor2  gate494(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate495(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate496(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate357(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate358(.a(gate35inter0), .b(s_28), .O(gate35inter1));
  and2  gate359(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate360(.a(s_28), .O(gate35inter3));
  inv1  gate361(.a(s_29), .O(gate35inter4));
  nand2 gate362(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate363(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate364(.a(N53), .O(gate35inter7));
  inv1  gate365(.a(N131), .O(gate35inter8));
  nand2 gate366(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate367(.a(s_29), .b(gate35inter3), .O(gate35inter10));
  nor2  gate368(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate369(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate370(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate651(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate652(.a(gate43inter0), .b(s_70), .O(gate43inter1));
  and2  gate653(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate654(.a(s_70), .O(gate43inter3));
  inv1  gate655(.a(s_71), .O(gate43inter4));
  nand2 gate656(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate657(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate658(.a(N105), .O(gate43inter7));
  inv1  gate659(.a(N147), .O(gate43inter8));
  nand2 gate660(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate661(.a(s_71), .b(gate43inter3), .O(gate43inter10));
  nor2  gate662(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate663(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate664(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );

  xor2  gate399(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate400(.a(gate45inter0), .b(s_34), .O(gate45inter1));
  and2  gate401(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate402(.a(s_34), .O(gate45inter3));
  inv1  gate403(.a(s_35), .O(gate45inter4));
  nand2 gate404(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate405(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate406(.a(N115), .O(gate45inter7));
  inv1  gate407(.a(N151), .O(gate45inter8));
  nand2 gate408(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate409(.a(s_35), .b(gate45inter3), .O(gate45inter10));
  nor2  gate410(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate411(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate412(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate497(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate498(.a(gate50inter0), .b(s_48), .O(gate50inter1));
  and2  gate499(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate500(.a(s_48), .O(gate50inter3));
  inv1  gate501(.a(s_49), .O(gate50inter4));
  nand2 gate502(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate503(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate504(.a(N203), .O(gate50inter7));
  inv1  gate505(.a(N154), .O(gate50inter8));
  nand2 gate506(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate507(.a(s_49), .b(gate50inter3), .O(gate50inter10));
  nor2  gate508(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate509(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate510(.a(gate50inter12), .b(gate50inter1), .O(N224));
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );

  xor2  gate525(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate526(.a(gate53inter0), .b(s_52), .O(gate53inter1));
  and2  gate527(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate528(.a(s_52), .O(gate53inter3));
  inv1  gate529(.a(s_53), .O(gate53inter4));
  nand2 gate530(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate531(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate532(.a(N203), .O(gate53inter7));
  inv1  gate533(.a(N165), .O(gate53inter8));
  nand2 gate534(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate535(.a(s_53), .b(gate53inter3), .O(gate53inter10));
  nor2  gate536(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate537(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate538(.a(gate53inter12), .b(gate53inter1), .O(N233));

  xor2  gate623(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate624(.a(gate54inter0), .b(s_66), .O(gate54inter1));
  and2  gate625(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate626(.a(s_66), .O(gate54inter3));
  inv1  gate627(.a(s_67), .O(gate54inter4));
  nand2 gate628(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate629(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate630(.a(N203), .O(gate54inter7));
  inv1  gate631(.a(N168), .O(gate54inter8));
  nand2 gate632(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate633(.a(s_67), .b(gate54inter3), .O(gate54inter10));
  nor2  gate634(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate635(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate636(.a(gate54inter12), .b(gate54inter1), .O(N236));

  xor2  gate693(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate694(.a(gate55inter0), .b(s_76), .O(gate55inter1));
  and2  gate695(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate696(.a(s_76), .O(gate55inter3));
  inv1  gate697(.a(s_77), .O(gate55inter4));
  nand2 gate698(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate699(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate700(.a(N203), .O(gate55inter7));
  inv1  gate701(.a(N171), .O(gate55inter8));
  nand2 gate702(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate703(.a(s_77), .b(gate55inter3), .O(gate55inter10));
  nor2  gate704(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate705(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate706(.a(gate55inter12), .b(gate55inter1), .O(N239));
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate581(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate582(.a(gate57inter0), .b(s_60), .O(gate57inter1));
  and2  gate583(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate584(.a(s_60), .O(gate57inter3));
  inv1  gate585(.a(s_61), .O(gate57inter4));
  nand2 gate586(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate587(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate588(.a(N203), .O(gate57inter7));
  inv1  gate589(.a(N174), .O(gate57inter8));
  nand2 gate590(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate591(.a(s_61), .b(gate57inter3), .O(gate57inter10));
  nor2  gate592(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate593(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate594(.a(gate57inter12), .b(gate57inter1), .O(N243));

  xor2  gate287(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate288(.a(gate58inter0), .b(s_18), .O(gate58inter1));
  and2  gate289(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate290(.a(s_18), .O(gate58inter3));
  inv1  gate291(.a(s_19), .O(gate58inter4));
  nand2 gate292(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate293(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate294(.a(N213), .O(gate58inter7));
  inv1  gate295(.a(N11), .O(gate58inter8));
  nand2 gate296(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate297(.a(s_19), .b(gate58inter3), .O(gate58inter10));
  nor2  gate298(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate299(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate300(.a(gate58inter12), .b(gate58inter1), .O(N246));
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate511(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate512(.a(gate60inter0), .b(s_50), .O(gate60inter1));
  and2  gate513(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate514(.a(s_50), .O(gate60inter3));
  inv1  gate515(.a(s_51), .O(gate60inter4));
  nand2 gate516(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate517(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate518(.a(N213), .O(gate60inter7));
  inv1  gate519(.a(N24), .O(gate60inter8));
  nand2 gate520(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate521(.a(s_51), .b(gate60inter3), .O(gate60inter10));
  nor2  gate522(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate523(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate524(.a(gate60inter12), .b(gate60inter1), .O(N250));
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );

  xor2  gate567(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate568(.a(gate64inter0), .b(s_58), .O(gate64inter1));
  and2  gate569(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate570(.a(s_58), .O(gate64inter3));
  inv1  gate571(.a(s_59), .O(gate64inter4));
  nand2 gate572(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate573(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate574(.a(N213), .O(gate64inter7));
  inv1  gate575(.a(N63), .O(gate64inter8));
  nand2 gate576(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate577(.a(s_59), .b(gate64inter3), .O(gate64inter10));
  nor2  gate578(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate579(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate580(.a(gate64inter12), .b(gate64inter1), .O(N256));
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );

  xor2  gate259(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate260(.a(gate69inter0), .b(s_14), .O(gate69inter1));
  and2  gate261(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate262(.a(s_14), .O(gate69inter3));
  inv1  gate263(.a(s_15), .O(gate69inter4));
  nand2 gate264(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate265(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate266(.a(N224), .O(gate69inter7));
  inv1  gate267(.a(N158), .O(gate69inter8));
  nand2 gate268(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate269(.a(s_15), .b(gate69inter3), .O(gate69inter10));
  nor2  gate270(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate271(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate272(.a(gate69inter12), .b(gate69inter1), .O(N263));

  xor2  gate161(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate162(.a(gate70inter0), .b(s_0), .O(gate70inter1));
  and2  gate163(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate164(.a(s_0), .O(gate70inter3));
  inv1  gate165(.a(s_1), .O(gate70inter4));
  nand2 gate166(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate167(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate168(.a(N227), .O(gate70inter7));
  inv1  gate169(.a(N183), .O(gate70inter8));
  nand2 gate170(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate171(.a(s_1), .b(gate70inter3), .O(gate70inter10));
  nor2  gate172(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate173(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate174(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate343(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate344(.a(gate72inter0), .b(s_26), .O(gate72inter1));
  and2  gate345(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate346(.a(s_26), .O(gate72inter3));
  inv1  gate347(.a(s_27), .O(gate72inter4));
  nand2 gate348(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate349(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate350(.a(N233), .O(gate72inter7));
  inv1  gate351(.a(N187), .O(gate72inter8));
  nand2 gate352(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate353(.a(s_27), .b(gate72inter3), .O(gate72inter10));
  nor2  gate354(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate355(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate356(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate665(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate666(.a(gate77inter0), .b(s_72), .O(gate77inter1));
  and2  gate667(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate668(.a(s_72), .O(gate77inter3));
  inv1  gate669(.a(s_73), .O(gate77inter4));
  nand2 gate670(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate671(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate672(.a(N251), .O(gate77inter7));
  inv1  gate673(.a(N197), .O(gate77inter8));
  nand2 gate674(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate675(.a(s_73), .b(gate77inter3), .O(gate77inter10));
  nor2  gate676(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate677(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate678(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );

  xor2  gate553(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate554(.a(gate81inter0), .b(s_56), .O(gate81inter1));
  and2  gate555(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate556(.a(s_56), .O(gate81inter3));
  inv1  gate557(.a(s_57), .O(gate81inter4));
  nand2 gate558(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate559(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate560(.a(N236), .O(gate81inter7));
  inv1  gate561(.a(N190), .O(gate81inter8));
  nand2 gate562(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate563(.a(s_57), .b(gate81inter3), .O(gate81inter10));
  nor2  gate564(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate565(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate566(.a(gate81inter12), .b(gate81inter1), .O(N291));
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate371(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate372(.a(gate83inter0), .b(s_30), .O(gate83inter1));
  and2  gate373(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate374(.a(s_30), .O(gate83inter3));
  inv1  gate375(.a(s_31), .O(gate83inter4));
  nand2 gate376(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate377(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate378(.a(N243), .O(gate83inter7));
  inv1  gate379(.a(N194), .O(gate83inter8));
  nand2 gate380(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate381(.a(s_31), .b(gate83inter3), .O(gate83inter10));
  nor2  gate382(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate383(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate384(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );

  xor2  gate245(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate246(.a(gate85inter0), .b(s_12), .O(gate85inter1));
  and2  gate247(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate248(.a(s_12), .O(gate85inter3));
  inv1  gate249(.a(s_13), .O(gate85inter4));
  nand2 gate250(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate251(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate252(.a(N251), .O(gate85inter7));
  inv1  gate253(.a(N198), .O(gate85inter8));
  nand2 gate254(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate255(.a(s_13), .b(gate85inter3), .O(gate85inter10));
  nor2  gate256(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate257(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate258(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );

  xor2  gate231(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate232(.a(gate100inter0), .b(s_10), .O(gate100inter1));
  and2  gate233(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate234(.a(s_10), .O(gate100inter3));
  inv1  gate235(.a(s_11), .O(gate100inter4));
  nand2 gate236(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate237(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate238(.a(N309), .O(gate100inter7));
  inv1  gate239(.a(N264), .O(gate100inter8));
  nand2 gate240(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate241(.a(s_11), .b(gate100inter3), .O(gate100inter10));
  nor2  gate242(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate243(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate244(.a(gate100inter12), .b(gate100inter1), .O(N331));
xor2 gate101( .a(N309), .b(N267), .O(N332) );

  xor2  gate315(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate316(.a(gate102inter0), .b(s_22), .O(gate102inter1));
  and2  gate317(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate318(.a(s_22), .O(gate102inter3));
  inv1  gate319(.a(s_23), .O(gate102inter4));
  nand2 gate320(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate321(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate322(.a(N309), .O(gate102inter7));
  inv1  gate323(.a(N270), .O(gate102inter8));
  nand2 gate324(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate325(.a(s_23), .b(gate102inter3), .O(gate102inter10));
  nor2  gate326(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate327(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate328(.a(gate102inter12), .b(gate102inter1), .O(N333));
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );

  xor2  gate441(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate442(.a(gate106inter0), .b(s_40), .O(gate106inter1));
  and2  gate443(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate444(.a(s_40), .O(gate106inter3));
  inv1  gate445(.a(s_41), .O(gate106inter4));
  nand2 gate446(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate447(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate448(.a(N309), .O(gate106inter7));
  inv1  gate449(.a(N276), .O(gate106inter8));
  nand2 gate450(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate451(.a(s_41), .b(gate106inter3), .O(gate106inter10));
  nor2  gate452(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate453(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate454(.a(gate106inter12), .b(gate106inter1), .O(N337));
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate707(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate708(.a(gate110inter0), .b(s_78), .O(gate110inter1));
  and2  gate709(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate710(.a(s_78), .O(gate110inter3));
  inv1  gate711(.a(s_79), .O(gate110inter4));
  nand2 gate712(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate713(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate714(.a(N309), .O(gate110inter7));
  inv1  gate715(.a(N282), .O(gate110inter8));
  nand2 gate716(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate717(.a(s_79), .b(gate110inter3), .O(gate110inter10));
  nor2  gate718(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate719(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate720(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );

  xor2  gate609(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate610(.a(gate112inter0), .b(s_64), .O(gate112inter1));
  and2  gate611(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate612(.a(s_64), .O(gate112inter3));
  inv1  gate613(.a(s_65), .O(gate112inter4));
  nand2 gate614(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate615(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate616(.a(N309), .O(gate112inter7));
  inv1  gate617(.a(N285), .O(gate112inter8));
  nand2 gate618(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate619(.a(s_65), .b(gate112inter3), .O(gate112inter10));
  nor2  gate620(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate621(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate622(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate679(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate680(.a(gate120inter0), .b(s_74), .O(gate120inter1));
  and2  gate681(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate682(.a(s_74), .O(gate120inter3));
  inv1  gate683(.a(s_75), .O(gate120inter4));
  nand2 gate684(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate685(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate686(.a(N333), .O(gate120inter7));
  inv1  gate687(.a(N303), .O(gate120inter8));
  nand2 gate688(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate689(.a(s_75), .b(gate120inter3), .O(gate120inter10));
  nor2  gate690(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate691(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate692(.a(gate120inter12), .b(gate120inter1), .O(N351));

  xor2  gate385(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate386(.a(gate121inter0), .b(s_32), .O(gate121inter1));
  and2  gate387(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate388(.a(s_32), .O(gate121inter3));
  inv1  gate389(.a(s_33), .O(gate121inter4));
  nand2 gate390(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate391(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate392(.a(N335), .O(gate121inter7));
  inv1  gate393(.a(N304), .O(gate121inter8));
  nand2 gate394(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate395(.a(s_33), .b(gate121inter3), .O(gate121inter10));
  nor2  gate396(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate397(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate398(.a(gate121inter12), .b(gate121inter1), .O(N352));
nand2 gate122( .a(N337), .b(N305), .O(N353) );

  xor2  gate595(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate596(.a(gate123inter0), .b(s_62), .O(gate123inter1));
  and2  gate597(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate598(.a(s_62), .O(gate123inter3));
  inv1  gate599(.a(s_63), .O(gate123inter4));
  nand2 gate600(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate601(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate602(.a(N339), .O(gate123inter7));
  inv1  gate603(.a(N306), .O(gate123inter8));
  nand2 gate604(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate605(.a(s_63), .b(gate123inter3), .O(gate123inter10));
  nor2  gate606(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate607(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate608(.a(gate123inter12), .b(gate123inter1), .O(N354));

  xor2  gate721(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate722(.a(gate124inter0), .b(s_80), .O(gate124inter1));
  and2  gate723(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate724(.a(s_80), .O(gate124inter3));
  inv1  gate725(.a(s_81), .O(gate124inter4));
  nand2 gate726(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate727(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate728(.a(N341), .O(gate124inter7));
  inv1  gate729(.a(N307), .O(gate124inter8));
  nand2 gate730(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate731(.a(s_81), .b(gate124inter3), .O(gate124inter10));
  nor2  gate732(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate733(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate734(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate301(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate302(.a(gate131inter0), .b(s_20), .O(gate131inter1));
  and2  gate303(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate304(.a(s_20), .O(gate131inter3));
  inv1  gate305(.a(s_21), .O(gate131inter4));
  nand2 gate306(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate307(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate308(.a(N360), .O(gate131inter7));
  inv1  gate309(.a(N40), .O(gate131inter8));
  nand2 gate310(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate311(.a(s_21), .b(gate131inter3), .O(gate131inter10));
  nor2  gate312(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate313(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate314(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );

  xor2  gate455(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate456(.a(gate133inter0), .b(s_42), .O(gate133inter1));
  and2  gate457(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate458(.a(s_42), .O(gate133inter3));
  inv1  gate459(.a(s_43), .O(gate133inter4));
  nand2 gate460(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate461(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate462(.a(N360), .O(gate133inter7));
  inv1  gate463(.a(N66), .O(gate133inter8));
  nand2 gate464(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate465(.a(s_43), .b(gate133inter3), .O(gate133inter10));
  nor2  gate466(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate467(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate468(.a(gate133inter12), .b(gate133inter1), .O(N375));
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate539(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate540(.a(gate135inter0), .b(s_54), .O(gate135inter1));
  and2  gate541(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate542(.a(s_54), .O(gate135inter3));
  inv1  gate543(.a(s_55), .O(gate135inter4));
  nand2 gate544(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate545(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate546(.a(N360), .O(gate135inter7));
  inv1  gate547(.a(N92), .O(gate135inter8));
  nand2 gate548(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate549(.a(s_55), .b(gate135inter3), .O(gate135inter10));
  nor2  gate550(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate551(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate552(.a(gate135inter12), .b(gate135inter1), .O(N377));

  xor2  gate217(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate218(.a(gate136inter0), .b(s_8), .O(gate136inter1));
  and2  gate219(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate220(.a(s_8), .O(gate136inter3));
  inv1  gate221(.a(s_9), .O(gate136inter4));
  nand2 gate222(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate223(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate224(.a(N360), .O(gate136inter7));
  inv1  gate225(.a(N105), .O(gate136inter8));
  nand2 gate226(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate227(.a(s_9), .b(gate136inter3), .O(gate136inter10));
  nor2  gate228(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate229(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate230(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate469(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate470(.a(gate153inter0), .b(s_44), .O(gate153inter1));
  and2  gate471(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate472(.a(s_44), .O(gate153inter3));
  inv1  gate473(.a(s_45), .O(gate153inter4));
  nand2 gate474(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate475(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate476(.a(N415), .O(gate153inter7));
  inv1  gate477(.a(N416), .O(gate153inter8));
  nand2 gate478(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate479(.a(s_45), .b(gate153inter3), .O(gate153inter10));
  nor2  gate480(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate481(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate482(.a(gate153inter12), .b(gate153inter1), .O(N421));

  xor2  gate413(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate414(.a(gate154inter0), .b(s_36), .O(gate154inter1));
  and2  gate415(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate416(.a(s_36), .O(gate154inter3));
  inv1  gate417(.a(s_37), .O(gate154inter4));
  nand2 gate418(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate419(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate420(.a(N386), .O(gate154inter7));
  inv1  gate421(.a(N417), .O(gate154inter8));
  nand2 gate422(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate423(.a(s_37), .b(gate154inter3), .O(gate154inter10));
  nor2  gate424(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate425(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate426(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule