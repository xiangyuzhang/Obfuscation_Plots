
module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input  N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,      N99,N102,N105,N108,N112,N115,CONST1,CONST0 //RE__PI;

input D_0,D_1,D_2,D_3,D_4,D_5,D_6,D_7,D_8,D_9,D_10,D_11,D_12,D_13,D_14,D_15,D_16,D_17,D_18,D_19,D_20,D_21,D_22,D_23,D_24,D_25,D_26,D_27,D_28,D_29,D_30,D_31,D_32,D_33,D_34,D_35,D_36,D_37,D_38,D_39,D_40,D_41,D_42,D_43,D_44,D_45,D_46,D_47,D_48,D_49,D_50,D_51,D_52,D_53,D_54,D_55,D_56,D_57,D_58,D_59,D_60,D_61,D_62,D_63,D_64,D_65,D_66,D_67,D_68,D_69,D_70,D_71,D_72,D_73,D_74,D_75,D_76,D_77,D_78,D_79,D_80,D_81,D_82,D_83,D_84,D_85,D_86,D_87,D_88,D_89,D_90,D_91,D_92,D_93,D_94,D_95,D_96,D_97,D_98,D_99,D_100,D_101,D_102,D_103,D_104,D_105,D_106,D_107,D_108,D_109,D_110,D_111 //RE__ALLOW(00,01,10,11);

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429,D_0_NOT,D_1_NOT,N289_NOT,N289_OBF,ED_0,ED_1,ED_2,ED_3,ED_4,ED_5,ED_6,ED_7,ED_8,ED_9,D_2_NOT,D_3_NOT,N213_NOT,N213_OBF,ED_10,ED_11,ED_12,ED_13,ED_14,ED_15,ED_16,ED_17,ED_18,ED_19,D_4_NOT,D_5_NOT,N69_NOT,N69_OBF,ED_20,ED_21,ED_22,ED_23,ED_24,ED_25,ED_26,ED_27,ED_28,ED_29,D_6_NOT,D_7_NOT,N227_NOT,N227_OBF,ED_30,ED_31,ED_32,ED_33,ED_34,ED_35,ED_36,ED_37,ED_38,ED_39,D_8_NOT,D_9_NOT,N416_NOT,N416_OBF,ED_40,ED_41,ED_42,ED_43,ED_44,ED_45,ED_46,ED_47,ED_48,ED_49,D_10_NOT,D_11_NOT,N213_NOT,N213_OBF,ED_50,ED_51,ED_52,ED_53,ED_54,ED_55,ED_56,ED_57,ED_58,ED_59,D_12_NOT,D_13_NOT,N30_NOT,N30_OBF,ED_60,ED_61,ED_62,ED_63,ED_64,ED_65,ED_66,ED_67,ED_68,ED_69,D_14_NOT,D_15_NOT,N360_NOT,N360_OBF,ED_70,ED_71,ED_72,ED_73,ED_74,ED_75,ED_76,ED_77,ED_78,ED_79,D_16_NOT,D_17_NOT,N99_NOT,N99_OBF,ED_80,ED_81,ED_82,ED_83,ED_84,ED_85,ED_86,ED_87,ED_88,ED_89,D_18_NOT,D_19_NOT,N296_NOT,N296_OBF,ED_90,ED_91,ED_92,ED_93,ED_94,ED_95,ED_96,ED_97,ED_98,ED_99,D_20_NOT,D_21_NOT,N95_NOT,N95_OBF,ED_100,ED_101,ED_102,ED_103,ED_104,ED_105,ED_106,ED_107,ED_108,ED_109,D_22_NOT,D_23_NOT,N357_NOT,N357_OBF,ED_110,ED_111,ED_112,ED_113,ED_114,ED_115,ED_116,ED_117,ED_118,ED_119,D_24_NOT,D_25_NOT,N50_NOT,N50_OBF,ED_120,ED_121,ED_122,ED_123,ED_124,ED_125,ED_126,ED_127,ED_128,ED_129,D_26_NOT,D_27_NOT,N341_NOT,N341_OBF,ED_130,ED_131,ED_132,ED_133,ED_134,ED_135,ED_136,ED_137,ED_138,ED_139,D_28_NOT,D_29_NOT,N267_NOT,N267_OBF,ED_140,ED_141,ED_142,ED_143,ED_144,ED_145,ED_146,ED_147,ED_148,ED_149,D_30_NOT,D_31_NOT,N254_NOT,N254_OBF,ED_150,ED_151,ED_152,ED_153,ED_154,ED_155,ED_156,ED_157,ED_158,ED_159,D_32_NOT,D_33_NOT,N360_NOT,N360_OBF,ED_160,ED_161,ED_162,ED_163,ED_164,ED_165,ED_166,ED_167,ED_168,ED_169,D_34_NOT,D_35_NOT,N196_NOT,N196_OBF,ED_170,ED_171,ED_172,ED_173,ED_174,ED_175,ED_176,ED_177,ED_178,ED_179,D_36_NOT,D_37_NOT,N197_NOT,N197_OBF,ED_180,ED_181,ED_182,ED_183,ED_184,ED_185,ED_186,ED_187,ED_188,ED_189,D_38_NOT,D_39_NOT,N157_NOT,N157_OBF,ED_190,ED_191,ED_192,ED_193,ED_194,ED_195,ED_196,ED_197,ED_198,ED_199,D_40_NOT,D_41_NOT,N50_NOT,N50_OBF,ED_200,ED_201,ED_202,ED_203,ED_204,ED_205,ED_206,ED_207,ED_208,ED_209,D_42_NOT,D_43_NOT,N123_NOT,N123_OBF,ED_210,ED_211,ED_212,ED_213,ED_214,ED_215,ED_216,ED_217,ED_218,ED_219,D_44_NOT,D_45_NOT,N105_NOT,N105_OBF,ED_220,ED_221,ED_222,ED_223,ED_224,ED_225,ED_226,ED_227,ED_228,ED_229,D_46_NOT,D_47_NOT,N102_NOT,N102_OBF,ED_230,ED_231,ED_232,ED_233,ED_234,ED_235,ED_236,ED_237,ED_238,ED_239,D_48_NOT,D_49_NOT,N95_NOT,N95_OBF,ED_240,ED_241,ED_242,ED_243,ED_244,ED_245,ED_246,ED_247,ED_248,ED_249,D_50_NOT,D_51_NOT,N139_NOT,N139_OBF,ED_250,ED_251,ED_252,ED_253,ED_254,ED_255,ED_256,ED_257,ED_258,ED_259,D_52_NOT,D_53_NOT,N295_NOT,N295_OBF,ED_260,ED_261,ED_262,ED_263,ED_264,ED_265,ED_266,ED_267,ED_268,ED_269,D_54_NOT,D_55_NOT,N131_NOT,N131_OBF,ED_270,ED_271,ED_272,ED_273,ED_274,ED_275,ED_276,ED_277,ED_278,ED_279,D_56_NOT,D_57_NOT,N360_NOT,N360_OBF,ED_280,ED_281,ED_282,ED_283,ED_284,ED_285,ED_286,ED_287,ED_288,ED_289,D_58_NOT,D_59_NOT,N334_NOT,N334_OBF,ED_290,ED_291,ED_292,ED_293,ED_294,ED_295,ED_296,ED_297,ED_298,ED_299,D_60_NOT,D_61_NOT,N292_NOT,N292_OBF,ED_300,ED_301,ED_302,ED_303,ED_304,ED_305,ED_306,ED_307,ED_308,ED_309,D_62_NOT,D_63_NOT,N199_NOT,N199_OBF,ED_310,ED_311,ED_312,ED_313,ED_314,ED_315,ED_316,ED_317,ED_318,ED_319,D_64_NOT,D_65_NOT,N112_NOT,N112_OBF,ED_320,ED_321,ED_322,ED_323,ED_324,ED_325,ED_326,ED_327,ED_328,ED_329,D_66_NOT,D_67_NOT,N243_NOT,N243_OBF,ED_330,ED_331,ED_332,ED_333,ED_334,ED_335,ED_336,ED_337,ED_338,ED_339,D_68_NOT,D_69_NOT,N131_NOT,N131_OBF,ED_340,ED_341,ED_342,ED_343,ED_344,ED_345,ED_346,ED_347,ED_348,ED_349,D_70_NOT,D_71_NOT,N191_NOT,N191_OBF,ED_350,ED_351,ED_352,ED_353,ED_354,ED_355,ED_356,ED_357,ED_358,ED_359,D_72_NOT,D_73_NOT,N345_NOT,N345_OBF,ED_360,ED_361,ED_362,ED_363,ED_364,ED_365,ED_366,ED_367,ED_368,ED_369,D_74_NOT,D_75_NOT,N213_NOT,N213_OBF,ED_370,ED_371,ED_372,ED_373,ED_374,ED_375,ED_376,ED_377,ED_378,ED_379,D_76_NOT,D_77_NOT,N1_NOT,N1_OBF,ED_380,ED_381,ED_382,ED_383,ED_384,ED_385,ED_386,ED_387,ED_388,ED_389,D_78_NOT,D_79_NOT,N420_NOT,N420_OBF,ED_390,ED_391,ED_392,ED_393,ED_394,ED_395,ED_396,ED_397,ED_398,ED_399,D_80_NOT,D_81_NOT,N319_NOT,N319_OBF,ED_400,ED_401,ED_402,ED_403,ED_404,ED_405,ED_406,ED_407,ED_408,ED_409,D_82_NOT,D_83_NOT,N294_NOT,N294_OBF,ED_410,ED_411,ED_412,ED_413,ED_414,ED_415,ED_416,ED_417,ED_418,ED_419,D_84_NOT,D_85_NOT,N422_NOT,N422_OBF,ED_420,ED_421,ED_422,ED_423,ED_424,ED_425,ED_426,ED_427,ED_428,ED_429,D_86_NOT,D_87_NOT,N4_NOT,N4_OBF,ED_430,ED_431,ED_432,ED_433,ED_434,ED_435,ED_436,ED_437,ED_438,ED_439,D_88_NOT,D_89_NOT,N56_NOT,N56_OBF,ED_440,ED_441,ED_442,ED_443,ED_444,ED_445,ED_446,ED_447,ED_448,ED_449,D_90_NOT,D_91_NOT,N37_NOT,N37_OBF,ED_450,ED_451,ED_452,ED_453,ED_454,ED_455,ED_456,ED_457,ED_458,ED_459,D_92_NOT,D_93_NOT,N8_NOT,N8_OBF,ED_460,ED_461,ED_462,ED_463,ED_464,ED_465,ED_466,ED_467,ED_468,ED_469,D_94_NOT,D_95_NOT,N34_NOT,N34_OBF,ED_470,ED_471,ED_472,ED_473,ED_474,ED_475,ED_476,ED_477,ED_478,ED_479,D_96_NOT,D_97_NOT,N14_NOT,N14_OBF,ED_480,ED_481,ED_482,ED_483,ED_484,ED_485,ED_486,ED_487,ED_488,ED_489,D_98_NOT,D_99_NOT,N357_NOT,N357_OBF,ED_490,ED_491,ED_492,ED_493,ED_494,ED_495,ED_496,ED_497,ED_498,ED_499,D_100_NOT,D_101_NOT,N411_NOT,N411_OBF,ED_500,ED_501,ED_502,ED_503,ED_504,ED_505,ED_506,ED_507,ED_508,ED_509,D_102_NOT,D_103_NOT,N290_NOT,N290_OBF,ED_510,ED_511,ED_512,ED_513,ED_514,ED_515,ED_516,ED_517,ED_518,ED_519,D_104_NOT,D_105_NOT,N332_NOT,N332_OBF,ED_520,ED_521,ED_522,ED_523,ED_524,ED_525,ED_526,ED_527,ED_528,ED_529,D_106_NOT,D_107_NOT,N230_NOT,N230_OBF,ED_530,ED_531,ED_532,ED_533,ED_534,ED_535,ED_536,ED_537,ED_538,ED_539,D_108_NOT,D_109_NOT,N230_NOT,N230_OBF,ED_540,ED_541,ED_542,ED_543,ED_544,ED_545,ED_546,ED_547,ED_548,ED_549,D_110_NOT,D_111_NOT,N63_NOT,N63_OBF,ED_550,ED_551,ED_552,ED_553,ED_554,ED_555,ED_556,ED_557,ED_558,ED_559;


inv1 gate1( .a(N1_OBF), .O(N118) );
inv1 gate2( .a(N4_OBF), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30_OBF), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50_OBF), .O(N134) );
inv1 gate10( .a(N56_OBF), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69_OBF), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95_OBF), .O(N147) );
inv1 gate17( .a(N102_OBF), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95_OBF), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123_OBF), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131_OBF), .O(N187) );
nor2 gate35( .a(N53), .b(N131_OBF), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139_OBF), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199_OBF), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213_OBF), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213_OBF), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37_OBF), .O(N254) );
nand2 gate63( .a(N213), .b(N50_OBF), .O(N255) );
nand2 gate64( .a(N213), .b(N63_OBF), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213_OBF), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157_OBF), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227_OBF), .b(N183), .O(N264) );
nand2 gate71( .a(N230_OBF), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191_OBF), .O(N276) );
nand2 gate75( .a(N243_OBF), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197_OBF), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230_OBF), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196_OBF), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267_OBF), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289_OBF), .O(N302) );
inv1 gate90( .a(N290_OBF), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292_OBF), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294_OBF), .O(N307) );
inv1 gate95( .a(N295_OBF), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296_OBF), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8_OBF), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34_OBF), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319_OBF), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99_OBF), .O(N346) );
nand2 gate116( .a(N319), .b(N112_OBF), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332_OBF), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341_OBF), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357_OBF), .O(N360) );
inv1 gate128( .a(N357_OBF), .O(N370) );
nand2 gate129( .a(N14_OBF), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360_OBF), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360_OBF), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105_OBF), .O(N378) );
nand2 gate137( .a(N360_OBF), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334_OBF), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254_OBF), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345_OBF), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411_OBF), .O(N420) );
nor2 gate153( .a(N415), .b(N416_OBF), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420_OBF), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422_OBF), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );
inv1 gate( .a(D_0), .O(D_0_NOT) );
inv1 gate( .a(D_1), .O(D_1_NOT) );
inv1 gate( .a(N289), .O(N289_NOT) );
and2 gate( .a(N289), .b(D_0_NOT), .O(ED_0) );
and2 gate( .a(N289_NOT), .b(D_0_NOT), .O(ED_1) );
and2 gate( .a(CONST1), .b(D_0), .O(ED_2) );
and2 gate( .a(CONST0), .b(D_0), .O(ED_3) );
and2 gate( .a(ED_0), .b(D_1_NOT), .O(ED_9) );
and2 gate( .a(ED_1), .b(D_1), .O(ED_7) );
and2 gate( .a(ED_2), .b(D_1_NOT), .O(ED_5) );
and2 gate( .a(ED_3), .b(D_1), .O(ED_4) );
or2  gate( .a(ED_4), .b(ED_5), .O(ED_6) );
or2  gate( .a(ED_6), .b(ED_7), .O(ED_8) );
or2  gate( .a(ED_9), .b(ED_8), .O(N289_OBF) );
inv1 gate( .a(D_2), .O(D_2_NOT) );
inv1 gate( .a(D_3), .O(D_3_NOT) );
inv1 gate( .a(N213), .O(N213_NOT) );
and2 gate( .a(N213), .b(D_2_NOT), .O(ED_10) );
and2 gate( .a(N213_NOT), .b(D_2_NOT), .O(ED_11) );
and2 gate( .a(CONST1), .b(D_2), .O(ED_12) );
and2 gate( .a(CONST0), .b(D_2), .O(ED_13) );
and2 gate( .a(ED_10), .b(D_3_NOT), .O(ED_19) );
and2 gate( .a(ED_11), .b(D_3), .O(ED_17) );
and2 gate( .a(ED_12), .b(D_3_NOT), .O(ED_15) );
and2 gate( .a(ED_13), .b(D_3), .O(ED_14) );
or2  gate( .a(ED_14), .b(ED_15), .O(ED_16) );
or2  gate( .a(ED_16), .b(ED_17), .O(ED_18) );
or2  gate( .a(ED_19), .b(ED_18), .O(N213_OBF) );
inv1 gate( .a(D_4), .O(D_4_NOT) );
inv1 gate( .a(D_5), .O(D_5_NOT) );
inv1 gate( .a(N69), .O(N69_NOT) );
and2 gate( .a(N69), .b(D_4_NOT), .O(ED_20) );
and2 gate( .a(N69_NOT), .b(D_4_NOT), .O(ED_21) );
and2 gate( .a(CONST1), .b(D_4), .O(ED_22) );
and2 gate( .a(CONST0), .b(D_4), .O(ED_23) );
and2 gate( .a(ED_20), .b(D_5_NOT), .O(ED_29) );
and2 gate( .a(ED_21), .b(D_5), .O(ED_27) );
and2 gate( .a(ED_22), .b(D_5_NOT), .O(ED_25) );
and2 gate( .a(ED_23), .b(D_5), .O(ED_24) );
or2  gate( .a(ED_24), .b(ED_25), .O(ED_26) );
or2  gate( .a(ED_26), .b(ED_27), .O(ED_28) );
or2  gate( .a(ED_29), .b(ED_28), .O(N69_OBF) );
inv1 gate( .a(D_6), .O(D_6_NOT) );
inv1 gate( .a(D_7), .O(D_7_NOT) );
inv1 gate( .a(N227), .O(N227_NOT) );
and2 gate( .a(N227), .b(D_6_NOT), .O(ED_30) );
and2 gate( .a(N227_NOT), .b(D_6_NOT), .O(ED_31) );
and2 gate( .a(CONST1), .b(D_6), .O(ED_32) );
and2 gate( .a(CONST0), .b(D_6), .O(ED_33) );
and2 gate( .a(ED_30), .b(D_7_NOT), .O(ED_39) );
and2 gate( .a(ED_31), .b(D_7), .O(ED_37) );
and2 gate( .a(ED_32), .b(D_7_NOT), .O(ED_35) );
and2 gate( .a(ED_33), .b(D_7), .O(ED_34) );
or2  gate( .a(ED_34), .b(ED_35), .O(ED_36) );
or2  gate( .a(ED_36), .b(ED_37), .O(ED_38) );
or2  gate( .a(ED_39), .b(ED_38), .O(N227_OBF) );
inv1 gate( .a(D_8), .O(D_8_NOT) );
inv1 gate( .a(D_9), .O(D_9_NOT) );
inv1 gate( .a(N416), .O(N416_NOT) );
and2 gate( .a(N416), .b(D_8_NOT), .O(ED_40) );
and2 gate( .a(N416_NOT), .b(D_8_NOT), .O(ED_41) );
and2 gate( .a(CONST1), .b(D_8), .O(ED_42) );
and2 gate( .a(CONST0), .b(D_8), .O(ED_43) );
and2 gate( .a(ED_40), .b(D_9_NOT), .O(ED_49) );
and2 gate( .a(ED_41), .b(D_9), .O(ED_47) );
and2 gate( .a(ED_42), .b(D_9_NOT), .O(ED_45) );
and2 gate( .a(ED_43), .b(D_9), .O(ED_44) );
or2  gate( .a(ED_44), .b(ED_45), .O(ED_46) );
or2  gate( .a(ED_46), .b(ED_47), .O(ED_48) );
or2  gate( .a(ED_49), .b(ED_48), .O(N416_OBF) );
inv1 gate( .a(D_10), .O(D_10_NOT) );
inv1 gate( .a(D_11), .O(D_11_NOT) );
inv1 gate( .a(N213), .O(N213_NOT) );
and2 gate( .a(N213), .b(D_10_NOT), .O(ED_50) );
and2 gate( .a(N213_NOT), .b(D_10_NOT), .O(ED_51) );
and2 gate( .a(CONST1), .b(D_10), .O(ED_52) );
and2 gate( .a(CONST0), .b(D_10), .O(ED_53) );
and2 gate( .a(ED_50), .b(D_11_NOT), .O(ED_59) );
and2 gate( .a(ED_51), .b(D_11), .O(ED_57) );
and2 gate( .a(ED_52), .b(D_11_NOT), .O(ED_55) );
and2 gate( .a(ED_53), .b(D_11), .O(ED_54) );
or2  gate( .a(ED_54), .b(ED_55), .O(ED_56) );
or2  gate( .a(ED_56), .b(ED_57), .O(ED_58) );
or2  gate( .a(ED_59), .b(ED_58), .O(N213_OBF) );
inv1 gate( .a(D_12), .O(D_12_NOT) );
inv1 gate( .a(D_13), .O(D_13_NOT) );
inv1 gate( .a(N30), .O(N30_NOT) );
and2 gate( .a(N30), .b(D_12_NOT), .O(ED_60) );
and2 gate( .a(N30_NOT), .b(D_12_NOT), .O(ED_61) );
and2 gate( .a(CONST1), .b(D_12), .O(ED_62) );
and2 gate( .a(CONST0), .b(D_12), .O(ED_63) );
and2 gate( .a(ED_60), .b(D_13_NOT), .O(ED_69) );
and2 gate( .a(ED_61), .b(D_13), .O(ED_67) );
and2 gate( .a(ED_62), .b(D_13_NOT), .O(ED_65) );
and2 gate( .a(ED_63), .b(D_13), .O(ED_64) );
or2  gate( .a(ED_64), .b(ED_65), .O(ED_66) );
or2  gate( .a(ED_66), .b(ED_67), .O(ED_68) );
or2  gate( .a(ED_69), .b(ED_68), .O(N30_OBF) );
inv1 gate( .a(D_14), .O(D_14_NOT) );
inv1 gate( .a(D_15), .O(D_15_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_14_NOT), .O(ED_70) );
and2 gate( .a(N360_NOT), .b(D_14_NOT), .O(ED_71) );
and2 gate( .a(CONST1), .b(D_14), .O(ED_72) );
and2 gate( .a(CONST0), .b(D_14), .O(ED_73) );
and2 gate( .a(ED_70), .b(D_15_NOT), .O(ED_79) );
and2 gate( .a(ED_71), .b(D_15), .O(ED_77) );
and2 gate( .a(ED_72), .b(D_15_NOT), .O(ED_75) );
and2 gate( .a(ED_73), .b(D_15), .O(ED_74) );
or2  gate( .a(ED_74), .b(ED_75), .O(ED_76) );
or2  gate( .a(ED_76), .b(ED_77), .O(ED_78) );
or2  gate( .a(ED_79), .b(ED_78), .O(N360_OBF) );
inv1 gate( .a(D_16), .O(D_16_NOT) );
inv1 gate( .a(D_17), .O(D_17_NOT) );
inv1 gate( .a(N99), .O(N99_NOT) );
and2 gate( .a(N99), .b(D_16_NOT), .O(ED_80) );
and2 gate( .a(N99_NOT), .b(D_16_NOT), .O(ED_81) );
and2 gate( .a(CONST1), .b(D_16), .O(ED_82) );
and2 gate( .a(CONST0), .b(D_16), .O(ED_83) );
and2 gate( .a(ED_80), .b(D_17_NOT), .O(ED_89) );
and2 gate( .a(ED_81), .b(D_17), .O(ED_87) );
and2 gate( .a(ED_82), .b(D_17_NOT), .O(ED_85) );
and2 gate( .a(ED_83), .b(D_17), .O(ED_84) );
or2  gate( .a(ED_84), .b(ED_85), .O(ED_86) );
or2  gate( .a(ED_86), .b(ED_87), .O(ED_88) );
or2  gate( .a(ED_89), .b(ED_88), .O(N99_OBF) );
inv1 gate( .a(D_18), .O(D_18_NOT) );
inv1 gate( .a(D_19), .O(D_19_NOT) );
inv1 gate( .a(N296), .O(N296_NOT) );
and2 gate( .a(N296), .b(D_18_NOT), .O(ED_90) );
and2 gate( .a(N296_NOT), .b(D_18_NOT), .O(ED_91) );
and2 gate( .a(CONST1), .b(D_18), .O(ED_92) );
and2 gate( .a(CONST0), .b(D_18), .O(ED_93) );
and2 gate( .a(ED_90), .b(D_19_NOT), .O(ED_99) );
and2 gate( .a(ED_91), .b(D_19), .O(ED_97) );
and2 gate( .a(ED_92), .b(D_19_NOT), .O(ED_95) );
and2 gate( .a(ED_93), .b(D_19), .O(ED_94) );
or2  gate( .a(ED_94), .b(ED_95), .O(ED_96) );
or2  gate( .a(ED_96), .b(ED_97), .O(ED_98) );
or2  gate( .a(ED_99), .b(ED_98), .O(N296_OBF) );
inv1 gate( .a(D_20), .O(D_20_NOT) );
inv1 gate( .a(D_21), .O(D_21_NOT) );
inv1 gate( .a(N95), .O(N95_NOT) );
and2 gate( .a(N95), .b(D_20_NOT), .O(ED_100) );
and2 gate( .a(N95_NOT), .b(D_20_NOT), .O(ED_101) );
and2 gate( .a(CONST1), .b(D_20), .O(ED_102) );
and2 gate( .a(CONST0), .b(D_20), .O(ED_103) );
and2 gate( .a(ED_100), .b(D_21_NOT), .O(ED_109) );
and2 gate( .a(ED_101), .b(D_21), .O(ED_107) );
and2 gate( .a(ED_102), .b(D_21_NOT), .O(ED_105) );
and2 gate( .a(ED_103), .b(D_21), .O(ED_104) );
or2  gate( .a(ED_104), .b(ED_105), .O(ED_106) );
or2  gate( .a(ED_106), .b(ED_107), .O(ED_108) );
or2  gate( .a(ED_109), .b(ED_108), .O(N95_OBF) );
inv1 gate( .a(D_22), .O(D_22_NOT) );
inv1 gate( .a(D_23), .O(D_23_NOT) );
inv1 gate( .a(N357), .O(N357_NOT) );
and2 gate( .a(N357), .b(D_22_NOT), .O(ED_110) );
and2 gate( .a(N357_NOT), .b(D_22_NOT), .O(ED_111) );
and2 gate( .a(CONST1), .b(D_22), .O(ED_112) );
and2 gate( .a(CONST0), .b(D_22), .O(ED_113) );
and2 gate( .a(ED_110), .b(D_23_NOT), .O(ED_119) );
and2 gate( .a(ED_111), .b(D_23), .O(ED_117) );
and2 gate( .a(ED_112), .b(D_23_NOT), .O(ED_115) );
and2 gate( .a(ED_113), .b(D_23), .O(ED_114) );
or2  gate( .a(ED_114), .b(ED_115), .O(ED_116) );
or2  gate( .a(ED_116), .b(ED_117), .O(ED_118) );
or2  gate( .a(ED_119), .b(ED_118), .O(N357_OBF) );
inv1 gate( .a(D_24), .O(D_24_NOT) );
inv1 gate( .a(D_25), .O(D_25_NOT) );
inv1 gate( .a(N50), .O(N50_NOT) );
and2 gate( .a(N50), .b(D_24_NOT), .O(ED_120) );
and2 gate( .a(N50_NOT), .b(D_24_NOT), .O(ED_121) );
and2 gate( .a(CONST1), .b(D_24), .O(ED_122) );
and2 gate( .a(CONST0), .b(D_24), .O(ED_123) );
and2 gate( .a(ED_120), .b(D_25_NOT), .O(ED_129) );
and2 gate( .a(ED_121), .b(D_25), .O(ED_127) );
and2 gate( .a(ED_122), .b(D_25_NOT), .O(ED_125) );
and2 gate( .a(ED_123), .b(D_25), .O(ED_124) );
or2  gate( .a(ED_124), .b(ED_125), .O(ED_126) );
or2  gate( .a(ED_126), .b(ED_127), .O(ED_128) );
or2  gate( .a(ED_129), .b(ED_128), .O(N50_OBF) );
inv1 gate( .a(D_26), .O(D_26_NOT) );
inv1 gate( .a(D_27), .O(D_27_NOT) );
inv1 gate( .a(N341), .O(N341_NOT) );
and2 gate( .a(N341), .b(D_26_NOT), .O(ED_130) );
and2 gate( .a(N341_NOT), .b(D_26_NOT), .O(ED_131) );
and2 gate( .a(CONST1), .b(D_26), .O(ED_132) );
and2 gate( .a(CONST0), .b(D_26), .O(ED_133) );
and2 gate( .a(ED_130), .b(D_27_NOT), .O(ED_139) );
and2 gate( .a(ED_131), .b(D_27), .O(ED_137) );
and2 gate( .a(ED_132), .b(D_27_NOT), .O(ED_135) );
and2 gate( .a(ED_133), .b(D_27), .O(ED_134) );
or2  gate( .a(ED_134), .b(ED_135), .O(ED_136) );
or2  gate( .a(ED_136), .b(ED_137), .O(ED_138) );
or2  gate( .a(ED_139), .b(ED_138), .O(N341_OBF) );
inv1 gate( .a(D_28), .O(D_28_NOT) );
inv1 gate( .a(D_29), .O(D_29_NOT) );
inv1 gate( .a(N267), .O(N267_NOT) );
and2 gate( .a(N267), .b(D_28_NOT), .O(ED_140) );
and2 gate( .a(N267_NOT), .b(D_28_NOT), .O(ED_141) );
and2 gate( .a(CONST1), .b(D_28), .O(ED_142) );
and2 gate( .a(CONST0), .b(D_28), .O(ED_143) );
and2 gate( .a(ED_140), .b(D_29_NOT), .O(ED_149) );
and2 gate( .a(ED_141), .b(D_29), .O(ED_147) );
and2 gate( .a(ED_142), .b(D_29_NOT), .O(ED_145) );
and2 gate( .a(ED_143), .b(D_29), .O(ED_144) );
or2  gate( .a(ED_144), .b(ED_145), .O(ED_146) );
or2  gate( .a(ED_146), .b(ED_147), .O(ED_148) );
or2  gate( .a(ED_149), .b(ED_148), .O(N267_OBF) );
inv1 gate( .a(D_30), .O(D_30_NOT) );
inv1 gate( .a(D_31), .O(D_31_NOT) );
inv1 gate( .a(N254), .O(N254_NOT) );
and2 gate( .a(N254), .b(D_30_NOT), .O(ED_150) );
and2 gate( .a(N254_NOT), .b(D_30_NOT), .O(ED_151) );
and2 gate( .a(CONST1), .b(D_30), .O(ED_152) );
and2 gate( .a(CONST0), .b(D_30), .O(ED_153) );
and2 gate( .a(ED_150), .b(D_31_NOT), .O(ED_159) );
and2 gate( .a(ED_151), .b(D_31), .O(ED_157) );
and2 gate( .a(ED_152), .b(D_31_NOT), .O(ED_155) );
and2 gate( .a(ED_153), .b(D_31), .O(ED_154) );
or2  gate( .a(ED_154), .b(ED_155), .O(ED_156) );
or2  gate( .a(ED_156), .b(ED_157), .O(ED_158) );
or2  gate( .a(ED_159), .b(ED_158), .O(N254_OBF) );
inv1 gate( .a(D_32), .O(D_32_NOT) );
inv1 gate( .a(D_33), .O(D_33_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_32_NOT), .O(ED_160) );
and2 gate( .a(N360_NOT), .b(D_32_NOT), .O(ED_161) );
and2 gate( .a(CONST1), .b(D_32), .O(ED_162) );
and2 gate( .a(CONST0), .b(D_32), .O(ED_163) );
and2 gate( .a(ED_160), .b(D_33_NOT), .O(ED_169) );
and2 gate( .a(ED_161), .b(D_33), .O(ED_167) );
and2 gate( .a(ED_162), .b(D_33_NOT), .O(ED_165) );
and2 gate( .a(ED_163), .b(D_33), .O(ED_164) );
or2  gate( .a(ED_164), .b(ED_165), .O(ED_166) );
or2  gate( .a(ED_166), .b(ED_167), .O(ED_168) );
or2  gate( .a(ED_169), .b(ED_168), .O(N360_OBF) );
inv1 gate( .a(D_34), .O(D_34_NOT) );
inv1 gate( .a(D_35), .O(D_35_NOT) );
inv1 gate( .a(N196), .O(N196_NOT) );
and2 gate( .a(N196), .b(D_34_NOT), .O(ED_170) );
and2 gate( .a(N196_NOT), .b(D_34_NOT), .O(ED_171) );
and2 gate( .a(CONST1), .b(D_34), .O(ED_172) );
and2 gate( .a(CONST0), .b(D_34), .O(ED_173) );
and2 gate( .a(ED_170), .b(D_35_NOT), .O(ED_179) );
and2 gate( .a(ED_171), .b(D_35), .O(ED_177) );
and2 gate( .a(ED_172), .b(D_35_NOT), .O(ED_175) );
and2 gate( .a(ED_173), .b(D_35), .O(ED_174) );
or2  gate( .a(ED_174), .b(ED_175), .O(ED_176) );
or2  gate( .a(ED_176), .b(ED_177), .O(ED_178) );
or2  gate( .a(ED_179), .b(ED_178), .O(N196_OBF) );
inv1 gate( .a(D_36), .O(D_36_NOT) );
inv1 gate( .a(D_37), .O(D_37_NOT) );
inv1 gate( .a(N197), .O(N197_NOT) );
and2 gate( .a(N197), .b(D_36_NOT), .O(ED_180) );
and2 gate( .a(N197_NOT), .b(D_36_NOT), .O(ED_181) );
and2 gate( .a(CONST1), .b(D_36), .O(ED_182) );
and2 gate( .a(CONST0), .b(D_36), .O(ED_183) );
and2 gate( .a(ED_180), .b(D_37_NOT), .O(ED_189) );
and2 gate( .a(ED_181), .b(D_37), .O(ED_187) );
and2 gate( .a(ED_182), .b(D_37_NOT), .O(ED_185) );
and2 gate( .a(ED_183), .b(D_37), .O(ED_184) );
or2  gate( .a(ED_184), .b(ED_185), .O(ED_186) );
or2  gate( .a(ED_186), .b(ED_187), .O(ED_188) );
or2  gate( .a(ED_189), .b(ED_188), .O(N197_OBF) );
inv1 gate( .a(D_38), .O(D_38_NOT) );
inv1 gate( .a(D_39), .O(D_39_NOT) );
inv1 gate( .a(N157), .O(N157_NOT) );
and2 gate( .a(N157), .b(D_38_NOT), .O(ED_190) );
and2 gate( .a(N157_NOT), .b(D_38_NOT), .O(ED_191) );
and2 gate( .a(CONST1), .b(D_38), .O(ED_192) );
and2 gate( .a(CONST0), .b(D_38), .O(ED_193) );
and2 gate( .a(ED_190), .b(D_39_NOT), .O(ED_199) );
and2 gate( .a(ED_191), .b(D_39), .O(ED_197) );
and2 gate( .a(ED_192), .b(D_39_NOT), .O(ED_195) );
and2 gate( .a(ED_193), .b(D_39), .O(ED_194) );
or2  gate( .a(ED_194), .b(ED_195), .O(ED_196) );
or2  gate( .a(ED_196), .b(ED_197), .O(ED_198) );
or2  gate( .a(ED_199), .b(ED_198), .O(N157_OBF) );
inv1 gate( .a(D_40), .O(D_40_NOT) );
inv1 gate( .a(D_41), .O(D_41_NOT) );
inv1 gate( .a(N50), .O(N50_NOT) );
and2 gate( .a(N50), .b(D_40_NOT), .O(ED_200) );
and2 gate( .a(N50_NOT), .b(D_40_NOT), .O(ED_201) );
and2 gate( .a(CONST1), .b(D_40), .O(ED_202) );
and2 gate( .a(CONST0), .b(D_40), .O(ED_203) );
and2 gate( .a(ED_200), .b(D_41_NOT), .O(ED_209) );
and2 gate( .a(ED_201), .b(D_41), .O(ED_207) );
and2 gate( .a(ED_202), .b(D_41_NOT), .O(ED_205) );
and2 gate( .a(ED_203), .b(D_41), .O(ED_204) );
or2  gate( .a(ED_204), .b(ED_205), .O(ED_206) );
or2  gate( .a(ED_206), .b(ED_207), .O(ED_208) );
or2  gate( .a(ED_209), .b(ED_208), .O(N50_OBF) );
inv1 gate( .a(D_42), .O(D_42_NOT) );
inv1 gate( .a(D_43), .O(D_43_NOT) );
inv1 gate( .a(N123), .O(N123_NOT) );
and2 gate( .a(N123), .b(D_42_NOT), .O(ED_210) );
and2 gate( .a(N123_NOT), .b(D_42_NOT), .O(ED_211) );
and2 gate( .a(CONST1), .b(D_42), .O(ED_212) );
and2 gate( .a(CONST0), .b(D_42), .O(ED_213) );
and2 gate( .a(ED_210), .b(D_43_NOT), .O(ED_219) );
and2 gate( .a(ED_211), .b(D_43), .O(ED_217) );
and2 gate( .a(ED_212), .b(D_43_NOT), .O(ED_215) );
and2 gate( .a(ED_213), .b(D_43), .O(ED_214) );
or2  gate( .a(ED_214), .b(ED_215), .O(ED_216) );
or2  gate( .a(ED_216), .b(ED_217), .O(ED_218) );
or2  gate( .a(ED_219), .b(ED_218), .O(N123_OBF) );
inv1 gate( .a(D_44), .O(D_44_NOT) );
inv1 gate( .a(D_45), .O(D_45_NOT) );
inv1 gate( .a(N105), .O(N105_NOT) );
and2 gate( .a(N105), .b(D_44_NOT), .O(ED_220) );
and2 gate( .a(N105_NOT), .b(D_44_NOT), .O(ED_221) );
and2 gate( .a(CONST1), .b(D_44), .O(ED_222) );
and2 gate( .a(CONST0), .b(D_44), .O(ED_223) );
and2 gate( .a(ED_220), .b(D_45_NOT), .O(ED_229) );
and2 gate( .a(ED_221), .b(D_45), .O(ED_227) );
and2 gate( .a(ED_222), .b(D_45_NOT), .O(ED_225) );
and2 gate( .a(ED_223), .b(D_45), .O(ED_224) );
or2  gate( .a(ED_224), .b(ED_225), .O(ED_226) );
or2  gate( .a(ED_226), .b(ED_227), .O(ED_228) );
or2  gate( .a(ED_229), .b(ED_228), .O(N105_OBF) );
inv1 gate( .a(D_46), .O(D_46_NOT) );
inv1 gate( .a(D_47), .O(D_47_NOT) );
inv1 gate( .a(N102), .O(N102_NOT) );
and2 gate( .a(N102), .b(D_46_NOT), .O(ED_230) );
and2 gate( .a(N102_NOT), .b(D_46_NOT), .O(ED_231) );
and2 gate( .a(CONST1), .b(D_46), .O(ED_232) );
and2 gate( .a(CONST0), .b(D_46), .O(ED_233) );
and2 gate( .a(ED_230), .b(D_47_NOT), .O(ED_239) );
and2 gate( .a(ED_231), .b(D_47), .O(ED_237) );
and2 gate( .a(ED_232), .b(D_47_NOT), .O(ED_235) );
and2 gate( .a(ED_233), .b(D_47), .O(ED_234) );
or2  gate( .a(ED_234), .b(ED_235), .O(ED_236) );
or2  gate( .a(ED_236), .b(ED_237), .O(ED_238) );
or2  gate( .a(ED_239), .b(ED_238), .O(N102_OBF) );
inv1 gate( .a(D_48), .O(D_48_NOT) );
inv1 gate( .a(D_49), .O(D_49_NOT) );
inv1 gate( .a(N95), .O(N95_NOT) );
and2 gate( .a(N95), .b(D_48_NOT), .O(ED_240) );
and2 gate( .a(N95_NOT), .b(D_48_NOT), .O(ED_241) );
and2 gate( .a(CONST1), .b(D_48), .O(ED_242) );
and2 gate( .a(CONST0), .b(D_48), .O(ED_243) );
and2 gate( .a(ED_240), .b(D_49_NOT), .O(ED_249) );
and2 gate( .a(ED_241), .b(D_49), .O(ED_247) );
and2 gate( .a(ED_242), .b(D_49_NOT), .O(ED_245) );
and2 gate( .a(ED_243), .b(D_49), .O(ED_244) );
or2  gate( .a(ED_244), .b(ED_245), .O(ED_246) );
or2  gate( .a(ED_246), .b(ED_247), .O(ED_248) );
or2  gate( .a(ED_249), .b(ED_248), .O(N95_OBF) );
inv1 gate( .a(D_50), .O(D_50_NOT) );
inv1 gate( .a(D_51), .O(D_51_NOT) );
inv1 gate( .a(N139), .O(N139_NOT) );
and2 gate( .a(N139), .b(D_50_NOT), .O(ED_250) );
and2 gate( .a(N139_NOT), .b(D_50_NOT), .O(ED_251) );
and2 gate( .a(CONST1), .b(D_50), .O(ED_252) );
and2 gate( .a(CONST0), .b(D_50), .O(ED_253) );
and2 gate( .a(ED_250), .b(D_51_NOT), .O(ED_259) );
and2 gate( .a(ED_251), .b(D_51), .O(ED_257) );
and2 gate( .a(ED_252), .b(D_51_NOT), .O(ED_255) );
and2 gate( .a(ED_253), .b(D_51), .O(ED_254) );
or2  gate( .a(ED_254), .b(ED_255), .O(ED_256) );
or2  gate( .a(ED_256), .b(ED_257), .O(ED_258) );
or2  gate( .a(ED_259), .b(ED_258), .O(N139_OBF) );
inv1 gate( .a(D_52), .O(D_52_NOT) );
inv1 gate( .a(D_53), .O(D_53_NOT) );
inv1 gate( .a(N295), .O(N295_NOT) );
and2 gate( .a(N295), .b(D_52_NOT), .O(ED_260) );
and2 gate( .a(N295_NOT), .b(D_52_NOT), .O(ED_261) );
and2 gate( .a(CONST1), .b(D_52), .O(ED_262) );
and2 gate( .a(CONST0), .b(D_52), .O(ED_263) );
and2 gate( .a(ED_260), .b(D_53_NOT), .O(ED_269) );
and2 gate( .a(ED_261), .b(D_53), .O(ED_267) );
and2 gate( .a(ED_262), .b(D_53_NOT), .O(ED_265) );
and2 gate( .a(ED_263), .b(D_53), .O(ED_264) );
or2  gate( .a(ED_264), .b(ED_265), .O(ED_266) );
or2  gate( .a(ED_266), .b(ED_267), .O(ED_268) );
or2  gate( .a(ED_269), .b(ED_268), .O(N295_OBF) );
inv1 gate( .a(D_54), .O(D_54_NOT) );
inv1 gate( .a(D_55), .O(D_55_NOT) );
inv1 gate( .a(N131), .O(N131_NOT) );
and2 gate( .a(N131), .b(D_54_NOT), .O(ED_270) );
and2 gate( .a(N131_NOT), .b(D_54_NOT), .O(ED_271) );
and2 gate( .a(CONST1), .b(D_54), .O(ED_272) );
and2 gate( .a(CONST0), .b(D_54), .O(ED_273) );
and2 gate( .a(ED_270), .b(D_55_NOT), .O(ED_279) );
and2 gate( .a(ED_271), .b(D_55), .O(ED_277) );
and2 gate( .a(ED_272), .b(D_55_NOT), .O(ED_275) );
and2 gate( .a(ED_273), .b(D_55), .O(ED_274) );
or2  gate( .a(ED_274), .b(ED_275), .O(ED_276) );
or2  gate( .a(ED_276), .b(ED_277), .O(ED_278) );
or2  gate( .a(ED_279), .b(ED_278), .O(N131_OBF) );
inv1 gate( .a(D_56), .O(D_56_NOT) );
inv1 gate( .a(D_57), .O(D_57_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_56_NOT), .O(ED_280) );
and2 gate( .a(N360_NOT), .b(D_56_NOT), .O(ED_281) );
and2 gate( .a(CONST1), .b(D_56), .O(ED_282) );
and2 gate( .a(CONST0), .b(D_56), .O(ED_283) );
and2 gate( .a(ED_280), .b(D_57_NOT), .O(ED_289) );
and2 gate( .a(ED_281), .b(D_57), .O(ED_287) );
and2 gate( .a(ED_282), .b(D_57_NOT), .O(ED_285) );
and2 gate( .a(ED_283), .b(D_57), .O(ED_284) );
or2  gate( .a(ED_284), .b(ED_285), .O(ED_286) );
or2  gate( .a(ED_286), .b(ED_287), .O(ED_288) );
or2  gate( .a(ED_289), .b(ED_288), .O(N360_OBF) );
inv1 gate( .a(D_58), .O(D_58_NOT) );
inv1 gate( .a(D_59), .O(D_59_NOT) );
inv1 gate( .a(N334), .O(N334_NOT) );
and2 gate( .a(N334), .b(D_58_NOT), .O(ED_290) );
and2 gate( .a(N334_NOT), .b(D_58_NOT), .O(ED_291) );
and2 gate( .a(CONST1), .b(D_58), .O(ED_292) );
and2 gate( .a(CONST0), .b(D_58), .O(ED_293) );
and2 gate( .a(ED_290), .b(D_59_NOT), .O(ED_299) );
and2 gate( .a(ED_291), .b(D_59), .O(ED_297) );
and2 gate( .a(ED_292), .b(D_59_NOT), .O(ED_295) );
and2 gate( .a(ED_293), .b(D_59), .O(ED_294) );
or2  gate( .a(ED_294), .b(ED_295), .O(ED_296) );
or2  gate( .a(ED_296), .b(ED_297), .O(ED_298) );
or2  gate( .a(ED_299), .b(ED_298), .O(N334_OBF) );
inv1 gate( .a(D_60), .O(D_60_NOT) );
inv1 gate( .a(D_61), .O(D_61_NOT) );
inv1 gate( .a(N292), .O(N292_NOT) );
and2 gate( .a(N292), .b(D_60_NOT), .O(ED_300) );
and2 gate( .a(N292_NOT), .b(D_60_NOT), .O(ED_301) );
and2 gate( .a(CONST1), .b(D_60), .O(ED_302) );
and2 gate( .a(CONST0), .b(D_60), .O(ED_303) );
and2 gate( .a(ED_300), .b(D_61_NOT), .O(ED_309) );
and2 gate( .a(ED_301), .b(D_61), .O(ED_307) );
and2 gate( .a(ED_302), .b(D_61_NOT), .O(ED_305) );
and2 gate( .a(ED_303), .b(D_61), .O(ED_304) );
or2  gate( .a(ED_304), .b(ED_305), .O(ED_306) );
or2  gate( .a(ED_306), .b(ED_307), .O(ED_308) );
or2  gate( .a(ED_309), .b(ED_308), .O(N292_OBF) );
inv1 gate( .a(D_62), .O(D_62_NOT) );
inv1 gate( .a(D_63), .O(D_63_NOT) );
inv1 gate( .a(N199), .O(N199_NOT) );
and2 gate( .a(N199), .b(D_62_NOT), .O(ED_310) );
and2 gate( .a(N199_NOT), .b(D_62_NOT), .O(ED_311) );
and2 gate( .a(CONST1), .b(D_62), .O(ED_312) );
and2 gate( .a(CONST0), .b(D_62), .O(ED_313) );
and2 gate( .a(ED_310), .b(D_63_NOT), .O(ED_319) );
and2 gate( .a(ED_311), .b(D_63), .O(ED_317) );
and2 gate( .a(ED_312), .b(D_63_NOT), .O(ED_315) );
and2 gate( .a(ED_313), .b(D_63), .O(ED_314) );
or2  gate( .a(ED_314), .b(ED_315), .O(ED_316) );
or2  gate( .a(ED_316), .b(ED_317), .O(ED_318) );
or2  gate( .a(ED_319), .b(ED_318), .O(N199_OBF) );
inv1 gate( .a(D_64), .O(D_64_NOT) );
inv1 gate( .a(D_65), .O(D_65_NOT) );
inv1 gate( .a(N112), .O(N112_NOT) );
and2 gate( .a(N112), .b(D_64_NOT), .O(ED_320) );
and2 gate( .a(N112_NOT), .b(D_64_NOT), .O(ED_321) );
and2 gate( .a(CONST1), .b(D_64), .O(ED_322) );
and2 gate( .a(CONST0), .b(D_64), .O(ED_323) );
and2 gate( .a(ED_320), .b(D_65_NOT), .O(ED_329) );
and2 gate( .a(ED_321), .b(D_65), .O(ED_327) );
and2 gate( .a(ED_322), .b(D_65_NOT), .O(ED_325) );
and2 gate( .a(ED_323), .b(D_65), .O(ED_324) );
or2  gate( .a(ED_324), .b(ED_325), .O(ED_326) );
or2  gate( .a(ED_326), .b(ED_327), .O(ED_328) );
or2  gate( .a(ED_329), .b(ED_328), .O(N112_OBF) );
inv1 gate( .a(D_66), .O(D_66_NOT) );
inv1 gate( .a(D_67), .O(D_67_NOT) );
inv1 gate( .a(N243), .O(N243_NOT) );
and2 gate( .a(N243), .b(D_66_NOT), .O(ED_330) );
and2 gate( .a(N243_NOT), .b(D_66_NOT), .O(ED_331) );
and2 gate( .a(CONST1), .b(D_66), .O(ED_332) );
and2 gate( .a(CONST0), .b(D_66), .O(ED_333) );
and2 gate( .a(ED_330), .b(D_67_NOT), .O(ED_339) );
and2 gate( .a(ED_331), .b(D_67), .O(ED_337) );
and2 gate( .a(ED_332), .b(D_67_NOT), .O(ED_335) );
and2 gate( .a(ED_333), .b(D_67), .O(ED_334) );
or2  gate( .a(ED_334), .b(ED_335), .O(ED_336) );
or2  gate( .a(ED_336), .b(ED_337), .O(ED_338) );
or2  gate( .a(ED_339), .b(ED_338), .O(N243_OBF) );
inv1 gate( .a(D_68), .O(D_68_NOT) );
inv1 gate( .a(D_69), .O(D_69_NOT) );
inv1 gate( .a(N131), .O(N131_NOT) );
and2 gate( .a(N131), .b(D_68_NOT), .O(ED_340) );
and2 gate( .a(N131_NOT), .b(D_68_NOT), .O(ED_341) );
and2 gate( .a(CONST1), .b(D_68), .O(ED_342) );
and2 gate( .a(CONST0), .b(D_68), .O(ED_343) );
and2 gate( .a(ED_340), .b(D_69_NOT), .O(ED_349) );
and2 gate( .a(ED_341), .b(D_69), .O(ED_347) );
and2 gate( .a(ED_342), .b(D_69_NOT), .O(ED_345) );
and2 gate( .a(ED_343), .b(D_69), .O(ED_344) );
or2  gate( .a(ED_344), .b(ED_345), .O(ED_346) );
or2  gate( .a(ED_346), .b(ED_347), .O(ED_348) );
or2  gate( .a(ED_349), .b(ED_348), .O(N131_OBF) );
inv1 gate( .a(D_70), .O(D_70_NOT) );
inv1 gate( .a(D_71), .O(D_71_NOT) );
inv1 gate( .a(N191), .O(N191_NOT) );
and2 gate( .a(N191), .b(D_70_NOT), .O(ED_350) );
and2 gate( .a(N191_NOT), .b(D_70_NOT), .O(ED_351) );
and2 gate( .a(CONST1), .b(D_70), .O(ED_352) );
and2 gate( .a(CONST0), .b(D_70), .O(ED_353) );
and2 gate( .a(ED_350), .b(D_71_NOT), .O(ED_359) );
and2 gate( .a(ED_351), .b(D_71), .O(ED_357) );
and2 gate( .a(ED_352), .b(D_71_NOT), .O(ED_355) );
and2 gate( .a(ED_353), .b(D_71), .O(ED_354) );
or2  gate( .a(ED_354), .b(ED_355), .O(ED_356) );
or2  gate( .a(ED_356), .b(ED_357), .O(ED_358) );
or2  gate( .a(ED_359), .b(ED_358), .O(N191_OBF) );
inv1 gate( .a(D_72), .O(D_72_NOT) );
inv1 gate( .a(D_73), .O(D_73_NOT) );
inv1 gate( .a(N345), .O(N345_NOT) );
and2 gate( .a(N345), .b(D_72_NOT), .O(ED_360) );
and2 gate( .a(N345_NOT), .b(D_72_NOT), .O(ED_361) );
and2 gate( .a(CONST1), .b(D_72), .O(ED_362) );
and2 gate( .a(CONST0), .b(D_72), .O(ED_363) );
and2 gate( .a(ED_360), .b(D_73_NOT), .O(ED_369) );
and2 gate( .a(ED_361), .b(D_73), .O(ED_367) );
and2 gate( .a(ED_362), .b(D_73_NOT), .O(ED_365) );
and2 gate( .a(ED_363), .b(D_73), .O(ED_364) );
or2  gate( .a(ED_364), .b(ED_365), .O(ED_366) );
or2  gate( .a(ED_366), .b(ED_367), .O(ED_368) );
or2  gate( .a(ED_369), .b(ED_368), .O(N345_OBF) );
inv1 gate( .a(D_74), .O(D_74_NOT) );
inv1 gate( .a(D_75), .O(D_75_NOT) );
inv1 gate( .a(N213), .O(N213_NOT) );
and2 gate( .a(N213), .b(D_74_NOT), .O(ED_370) );
and2 gate( .a(N213_NOT), .b(D_74_NOT), .O(ED_371) );
and2 gate( .a(CONST1), .b(D_74), .O(ED_372) );
and2 gate( .a(CONST0), .b(D_74), .O(ED_373) );
and2 gate( .a(ED_370), .b(D_75_NOT), .O(ED_379) );
and2 gate( .a(ED_371), .b(D_75), .O(ED_377) );
and2 gate( .a(ED_372), .b(D_75_NOT), .O(ED_375) );
and2 gate( .a(ED_373), .b(D_75), .O(ED_374) );
or2  gate( .a(ED_374), .b(ED_375), .O(ED_376) );
or2  gate( .a(ED_376), .b(ED_377), .O(ED_378) );
or2  gate( .a(ED_379), .b(ED_378), .O(N213_OBF) );
inv1 gate( .a(D_76), .O(D_76_NOT) );
inv1 gate( .a(D_77), .O(D_77_NOT) );
inv1 gate( .a(N1), .O(N1_NOT) );
and2 gate( .a(N1), .b(D_76_NOT), .O(ED_380) );
and2 gate( .a(N1_NOT), .b(D_76_NOT), .O(ED_381) );
and2 gate( .a(CONST1), .b(D_76), .O(ED_382) );
and2 gate( .a(CONST0), .b(D_76), .O(ED_383) );
and2 gate( .a(ED_380), .b(D_77_NOT), .O(ED_389) );
and2 gate( .a(ED_381), .b(D_77), .O(ED_387) );
and2 gate( .a(ED_382), .b(D_77_NOT), .O(ED_385) );
and2 gate( .a(ED_383), .b(D_77), .O(ED_384) );
or2  gate( .a(ED_384), .b(ED_385), .O(ED_386) );
or2  gate( .a(ED_386), .b(ED_387), .O(ED_388) );
or2  gate( .a(ED_389), .b(ED_388), .O(N1_OBF) );
inv1 gate( .a(D_78), .O(D_78_NOT) );
inv1 gate( .a(D_79), .O(D_79_NOT) );
inv1 gate( .a(N420), .O(N420_NOT) );
and2 gate( .a(N420), .b(D_78_NOT), .O(ED_390) );
and2 gate( .a(N420_NOT), .b(D_78_NOT), .O(ED_391) );
and2 gate( .a(CONST1), .b(D_78), .O(ED_392) );
and2 gate( .a(CONST0), .b(D_78), .O(ED_393) );
and2 gate( .a(ED_390), .b(D_79_NOT), .O(ED_399) );
and2 gate( .a(ED_391), .b(D_79), .O(ED_397) );
and2 gate( .a(ED_392), .b(D_79_NOT), .O(ED_395) );
and2 gate( .a(ED_393), .b(D_79), .O(ED_394) );
or2  gate( .a(ED_394), .b(ED_395), .O(ED_396) );
or2  gate( .a(ED_396), .b(ED_397), .O(ED_398) );
or2  gate( .a(ED_399), .b(ED_398), .O(N420_OBF) );
inv1 gate( .a(D_80), .O(D_80_NOT) );
inv1 gate( .a(D_81), .O(D_81_NOT) );
inv1 gate( .a(N319), .O(N319_NOT) );
and2 gate( .a(N319), .b(D_80_NOT), .O(ED_400) );
and2 gate( .a(N319_NOT), .b(D_80_NOT), .O(ED_401) );
and2 gate( .a(CONST1), .b(D_80), .O(ED_402) );
and2 gate( .a(CONST0), .b(D_80), .O(ED_403) );
and2 gate( .a(ED_400), .b(D_81_NOT), .O(ED_409) );
and2 gate( .a(ED_401), .b(D_81), .O(ED_407) );
and2 gate( .a(ED_402), .b(D_81_NOT), .O(ED_405) );
and2 gate( .a(ED_403), .b(D_81), .O(ED_404) );
or2  gate( .a(ED_404), .b(ED_405), .O(ED_406) );
or2  gate( .a(ED_406), .b(ED_407), .O(ED_408) );
or2  gate( .a(ED_409), .b(ED_408), .O(N319_OBF) );
inv1 gate( .a(D_82), .O(D_82_NOT) );
inv1 gate( .a(D_83), .O(D_83_NOT) );
inv1 gate( .a(N294), .O(N294_NOT) );
and2 gate( .a(N294), .b(D_82_NOT), .O(ED_410) );
and2 gate( .a(N294_NOT), .b(D_82_NOT), .O(ED_411) );
and2 gate( .a(CONST1), .b(D_82), .O(ED_412) );
and2 gate( .a(CONST0), .b(D_82), .O(ED_413) );
and2 gate( .a(ED_410), .b(D_83_NOT), .O(ED_419) );
and2 gate( .a(ED_411), .b(D_83), .O(ED_417) );
and2 gate( .a(ED_412), .b(D_83_NOT), .O(ED_415) );
and2 gate( .a(ED_413), .b(D_83), .O(ED_414) );
or2  gate( .a(ED_414), .b(ED_415), .O(ED_416) );
or2  gate( .a(ED_416), .b(ED_417), .O(ED_418) );
or2  gate( .a(ED_419), .b(ED_418), .O(N294_OBF) );
inv1 gate( .a(D_84), .O(D_84_NOT) );
inv1 gate( .a(D_85), .O(D_85_NOT) );
inv1 gate( .a(N422), .O(N422_NOT) );
and2 gate( .a(N422), .b(D_84_NOT), .O(ED_420) );
and2 gate( .a(N422_NOT), .b(D_84_NOT), .O(ED_421) );
and2 gate( .a(CONST1), .b(D_84), .O(ED_422) );
and2 gate( .a(CONST0), .b(D_84), .O(ED_423) );
and2 gate( .a(ED_420), .b(D_85_NOT), .O(ED_429) );
and2 gate( .a(ED_421), .b(D_85), .O(ED_427) );
and2 gate( .a(ED_422), .b(D_85_NOT), .O(ED_425) );
and2 gate( .a(ED_423), .b(D_85), .O(ED_424) );
or2  gate( .a(ED_424), .b(ED_425), .O(ED_426) );
or2  gate( .a(ED_426), .b(ED_427), .O(ED_428) );
or2  gate( .a(ED_429), .b(ED_428), .O(N422_OBF) );
inv1 gate( .a(D_86), .O(D_86_NOT) );
inv1 gate( .a(D_87), .O(D_87_NOT) );
inv1 gate( .a(N4), .O(N4_NOT) );
and2 gate( .a(N4), .b(D_86_NOT), .O(ED_430) );
and2 gate( .a(N4_NOT), .b(D_86_NOT), .O(ED_431) );
and2 gate( .a(CONST1), .b(D_86), .O(ED_432) );
and2 gate( .a(CONST0), .b(D_86), .O(ED_433) );
and2 gate( .a(ED_430), .b(D_87_NOT), .O(ED_439) );
and2 gate( .a(ED_431), .b(D_87), .O(ED_437) );
and2 gate( .a(ED_432), .b(D_87_NOT), .O(ED_435) );
and2 gate( .a(ED_433), .b(D_87), .O(ED_434) );
or2  gate( .a(ED_434), .b(ED_435), .O(ED_436) );
or2  gate( .a(ED_436), .b(ED_437), .O(ED_438) );
or2  gate( .a(ED_439), .b(ED_438), .O(N4_OBF) );
inv1 gate( .a(D_88), .O(D_88_NOT) );
inv1 gate( .a(D_89), .O(D_89_NOT) );
inv1 gate( .a(N56), .O(N56_NOT) );
and2 gate( .a(N56), .b(D_88_NOT), .O(ED_440) );
and2 gate( .a(N56_NOT), .b(D_88_NOT), .O(ED_441) );
and2 gate( .a(CONST1), .b(D_88), .O(ED_442) );
and2 gate( .a(CONST0), .b(D_88), .O(ED_443) );
and2 gate( .a(ED_440), .b(D_89_NOT), .O(ED_449) );
and2 gate( .a(ED_441), .b(D_89), .O(ED_447) );
and2 gate( .a(ED_442), .b(D_89_NOT), .O(ED_445) );
and2 gate( .a(ED_443), .b(D_89), .O(ED_444) );
or2  gate( .a(ED_444), .b(ED_445), .O(ED_446) );
or2  gate( .a(ED_446), .b(ED_447), .O(ED_448) );
or2  gate( .a(ED_449), .b(ED_448), .O(N56_OBF) );
inv1 gate( .a(D_90), .O(D_90_NOT) );
inv1 gate( .a(D_91), .O(D_91_NOT) );
inv1 gate( .a(N37), .O(N37_NOT) );
and2 gate( .a(N37), .b(D_90_NOT), .O(ED_450) );
and2 gate( .a(N37_NOT), .b(D_90_NOT), .O(ED_451) );
and2 gate( .a(CONST1), .b(D_90), .O(ED_452) );
and2 gate( .a(CONST0), .b(D_90), .O(ED_453) );
and2 gate( .a(ED_450), .b(D_91_NOT), .O(ED_459) );
and2 gate( .a(ED_451), .b(D_91), .O(ED_457) );
and2 gate( .a(ED_452), .b(D_91_NOT), .O(ED_455) );
and2 gate( .a(ED_453), .b(D_91), .O(ED_454) );
or2  gate( .a(ED_454), .b(ED_455), .O(ED_456) );
or2  gate( .a(ED_456), .b(ED_457), .O(ED_458) );
or2  gate( .a(ED_459), .b(ED_458), .O(N37_OBF) );
inv1 gate( .a(D_92), .O(D_92_NOT) );
inv1 gate( .a(D_93), .O(D_93_NOT) );
inv1 gate( .a(N8), .O(N8_NOT) );
and2 gate( .a(N8), .b(D_92_NOT), .O(ED_460) );
and2 gate( .a(N8_NOT), .b(D_92_NOT), .O(ED_461) );
and2 gate( .a(CONST1), .b(D_92), .O(ED_462) );
and2 gate( .a(CONST0), .b(D_92), .O(ED_463) );
and2 gate( .a(ED_460), .b(D_93_NOT), .O(ED_469) );
and2 gate( .a(ED_461), .b(D_93), .O(ED_467) );
and2 gate( .a(ED_462), .b(D_93_NOT), .O(ED_465) );
and2 gate( .a(ED_463), .b(D_93), .O(ED_464) );
or2  gate( .a(ED_464), .b(ED_465), .O(ED_466) );
or2  gate( .a(ED_466), .b(ED_467), .O(ED_468) );
or2  gate( .a(ED_469), .b(ED_468), .O(N8_OBF) );
inv1 gate( .a(D_94), .O(D_94_NOT) );
inv1 gate( .a(D_95), .O(D_95_NOT) );
inv1 gate( .a(N34), .O(N34_NOT) );
and2 gate( .a(N34), .b(D_94_NOT), .O(ED_470) );
and2 gate( .a(N34_NOT), .b(D_94_NOT), .O(ED_471) );
and2 gate( .a(CONST1), .b(D_94), .O(ED_472) );
and2 gate( .a(CONST0), .b(D_94), .O(ED_473) );
and2 gate( .a(ED_470), .b(D_95_NOT), .O(ED_479) );
and2 gate( .a(ED_471), .b(D_95), .O(ED_477) );
and2 gate( .a(ED_472), .b(D_95_NOT), .O(ED_475) );
and2 gate( .a(ED_473), .b(D_95), .O(ED_474) );
or2  gate( .a(ED_474), .b(ED_475), .O(ED_476) );
or2  gate( .a(ED_476), .b(ED_477), .O(ED_478) );
or2  gate( .a(ED_479), .b(ED_478), .O(N34_OBF) );
inv1 gate( .a(D_96), .O(D_96_NOT) );
inv1 gate( .a(D_97), .O(D_97_NOT) );
inv1 gate( .a(N14), .O(N14_NOT) );
and2 gate( .a(N14), .b(D_96_NOT), .O(ED_480) );
and2 gate( .a(N14_NOT), .b(D_96_NOT), .O(ED_481) );
and2 gate( .a(CONST1), .b(D_96), .O(ED_482) );
and2 gate( .a(CONST0), .b(D_96), .O(ED_483) );
and2 gate( .a(ED_480), .b(D_97_NOT), .O(ED_489) );
and2 gate( .a(ED_481), .b(D_97), .O(ED_487) );
and2 gate( .a(ED_482), .b(D_97_NOT), .O(ED_485) );
and2 gate( .a(ED_483), .b(D_97), .O(ED_484) );
or2  gate( .a(ED_484), .b(ED_485), .O(ED_486) );
or2  gate( .a(ED_486), .b(ED_487), .O(ED_488) );
or2  gate( .a(ED_489), .b(ED_488), .O(N14_OBF) );
inv1 gate( .a(D_98), .O(D_98_NOT) );
inv1 gate( .a(D_99), .O(D_99_NOT) );
inv1 gate( .a(N357), .O(N357_NOT) );
and2 gate( .a(N357), .b(D_98_NOT), .O(ED_490) );
and2 gate( .a(N357_NOT), .b(D_98_NOT), .O(ED_491) );
and2 gate( .a(CONST1), .b(D_98), .O(ED_492) );
and2 gate( .a(CONST0), .b(D_98), .O(ED_493) );
and2 gate( .a(ED_490), .b(D_99_NOT), .O(ED_499) );
and2 gate( .a(ED_491), .b(D_99), .O(ED_497) );
and2 gate( .a(ED_492), .b(D_99_NOT), .O(ED_495) );
and2 gate( .a(ED_493), .b(D_99), .O(ED_494) );
or2  gate( .a(ED_494), .b(ED_495), .O(ED_496) );
or2  gate( .a(ED_496), .b(ED_497), .O(ED_498) );
or2  gate( .a(ED_499), .b(ED_498), .O(N357_OBF) );
inv1 gate( .a(D_100), .O(D_100_NOT) );
inv1 gate( .a(D_101), .O(D_101_NOT) );
inv1 gate( .a(N411), .O(N411_NOT) );
and2 gate( .a(N411), .b(D_100_NOT), .O(ED_500) );
and2 gate( .a(N411_NOT), .b(D_100_NOT), .O(ED_501) );
and2 gate( .a(CONST1), .b(D_100), .O(ED_502) );
and2 gate( .a(CONST0), .b(D_100), .O(ED_503) );
and2 gate( .a(ED_500), .b(D_101_NOT), .O(ED_509) );
and2 gate( .a(ED_501), .b(D_101), .O(ED_507) );
and2 gate( .a(ED_502), .b(D_101_NOT), .O(ED_505) );
and2 gate( .a(ED_503), .b(D_101), .O(ED_504) );
or2  gate( .a(ED_504), .b(ED_505), .O(ED_506) );
or2  gate( .a(ED_506), .b(ED_507), .O(ED_508) );
or2  gate( .a(ED_509), .b(ED_508), .O(N411_OBF) );
inv1 gate( .a(D_102), .O(D_102_NOT) );
inv1 gate( .a(D_103), .O(D_103_NOT) );
inv1 gate( .a(N290), .O(N290_NOT) );
and2 gate( .a(N290), .b(D_102_NOT), .O(ED_510) );
and2 gate( .a(N290_NOT), .b(D_102_NOT), .O(ED_511) );
and2 gate( .a(CONST1), .b(D_102), .O(ED_512) );
and2 gate( .a(CONST0), .b(D_102), .O(ED_513) );
and2 gate( .a(ED_510), .b(D_103_NOT), .O(ED_519) );
and2 gate( .a(ED_511), .b(D_103), .O(ED_517) );
and2 gate( .a(ED_512), .b(D_103_NOT), .O(ED_515) );
and2 gate( .a(ED_513), .b(D_103), .O(ED_514) );
or2  gate( .a(ED_514), .b(ED_515), .O(ED_516) );
or2  gate( .a(ED_516), .b(ED_517), .O(ED_518) );
or2  gate( .a(ED_519), .b(ED_518), .O(N290_OBF) );
inv1 gate( .a(D_104), .O(D_104_NOT) );
inv1 gate( .a(D_105), .O(D_105_NOT) );
inv1 gate( .a(N332), .O(N332_NOT) );
and2 gate( .a(N332), .b(D_104_NOT), .O(ED_520) );
and2 gate( .a(N332_NOT), .b(D_104_NOT), .O(ED_521) );
and2 gate( .a(CONST1), .b(D_104), .O(ED_522) );
and2 gate( .a(CONST0), .b(D_104), .O(ED_523) );
and2 gate( .a(ED_520), .b(D_105_NOT), .O(ED_529) );
and2 gate( .a(ED_521), .b(D_105), .O(ED_527) );
and2 gate( .a(ED_522), .b(D_105_NOT), .O(ED_525) );
and2 gate( .a(ED_523), .b(D_105), .O(ED_524) );
or2  gate( .a(ED_524), .b(ED_525), .O(ED_526) );
or2  gate( .a(ED_526), .b(ED_527), .O(ED_528) );
or2  gate( .a(ED_529), .b(ED_528), .O(N332_OBF) );
inv1 gate( .a(D_106), .O(D_106_NOT) );
inv1 gate( .a(D_107), .O(D_107_NOT) );
inv1 gate( .a(N230), .O(N230_NOT) );
and2 gate( .a(N230), .b(D_106_NOT), .O(ED_530) );
and2 gate( .a(N230_NOT), .b(D_106_NOT), .O(ED_531) );
and2 gate( .a(CONST1), .b(D_106), .O(ED_532) );
and2 gate( .a(CONST0), .b(D_106), .O(ED_533) );
and2 gate( .a(ED_530), .b(D_107_NOT), .O(ED_539) );
and2 gate( .a(ED_531), .b(D_107), .O(ED_537) );
and2 gate( .a(ED_532), .b(D_107_NOT), .O(ED_535) );
and2 gate( .a(ED_533), .b(D_107), .O(ED_534) );
or2  gate( .a(ED_534), .b(ED_535), .O(ED_536) );
or2  gate( .a(ED_536), .b(ED_537), .O(ED_538) );
or2  gate( .a(ED_539), .b(ED_538), .O(N230_OBF) );
inv1 gate( .a(D_108), .O(D_108_NOT) );
inv1 gate( .a(D_109), .O(D_109_NOT) );
inv1 gate( .a(N230), .O(N230_NOT) );
and2 gate( .a(N230), .b(D_108_NOT), .O(ED_540) );
and2 gate( .a(N230_NOT), .b(D_108_NOT), .O(ED_541) );
and2 gate( .a(CONST1), .b(D_108), .O(ED_542) );
and2 gate( .a(CONST0), .b(D_108), .O(ED_543) );
and2 gate( .a(ED_540), .b(D_109_NOT), .O(ED_549) );
and2 gate( .a(ED_541), .b(D_109), .O(ED_547) );
and2 gate( .a(ED_542), .b(D_109_NOT), .O(ED_545) );
and2 gate( .a(ED_543), .b(D_109), .O(ED_544) );
or2  gate( .a(ED_544), .b(ED_545), .O(ED_546) );
or2  gate( .a(ED_546), .b(ED_547), .O(ED_548) );
or2  gate( .a(ED_549), .b(ED_548), .O(N230_OBF) );
inv1 gate( .a(D_110), .O(D_110_NOT) );
inv1 gate( .a(D_111), .O(D_111_NOT) );
inv1 gate( .a(N63), .O(N63_NOT) );
and2 gate( .a(N63), .b(D_110_NOT), .O(ED_550) );
and2 gate( .a(N63_NOT), .b(D_110_NOT), .O(ED_551) );
and2 gate( .a(CONST1), .b(D_110), .O(ED_552) );
and2 gate( .a(CONST0), .b(D_110), .O(ED_553) );
and2 gate( .a(ED_550), .b(D_111_NOT), .O(ED_559) );
and2 gate( .a(ED_551), .b(D_111), .O(ED_557) );
and2 gate( .a(ED_552), .b(D_111_NOT), .O(ED_555) );
and2 gate( .a(ED_553), .b(D_111), .O(ED_554) );
or2  gate( .a(ED_554), .b(ED_555), .O(ED_556) );
or2  gate( .a(ED_556), .b(ED_557), .O(ED_558) );
or2  gate( .a(ED_559), .b(ED_558), .O(N63_OBF) );

endmodule
