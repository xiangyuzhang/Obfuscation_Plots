module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );

  xor2  gate469(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate470(.a(gate20inter0), .b(s_44), .O(gate20inter1));
  and2  gate471(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate472(.a(s_44), .O(gate20inter3));
  inv1  gate473(.a(s_45), .O(gate20inter4));
  nand2 gate474(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate475(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate476(.a(N8), .O(gate20inter7));
  inv1  gate477(.a(N119), .O(gate20inter8));
  nand2 gate478(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate479(.a(s_45), .b(gate20inter3), .O(gate20inter10));
  nor2  gate480(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate481(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate482(.a(gate20inter12), .b(gate20inter1), .O(N157));

  xor2  gate623(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate624(.a(gate21inter0), .b(s_66), .O(gate21inter1));
  and2  gate625(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate626(.a(s_66), .O(gate21inter3));
  inv1  gate627(.a(s_67), .O(gate21inter4));
  nand2 gate628(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate629(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate630(.a(N14), .O(gate21inter7));
  inv1  gate631(.a(N119), .O(gate21inter8));
  nand2 gate632(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate633(.a(s_67), .b(gate21inter3), .O(gate21inter10));
  nor2  gate634(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate635(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate636(.a(gate21inter12), .b(gate21inter1), .O(N158));
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );

  xor2  gate399(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate400(.a(gate31inter0), .b(s_34), .O(gate31inter1));
  and2  gate401(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate402(.a(s_34), .O(gate31inter3));
  inv1  gate403(.a(s_35), .O(gate31inter4));
  nand2 gate404(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate405(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate406(.a(N27), .O(gate31inter7));
  inv1  gate407(.a(N123), .O(gate31inter8));
  nand2 gate408(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate409(.a(s_35), .b(gate31inter3), .O(gate31inter10));
  nor2  gate410(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate411(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate412(.a(gate31inter12), .b(gate31inter1), .O(N184));

  xor2  gate427(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate428(.a(gate32inter0), .b(s_38), .O(gate32inter1));
  and2  gate429(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate430(.a(s_38), .O(gate32inter3));
  inv1  gate431(.a(s_39), .O(gate32inter4));
  nand2 gate432(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate433(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate434(.a(N34), .O(gate32inter7));
  inv1  gate435(.a(N127), .O(gate32inter8));
  nand2 gate436(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate437(.a(s_39), .b(gate32inter3), .O(gate32inter10));
  nor2  gate438(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate439(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate440(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate161(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate162(.a(gate34inter0), .b(s_0), .O(gate34inter1));
  and2  gate163(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate164(.a(s_0), .O(gate34inter3));
  inv1  gate165(.a(s_1), .O(gate34inter4));
  nand2 gate166(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate167(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate168(.a(N47), .O(gate34inter7));
  inv1  gate169(.a(N131), .O(gate34inter8));
  nand2 gate170(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate171(.a(s_1), .b(gate34inter3), .O(gate34inter10));
  nor2  gate172(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate173(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate174(.a(gate34inter12), .b(gate34inter1), .O(N187));
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate525(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate526(.a(gate36inter0), .b(s_52), .O(gate36inter1));
  and2  gate527(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate528(.a(s_52), .O(gate36inter3));
  inv1  gate529(.a(s_53), .O(gate36inter4));
  nand2 gate530(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate531(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate532(.a(N60), .O(gate36inter7));
  inv1  gate533(.a(N135), .O(gate36inter8));
  nand2 gate534(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate535(.a(s_53), .b(gate36inter3), .O(gate36inter10));
  nor2  gate536(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate537(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate538(.a(gate36inter12), .b(gate36inter1), .O(N189));

  xor2  gate287(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate288(.a(gate37inter0), .b(s_18), .O(gate37inter1));
  and2  gate289(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate290(.a(s_18), .O(gate37inter3));
  inv1  gate291(.a(s_19), .O(gate37inter4));
  nand2 gate292(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate293(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate294(.a(N66), .O(gate37inter7));
  inv1  gate295(.a(N135), .O(gate37inter8));
  nand2 gate296(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate297(.a(s_19), .b(gate37inter3), .O(gate37inter10));
  nor2  gate298(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate299(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate300(.a(gate37inter12), .b(gate37inter1), .O(N190));
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate301(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate302(.a(gate41inter0), .b(s_20), .O(gate41inter1));
  and2  gate303(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate304(.a(s_20), .O(gate41inter3));
  inv1  gate305(.a(s_21), .O(gate41inter4));
  nand2 gate306(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate307(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate308(.a(N92), .O(gate41inter7));
  inv1  gate309(.a(N143), .O(gate41inter8));
  nand2 gate310(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate311(.a(s_21), .b(gate41inter3), .O(gate41inter10));
  nor2  gate312(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate313(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate314(.a(gate41inter12), .b(gate41inter1), .O(N194));

  xor2  gate511(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate512(.a(gate42inter0), .b(s_50), .O(gate42inter1));
  and2  gate513(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate514(.a(s_50), .O(gate42inter3));
  inv1  gate515(.a(s_51), .O(gate42inter4));
  nand2 gate516(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate517(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate518(.a(N99), .O(gate42inter7));
  inv1  gate519(.a(N147), .O(gate42inter8));
  nand2 gate520(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate521(.a(s_51), .b(gate42inter3), .O(gate42inter10));
  nor2  gate522(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate523(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate524(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate245(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate246(.a(gate52inter0), .b(s_12), .O(gate52inter1));
  and2  gate247(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate248(.a(s_12), .O(gate52inter3));
  inv1  gate249(.a(s_13), .O(gate52inter4));
  nand2 gate250(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate251(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate252(.a(N203), .O(gate52inter7));
  inv1  gate253(.a(N162), .O(gate52inter8));
  nand2 gate254(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate255(.a(s_13), .b(gate52inter3), .O(gate52inter10));
  nor2  gate256(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate257(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate258(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate413(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate414(.a(gate57inter0), .b(s_36), .O(gate57inter1));
  and2  gate415(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate416(.a(s_36), .O(gate57inter3));
  inv1  gate417(.a(s_37), .O(gate57inter4));
  nand2 gate418(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate419(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate420(.a(N203), .O(gate57inter7));
  inv1  gate421(.a(N174), .O(gate57inter8));
  nand2 gate422(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate423(.a(s_37), .b(gate57inter3), .O(gate57inter10));
  nor2  gate424(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate425(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate426(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate203(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate204(.a(gate60inter0), .b(s_6), .O(gate60inter1));
  and2  gate205(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate206(.a(s_6), .O(gate60inter3));
  inv1  gate207(.a(s_7), .O(gate60inter4));
  nand2 gate208(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate209(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate210(.a(N213), .O(gate60inter7));
  inv1  gate211(.a(N24), .O(gate60inter8));
  nand2 gate212(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate213(.a(s_7), .b(gate60inter3), .O(gate60inter10));
  nor2  gate214(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate215(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate216(.a(gate60inter12), .b(gate60inter1), .O(N250));

  xor2  gate609(.a(N180), .b(N203), .O(gate61inter0));
  nand2 gate610(.a(gate61inter0), .b(s_64), .O(gate61inter1));
  and2  gate611(.a(N180), .b(N203), .O(gate61inter2));
  inv1  gate612(.a(s_64), .O(gate61inter3));
  inv1  gate613(.a(s_65), .O(gate61inter4));
  nand2 gate614(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate615(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate616(.a(N203), .O(gate61inter7));
  inv1  gate617(.a(N180), .O(gate61inter8));
  nand2 gate618(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate619(.a(s_65), .b(gate61inter3), .O(gate61inter10));
  nor2  gate620(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate621(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate622(.a(gate61inter12), .b(gate61inter1), .O(N251));
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );

  xor2  gate343(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate344(.a(gate64inter0), .b(s_26), .O(gate64inter1));
  and2  gate345(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate346(.a(s_26), .O(gate64inter3));
  inv1  gate347(.a(s_27), .O(gate64inter4));
  nand2 gate348(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate349(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate350(.a(N213), .O(gate64inter7));
  inv1  gate351(.a(N63), .O(gate64inter8));
  nand2 gate352(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate353(.a(s_27), .b(gate64inter3), .O(gate64inter10));
  nor2  gate354(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate355(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate356(.a(gate64inter12), .b(gate64inter1), .O(N256));
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate259(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate260(.a(gate75inter0), .b(s_14), .O(gate75inter1));
  and2  gate261(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate262(.a(s_14), .O(gate75inter3));
  inv1  gate263(.a(s_15), .O(gate75inter4));
  nand2 gate264(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate265(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate266(.a(N243), .O(gate75inter7));
  inv1  gate267(.a(N193), .O(gate75inter8));
  nand2 gate268(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate269(.a(s_15), .b(gate75inter3), .O(gate75inter10));
  nor2  gate270(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate271(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate272(.a(gate75inter12), .b(gate75inter1), .O(N279));

  xor2  gate217(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate218(.a(gate76inter0), .b(s_8), .O(gate76inter1));
  and2  gate219(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate220(.a(s_8), .O(gate76inter3));
  inv1  gate221(.a(s_9), .O(gate76inter4));
  nand2 gate222(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate223(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate224(.a(N247), .O(gate76inter7));
  inv1  gate225(.a(N195), .O(gate76inter8));
  nand2 gate226(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate227(.a(s_9), .b(gate76inter3), .O(gate76inter10));
  nor2  gate228(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate229(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate230(.a(gate76inter12), .b(gate76inter1), .O(N282));
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate329(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate330(.a(gate80inter0), .b(s_24), .O(gate80inter1));
  and2  gate331(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate332(.a(s_24), .O(gate80inter3));
  inv1  gate333(.a(s_25), .O(gate80inter4));
  nand2 gate334(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate335(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate336(.a(N233), .O(gate80inter7));
  inv1  gate337(.a(N188), .O(gate80inter8));
  nand2 gate338(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate339(.a(s_25), .b(gate80inter3), .O(gate80inter10));
  nor2  gate340(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate341(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate342(.a(gate80inter12), .b(gate80inter1), .O(N290));

  xor2  gate581(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate582(.a(gate81inter0), .b(s_60), .O(gate81inter1));
  and2  gate583(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate584(.a(s_60), .O(gate81inter3));
  inv1  gate585(.a(s_61), .O(gate81inter4));
  nand2 gate586(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate587(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate588(.a(N236), .O(gate81inter7));
  inv1  gate589(.a(N190), .O(gate81inter8));
  nand2 gate590(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate591(.a(s_61), .b(gate81inter3), .O(gate81inter10));
  nor2  gate592(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate593(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate594(.a(gate81inter12), .b(gate81inter1), .O(N291));

  xor2  gate637(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate638(.a(gate82inter0), .b(s_68), .O(gate82inter1));
  and2  gate639(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate640(.a(s_68), .O(gate82inter3));
  inv1  gate641(.a(s_69), .O(gate82inter4));
  nand2 gate642(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate643(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate644(.a(N239), .O(gate82inter7));
  inv1  gate645(.a(N192), .O(gate82inter8));
  nand2 gate646(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate647(.a(s_69), .b(gate82inter3), .O(gate82inter10));
  nor2  gate648(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate649(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate650(.a(gate82inter12), .b(gate82inter1), .O(N292));
nand2 gate83( .a(N243), .b(N194), .O(N293) );

  xor2  gate651(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate652(.a(gate84inter0), .b(s_70), .O(gate84inter1));
  and2  gate653(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate654(.a(s_70), .O(gate84inter3));
  inv1  gate655(.a(s_71), .O(gate84inter4));
  nand2 gate656(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate657(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate658(.a(N247), .O(gate84inter7));
  inv1  gate659(.a(N196), .O(gate84inter8));
  nand2 gate660(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate661(.a(s_71), .b(gate84inter3), .O(gate84inter10));
  nor2  gate662(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate663(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate664(.a(gate84inter12), .b(gate84inter1), .O(N294));
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate567(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate568(.a(gate99inter0), .b(s_58), .O(gate99inter1));
  and2  gate569(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate570(.a(s_58), .O(gate99inter3));
  inv1  gate571(.a(s_59), .O(gate99inter4));
  nand2 gate572(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate573(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate574(.a(N309), .O(gate99inter7));
  inv1  gate575(.a(N260), .O(gate99inter8));
  nand2 gate576(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate577(.a(s_59), .b(gate99inter3), .O(gate99inter10));
  nor2  gate578(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate579(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate580(.a(gate99inter12), .b(gate99inter1), .O(N330));

  xor2  gate273(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate274(.a(gate100inter0), .b(s_16), .O(gate100inter1));
  and2  gate275(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate276(.a(s_16), .O(gate100inter3));
  inv1  gate277(.a(s_17), .O(gate100inter4));
  nand2 gate278(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate279(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate280(.a(N309), .O(gate100inter7));
  inv1  gate281(.a(N264), .O(gate100inter8));
  nand2 gate282(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate283(.a(s_17), .b(gate100inter3), .O(gate100inter10));
  nor2  gate284(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate285(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate286(.a(gate100inter12), .b(gate100inter1), .O(N331));
xor2 gate101( .a(N309), .b(N267), .O(N332) );

  xor2  gate497(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate498(.a(gate102inter0), .b(s_48), .O(gate102inter1));
  and2  gate499(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate500(.a(s_48), .O(gate102inter3));
  inv1  gate501(.a(s_49), .O(gate102inter4));
  nand2 gate502(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate503(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate504(.a(N309), .O(gate102inter7));
  inv1  gate505(.a(N270), .O(gate102inter8));
  nand2 gate506(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate507(.a(s_49), .b(gate102inter3), .O(gate102inter10));
  nor2  gate508(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate509(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate510(.a(gate102inter12), .b(gate102inter1), .O(N333));
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate315(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate316(.a(gate105inter0), .b(s_22), .O(gate105inter1));
  and2  gate317(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate318(.a(s_22), .O(gate105inter3));
  inv1  gate319(.a(s_23), .O(gate105inter4));
  nand2 gate320(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate321(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate322(.a(N319), .O(gate105inter7));
  inv1  gate323(.a(N21), .O(gate105inter8));
  nand2 gate324(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate325(.a(s_23), .b(gate105inter3), .O(gate105inter10));
  nor2  gate326(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate327(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate328(.a(gate105inter12), .b(gate105inter1), .O(N336));

  xor2  gate539(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate540(.a(gate106inter0), .b(s_54), .O(gate106inter1));
  and2  gate541(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate542(.a(s_54), .O(gate106inter3));
  inv1  gate543(.a(s_55), .O(gate106inter4));
  nand2 gate544(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate545(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate546(.a(N309), .O(gate106inter7));
  inv1  gate547(.a(N276), .O(gate106inter8));
  nand2 gate548(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate549(.a(s_55), .b(gate106inter3), .O(gate106inter10));
  nor2  gate550(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate551(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate552(.a(gate106inter12), .b(gate106inter1), .O(N337));
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );

  xor2  gate385(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate386(.a(gate109inter0), .b(s_32), .O(gate109inter1));
  and2  gate387(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate388(.a(s_32), .O(gate109inter3));
  inv1  gate389(.a(s_33), .O(gate109inter4));
  nand2 gate390(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate391(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate392(.a(N319), .O(gate109inter7));
  inv1  gate393(.a(N47), .O(gate109inter8));
  nand2 gate394(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate395(.a(s_33), .b(gate109inter3), .O(gate109inter10));
  nor2  gate396(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate397(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate398(.a(gate109inter12), .b(gate109inter1), .O(N340));

  xor2  gate231(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate232(.a(gate110inter0), .b(s_10), .O(gate110inter1));
  and2  gate233(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate234(.a(s_10), .O(gate110inter3));
  inv1  gate235(.a(s_11), .O(gate110inter4));
  nand2 gate236(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate237(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate238(.a(N309), .O(gate110inter7));
  inv1  gate239(.a(N282), .O(gate110inter8));
  nand2 gate240(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate241(.a(s_11), .b(gate110inter3), .O(gate110inter10));
  nor2  gate242(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate243(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate244(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );

  xor2  gate553(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate554(.a(gate114inter0), .b(s_56), .O(gate114inter1));
  and2  gate555(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate556(.a(s_56), .O(gate114inter3));
  inv1  gate557(.a(s_57), .O(gate114inter4));
  nand2 gate558(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate559(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate560(.a(N319), .O(gate114inter7));
  inv1  gate561(.a(N86), .O(gate114inter8));
  nand2 gate562(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate563(.a(s_57), .b(gate114inter3), .O(gate114inter10));
  nor2  gate564(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate565(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate566(.a(gate114inter12), .b(gate114inter1), .O(N345));

  xor2  gate595(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate596(.a(gate115inter0), .b(s_62), .O(gate115inter1));
  and2  gate597(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate598(.a(s_62), .O(gate115inter3));
  inv1  gate599(.a(s_63), .O(gate115inter4));
  nand2 gate600(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate601(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate602(.a(N319), .O(gate115inter7));
  inv1  gate603(.a(N99), .O(gate115inter8));
  nand2 gate604(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate605(.a(s_63), .b(gate115inter3), .O(gate115inter10));
  nor2  gate606(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate607(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate608(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate455(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate456(.a(gate121inter0), .b(s_42), .O(gate121inter1));
  and2  gate457(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate458(.a(s_42), .O(gate121inter3));
  inv1  gate459(.a(s_43), .O(gate121inter4));
  nand2 gate460(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate461(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate462(.a(N335), .O(gate121inter7));
  inv1  gate463(.a(N304), .O(gate121inter8));
  nand2 gate464(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate465(.a(s_43), .b(gate121inter3), .O(gate121inter10));
  nor2  gate466(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate467(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate468(.a(gate121inter12), .b(gate121inter1), .O(N352));

  xor2  gate357(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate358(.a(gate122inter0), .b(s_28), .O(gate122inter1));
  and2  gate359(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate360(.a(s_28), .O(gate122inter3));
  inv1  gate361(.a(s_29), .O(gate122inter4));
  nand2 gate362(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate363(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate364(.a(N337), .O(gate122inter7));
  inv1  gate365(.a(N305), .O(gate122inter8));
  nand2 gate366(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate367(.a(s_29), .b(gate122inter3), .O(gate122inter10));
  nor2  gate368(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate369(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate370(.a(gate122inter12), .b(gate122inter1), .O(N353));

  xor2  gate189(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate190(.a(gate123inter0), .b(s_4), .O(gate123inter1));
  and2  gate191(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate192(.a(s_4), .O(gate123inter3));
  inv1  gate193(.a(s_5), .O(gate123inter4));
  nand2 gate194(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate195(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate196(.a(N339), .O(gate123inter7));
  inv1  gate197(.a(N306), .O(gate123inter8));
  nand2 gate198(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate199(.a(s_5), .b(gate123inter3), .O(gate123inter10));
  nor2  gate200(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate201(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate202(.a(gate123inter12), .b(gate123inter1), .O(N354));

  xor2  gate371(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate372(.a(gate124inter0), .b(s_30), .O(gate124inter1));
  and2  gate373(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate374(.a(s_30), .O(gate124inter3));
  inv1  gate375(.a(s_31), .O(gate124inter4));
  nand2 gate376(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate377(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate378(.a(N341), .O(gate124inter7));
  inv1  gate379(.a(N307), .O(gate124inter8));
  nand2 gate380(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate381(.a(s_31), .b(gate124inter3), .O(gate124inter10));
  nor2  gate382(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate383(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate384(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate483(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate484(.a(gate129inter0), .b(s_46), .O(gate129inter1));
  and2  gate485(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate486(.a(s_46), .O(gate129inter3));
  inv1  gate487(.a(s_47), .O(gate129inter4));
  nand2 gate488(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate489(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate490(.a(N14), .O(gate129inter7));
  inv1  gate491(.a(N360), .O(gate129inter8));
  nand2 gate492(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate493(.a(s_47), .b(gate129inter3), .O(gate129inter10));
  nor2  gate494(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate495(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate496(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );

  xor2  gate175(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate176(.a(gate134inter0), .b(s_2), .O(gate134inter1));
  and2  gate177(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate178(.a(s_2), .O(gate134inter3));
  inv1  gate179(.a(s_3), .O(gate134inter4));
  nand2 gate180(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate181(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate182(.a(N360), .O(gate134inter7));
  inv1  gate183(.a(N79), .O(gate134inter8));
  nand2 gate184(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate185(.a(s_3), .b(gate134inter3), .O(gate134inter10));
  nor2  gate186(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate187(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate188(.a(gate134inter12), .b(gate134inter1), .O(N376));
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );

  xor2  gate441(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate442(.a(gate137inter0), .b(s_40), .O(gate137inter1));
  and2  gate443(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate444(.a(s_40), .O(gate137inter3));
  inv1  gate445(.a(s_41), .O(gate137inter4));
  nand2 gate446(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate447(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate448(.a(N360), .O(gate137inter7));
  inv1  gate449(.a(N115), .O(gate137inter8));
  nand2 gate450(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate451(.a(s_41), .b(gate137inter3), .O(gate137inter10));
  nor2  gate452(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate453(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate454(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule