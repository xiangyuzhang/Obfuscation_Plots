module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );

  xor2  gate287(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate288(.a(gate21inter0), .b(s_18), .O(gate21inter1));
  and2  gate289(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate290(.a(s_18), .O(gate21inter3));
  inv1  gate291(.a(s_19), .O(gate21inter4));
  nand2 gate292(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate293(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate294(.a(N14), .O(gate21inter7));
  inv1  gate295(.a(N119), .O(gate21inter8));
  nand2 gate296(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate297(.a(s_19), .b(gate21inter3), .O(gate21inter10));
  nor2  gate298(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate299(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate300(.a(gate21inter12), .b(gate21inter1), .O(N158));
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate343(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate344(.a(gate23inter0), .b(s_26), .O(gate23inter1));
  and2  gate345(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate346(.a(s_26), .O(gate23inter3));
  inv1  gate347(.a(s_27), .O(gate23inter4));
  nand2 gate348(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate349(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate350(.a(N126), .O(gate23inter7));
  inv1  gate351(.a(N30), .O(gate23inter8));
  nand2 gate352(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate353(.a(s_27), .b(gate23inter3), .O(gate23inter10));
  nor2  gate354(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate355(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate356(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate301(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate302(.a(gate38inter0), .b(s_20), .O(gate38inter1));
  and2  gate303(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate304(.a(s_20), .O(gate38inter3));
  inv1  gate305(.a(s_21), .O(gate38inter4));
  nand2 gate306(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate307(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate308(.a(N73), .O(gate38inter7));
  inv1  gate309(.a(N139), .O(gate38inter8));
  nand2 gate310(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate311(.a(s_21), .b(gate38inter3), .O(gate38inter10));
  nor2  gate312(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate313(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate314(.a(gate38inter12), .b(gate38inter1), .O(N191));

  xor2  gate231(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate232(.a(gate39inter0), .b(s_10), .O(gate39inter1));
  and2  gate233(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate234(.a(s_10), .O(gate39inter3));
  inv1  gate235(.a(s_11), .O(gate39inter4));
  nand2 gate236(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate237(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate238(.a(N79), .O(gate39inter7));
  inv1  gate239(.a(N139), .O(gate39inter8));
  nand2 gate240(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate241(.a(s_11), .b(gate39inter3), .O(gate39inter10));
  nor2  gate242(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate243(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate244(.a(gate39inter12), .b(gate39inter1), .O(N192));
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );

  xor2  gate273(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate274(.a(gate66inter0), .b(s_16), .O(gate66inter1));
  and2  gate275(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate276(.a(s_16), .O(gate66inter3));
  inv1  gate277(.a(s_17), .O(gate66inter4));
  nand2 gate278(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate279(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate280(.a(N213), .O(gate66inter7));
  inv1  gate281(.a(N89), .O(gate66inter8));
  nand2 gate282(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate283(.a(s_17), .b(gate66inter3), .O(gate66inter10));
  nor2  gate284(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate285(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate286(.a(gate66inter12), .b(gate66inter1), .O(N258));

  xor2  gate329(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate330(.a(gate67inter0), .b(s_24), .O(gate67inter1));
  and2  gate331(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate332(.a(s_24), .O(gate67inter3));
  inv1  gate333(.a(s_25), .O(gate67inter4));
  nand2 gate334(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate335(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate336(.a(N213), .O(gate67inter7));
  inv1  gate337(.a(N102), .O(gate67inter8));
  nand2 gate338(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate339(.a(s_25), .b(gate67inter3), .O(gate67inter10));
  nor2  gate340(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate341(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate342(.a(gate67inter12), .b(gate67inter1), .O(N259));
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate315(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate316(.a(gate70inter0), .b(s_22), .O(gate70inter1));
  and2  gate317(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate318(.a(s_22), .O(gate70inter3));
  inv1  gate319(.a(s_23), .O(gate70inter4));
  nand2 gate320(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate321(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate322(.a(N227), .O(gate70inter7));
  inv1  gate323(.a(N183), .O(gate70inter8));
  nand2 gate324(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate325(.a(s_23), .b(gate70inter3), .O(gate70inter10));
  nor2  gate326(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate327(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate328(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate175(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate176(.a(gate72inter0), .b(s_2), .O(gate72inter1));
  and2  gate177(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate178(.a(s_2), .O(gate72inter3));
  inv1  gate179(.a(s_3), .O(gate72inter4));
  nand2 gate180(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate181(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate182(.a(N233), .O(gate72inter7));
  inv1  gate183(.a(N187), .O(gate72inter8));
  nand2 gate184(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate185(.a(s_3), .b(gate72inter3), .O(gate72inter10));
  nor2  gate186(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate187(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate188(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );

  xor2  gate371(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate372(.a(gate74inter0), .b(s_30), .O(gate74inter1));
  and2  gate373(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate374(.a(s_30), .O(gate74inter3));
  inv1  gate375(.a(s_31), .O(gate74inter4));
  nand2 gate376(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate377(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate378(.a(N239), .O(gate74inter7));
  inv1  gate379(.a(N191), .O(gate74inter8));
  nand2 gate380(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate381(.a(s_31), .b(gate74inter3), .O(gate74inter10));
  nor2  gate382(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate383(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate384(.a(gate74inter12), .b(gate74inter1), .O(N276));
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate203(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate204(.a(gate83inter0), .b(s_6), .O(gate83inter1));
  and2  gate205(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate206(.a(s_6), .O(gate83inter3));
  inv1  gate207(.a(s_7), .O(gate83inter4));
  nand2 gate208(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate209(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate210(.a(N243), .O(gate83inter7));
  inv1  gate211(.a(N194), .O(gate83inter8));
  nand2 gate212(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate213(.a(s_7), .b(gate83inter3), .O(gate83inter10));
  nor2  gate214(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate215(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate216(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate161(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate162(.a(gate99inter0), .b(s_0), .O(gate99inter1));
  and2  gate163(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate164(.a(s_0), .O(gate99inter3));
  inv1  gate165(.a(s_1), .O(gate99inter4));
  nand2 gate166(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate167(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate168(.a(N309), .O(gate99inter7));
  inv1  gate169(.a(N260), .O(gate99inter8));
  nand2 gate170(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate171(.a(s_1), .b(gate99inter3), .O(gate99inter10));
  nor2  gate172(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate173(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate174(.a(gate99inter12), .b(gate99inter1), .O(N330));
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );

  xor2  gate245(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate246(.a(gate108inter0), .b(s_12), .O(gate108inter1));
  and2  gate247(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate248(.a(s_12), .O(gate108inter3));
  inv1  gate249(.a(s_13), .O(gate108inter4));
  nand2 gate250(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate251(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate252(.a(N309), .O(gate108inter7));
  inv1  gate253(.a(N279), .O(gate108inter8));
  nand2 gate254(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate255(.a(s_13), .b(gate108inter3), .O(gate108inter10));
  nor2  gate256(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate257(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate258(.a(gate108inter12), .b(gate108inter1), .O(N339));
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate189(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate190(.a(gate110inter0), .b(s_4), .O(gate110inter1));
  and2  gate191(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate192(.a(s_4), .O(gate110inter3));
  inv1  gate193(.a(s_5), .O(gate110inter4));
  nand2 gate194(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate195(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate196(.a(N309), .O(gate110inter7));
  inv1  gate197(.a(N282), .O(gate110inter8));
  nand2 gate198(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate199(.a(s_5), .b(gate110inter3), .O(gate110inter10));
  nor2  gate200(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate201(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate202(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate217(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate218(.a(gate115inter0), .b(s_8), .O(gate115inter1));
  and2  gate219(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate220(.a(s_8), .O(gate115inter3));
  inv1  gate221(.a(s_9), .O(gate115inter4));
  nand2 gate222(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate223(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate224(.a(N319), .O(gate115inter7));
  inv1  gate225(.a(N99), .O(gate115inter8));
  nand2 gate226(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate227(.a(s_9), .b(gate115inter3), .O(gate115inter10));
  nor2  gate228(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate229(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate230(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );

  xor2  gate357(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate358(.a(gate123inter0), .b(s_28), .O(gate123inter1));
  and2  gate359(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate360(.a(s_28), .O(gate123inter3));
  inv1  gate361(.a(s_29), .O(gate123inter4));
  nand2 gate362(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate363(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate364(.a(N339), .O(gate123inter7));
  inv1  gate365(.a(N306), .O(gate123inter8));
  nand2 gate366(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate367(.a(s_29), .b(gate123inter3), .O(gate123inter10));
  nor2  gate368(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate369(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate370(.a(gate123inter12), .b(gate123inter1), .O(N354));
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate259(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate260(.a(gate129inter0), .b(s_14), .O(gate129inter1));
  and2  gate261(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate262(.a(s_14), .O(gate129inter3));
  inv1  gate263(.a(s_15), .O(gate129inter4));
  nand2 gate264(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate265(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate266(.a(N14), .O(gate129inter7));
  inv1  gate267(.a(N360), .O(gate129inter8));
  nand2 gate268(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate269(.a(s_15), .b(gate129inter3), .O(gate129inter10));
  nor2  gate270(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate271(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate272(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule