
module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input  N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,      N99,N102,N105,N108,N112,N115,CONST1,CONST0 //RE__PI;

input D_0,D_1,D_2,D_3,D_4,D_5,D_6,D_7,D_8,D_9,D_10,D_11,D_12,D_13,D_14,D_15,D_16,D_17,D_18,D_19,D_20,D_21,D_22,D_23,D_24,D_25,D_26,D_27,D_28,D_29,D_30,D_31,D_32,D_33,D_34,D_35,D_36,D_37,D_38,D_39,D_40,D_41,D_42,D_43,D_44,D_45,D_46,D_47,D_48,D_49,D_50,D_51,D_52,D_53,D_54,D_55,D_56,D_57,D_58,D_59,D_60,D_61,D_62,D_63,D_64,D_65,D_66,D_67,D_68,D_69,D_70,D_71,D_72,D_73,D_74,D_75,D_76,D_77,D_78,D_79,D_80,D_81,D_82,D_83,D_84,D_85,D_86,D_87,D_88,D_89,D_90,D_91,D_92,D_93,D_94,D_95,D_96,D_97,D_98,D_99,D_100,D_101,D_102,D_103,D_104,D_105,D_106,D_107,D_108,D_109,D_110,D_111,D_112,D_113,D_114,D_115,D_116,D_117,D_118,D_119,D_120,D_121,D_122,D_123,D_124,D_125,D_126,D_127,D_128,D_129,D_130,D_131,D_132,D_133,D_134,D_135,D_136,D_137,D_138,D_139,D_140,D_141,D_142,D_143,D_144,D_145,D_146,D_147,D_148,D_149,D_150,D_151,D_152,D_153,D_154,D_155,D_156,D_157,D_158,D_159,D_160,D_161,D_162,D_163,D_164,D_165,D_166,D_167,D_168,D_169,D_170,D_171,D_172,D_173,D_174,D_175,D_176,D_177,D_178,D_179,D_180,D_181,D_182,D_183,D_184,D_185,D_186,D_187,D_188,D_189,D_190,D_191,D_192,D_193,D_194,D_195,D_196,D_197,D_198,D_199,D_200,D_201,D_202,D_203,D_204,D_205,D_206,D_207,D_208,D_209,D_210,D_211,D_212,D_213,D_214,D_215,D_216,D_217,D_218,D_219,D_220,D_221,D_222,D_223,D_224,D_225,D_226,D_227,D_228,D_229,D_230,D_231,D_232,D_233,D_234,D_235,D_236,D_237,D_238,D_239,D_240,D_241,D_242,D_243,D_244,D_245,D_246,D_247,D_248,D_249,D_250,D_251,D_252,D_253,D_254,D_255,D_256,D_257,D_258,D_259,D_260,D_261,D_262,D_263,D_264,D_265,D_266,D_267,D_268,D_269,D_270,D_271,D_272,D_273,D_274,D_275,D_276,D_277,D_278,D_279,D_280,D_281,D_282,D_283 //RE__ALLOW(00,01,10,11);

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429,D_0_NOT,D_1_NOT,N199_NOT,N199_OBF,ED_0,ED_1,ED_2,ED_3,ED_4,ED_5,ED_6,ED_7,ED_8,ED_9,D_2_NOT,D_3_NOT,N319_NOT,N319_OBF,ED_10,ED_11,ED_12,ED_13,ED_14,ED_15,ED_16,ED_17,ED_18,ED_19,D_4_NOT,D_5_NOT,N89_NOT,N89_OBF,ED_20,ED_21,ED_22,ED_23,ED_24,ED_25,ED_26,ED_27,ED_28,ED_29,D_6_NOT,D_7_NOT,N105_NOT,N105_OBF,ED_30,ED_31,ED_32,ED_33,ED_34,ED_35,ED_36,ED_37,ED_38,ED_39,D_8_NOT,D_9_NOT,N393_NOT,N393_OBF,ED_40,ED_41,ED_42,ED_43,ED_44,ED_45,ED_46,ED_47,ED_48,ED_49,D_10_NOT,D_11_NOT,N357_NOT,N357_OBF,ED_50,ED_51,ED_52,ED_53,ED_54,ED_55,ED_56,ED_57,ED_58,ED_59,D_12_NOT,D_13_NOT,N425_NOT,N425_OBF,ED_60,ED_61,ED_62,ED_63,ED_64,ED_65,ED_66,ED_67,ED_68,ED_69,D_14_NOT,D_15_NOT,N115_NOT,N115_OBF,ED_70,ED_71,ED_72,ED_73,ED_74,ED_75,ED_76,ED_77,ED_78,ED_79,D_16_NOT,D_17_NOT,N233_NOT,N233_OBF,ED_80,ED_81,ED_82,ED_83,ED_84,ED_85,ED_86,ED_87,ED_88,ED_89,D_18_NOT,D_19_NOT,N4_NOT,N4_OBF,ED_90,ED_91,ED_92,ED_93,ED_94,ED_95,ED_96,ED_97,ED_98,ED_99,D_20_NOT,D_21_NOT,N335_NOT,N335_OBF,ED_100,ED_101,ED_102,ED_103,ED_104,ED_105,ED_106,ED_107,ED_108,ED_109,D_22_NOT,D_23_NOT,N191_NOT,N191_OBF,ED_110,ED_111,ED_112,ED_113,ED_114,ED_115,ED_116,ED_117,ED_118,ED_119,D_24_NOT,D_25_NOT,N50_NOT,N50_OBF,ED_120,ED_121,ED_122,ED_123,ED_124,ED_125,ED_126,ED_127,ED_128,ED_129,D_26_NOT,D_27_NOT,N199_NOT,N199_OBF,ED_130,ED_131,ED_132,ED_133,ED_134,ED_135,ED_136,ED_137,ED_138,ED_139,D_28_NOT,D_29_NOT,N135_NOT,N135_OBF,ED_140,ED_141,ED_142,ED_143,ED_144,ED_145,ED_146,ED_147,ED_148,ED_149,D_30_NOT,D_31_NOT,N360_NOT,N360_OBF,ED_150,ED_151,ED_152,ED_153,ED_154,ED_155,ED_156,ED_157,ED_158,ED_159,D_32_NOT,D_33_NOT,N319_NOT,N319_OBF,ED_160,ED_161,ED_162,ED_163,ED_164,ED_165,ED_166,ED_167,ED_168,ED_169,D_34_NOT,D_35_NOT,N186_NOT,N186_OBF,ED_170,ED_171,ED_172,ED_173,ED_174,ED_175,ED_176,ED_177,ED_178,ED_179,D_36_NOT,D_37_NOT,N331_NOT,N331_OBF,ED_180,ED_181,ED_182,ED_183,ED_184,ED_185,ED_186,ED_187,ED_188,ED_189,D_38_NOT,D_39_NOT,N247_NOT,N247_OBF,ED_190,ED_191,ED_192,ED_193,ED_194,ED_195,ED_196,ED_197,ED_198,ED_199,D_40_NOT,D_41_NOT,N17_NOT,N17_OBF,ED_200,ED_201,ED_202,ED_203,ED_204,ED_205,ED_206,ED_207,ED_208,ED_209,D_42_NOT,D_43_NOT,N43_NOT,N43_OBF,ED_210,ED_211,ED_212,ED_213,ED_214,ED_215,ED_216,ED_217,ED_218,ED_219,D_44_NOT,D_45_NOT,N293_NOT,N293_OBF,ED_220,ED_221,ED_222,ED_223,ED_224,ED_225,ED_226,ED_227,ED_228,ED_229,D_46_NOT,D_47_NOT,N127_NOT,N127_OBF,ED_230,ED_231,ED_232,ED_233,ED_234,ED_235,ED_236,ED_237,ED_238,ED_239,D_48_NOT,D_49_NOT,N407_NOT,N407_OBF,ED_240,ED_241,ED_242,ED_243,ED_244,ED_245,ED_246,ED_247,ED_248,ED_249,D_50_NOT,D_51_NOT,N21_NOT,N21_OBF,ED_250,ED_251,ED_252,ED_253,ED_254,ED_255,ED_256,ED_257,ED_258,ED_259,D_52_NOT,D_53_NOT,N288_NOT,N288_OBF,ED_260,ED_261,ED_262,ED_263,ED_264,ED_265,ED_266,ED_267,ED_268,ED_269,D_54_NOT,D_55_NOT,N139_NOT,N139_OBF,ED_270,ED_271,ED_272,ED_273,ED_274,ED_275,ED_276,ED_277,ED_278,ED_279,D_56_NOT,D_57_NOT,N296_NOT,N296_OBF,ED_280,ED_281,ED_282,ED_283,ED_284,ED_285,ED_286,ED_287,ED_288,ED_289,D_58_NOT,D_59_NOT,N123_NOT,N123_OBF,ED_290,ED_291,ED_292,ED_293,ED_294,ED_295,ED_296,ED_297,ED_298,ED_299,D_60_NOT,D_61_NOT,N197_NOT,N197_OBF,ED_300,ED_301,ED_302,ED_303,ED_304,ED_305,ED_306,ED_307,ED_308,ED_309,D_62_NOT,D_63_NOT,N393_NOT,N393_OBF,ED_310,ED_311,ED_312,ED_313,ED_314,ED_315,ED_316,ED_317,ED_318,ED_319,D_64_NOT,D_65_NOT,N416_NOT,N416_OBF,ED_320,ED_321,ED_322,ED_323,ED_324,ED_325,ED_326,ED_327,ED_328,ED_329,D_66_NOT,D_67_NOT,N319_NOT,N319_OBF,ED_330,ED_331,ED_332,ED_333,ED_334,ED_335,ED_336,ED_337,ED_338,ED_339,D_68_NOT,D_69_NOT,N14_NOT,N14_OBF,ED_340,ED_341,ED_342,ED_343,ED_344,ED_345,ED_346,ED_347,ED_348,ED_349,D_70_NOT,D_71_NOT,N69_NOT,N69_OBF,ED_350,ED_351,ED_352,ED_353,ED_354,ED_355,ED_356,ED_357,ED_358,ED_359,D_72_NOT,D_73_NOT,N236_NOT,N236_OBF,ED_360,ED_361,ED_362,ED_363,ED_364,ED_365,ED_366,ED_367,ED_368,ED_369,D_74_NOT,D_75_NOT,N360_NOT,N360_OBF,ED_370,ED_371,ED_372,ED_373,ED_374,ED_375,ED_376,ED_377,ED_378,ED_379,D_76_NOT,D_77_NOT,N56_NOT,N56_OBF,ED_380,ED_381,ED_382,ED_383,ED_384,ED_385,ED_386,ED_387,ED_388,ED_389,D_78_NOT,D_79_NOT,N24_NOT,N24_OBF,ED_390,ED_391,ED_392,ED_393,ED_394,ED_395,ED_396,ED_397,ED_398,ED_399,D_80_NOT,D_81_NOT,N302_NOT,N302_OBF,ED_400,ED_401,ED_402,ED_403,ED_404,ED_405,ED_406,ED_407,ED_408,ED_409,D_82_NOT,D_83_NOT,N183_NOT,N183_OBF,ED_410,ED_411,ED_412,ED_413,ED_414,ED_415,ED_416,ED_417,ED_418,ED_419,D_84_NOT,D_85_NOT,N108_NOT,N108_OBF,ED_420,ED_421,ED_422,ED_423,ED_424,ED_425,ED_426,ED_427,ED_428,ED_429,D_86_NOT,D_87_NOT,N146_NOT,N146_OBF,ED_430,ED_431,ED_432,ED_433,ED_434,ED_435,ED_436,ED_437,ED_438,ED_439,D_88_NOT,D_89_NOT,N291_NOT,N291_OBF,ED_440,ED_441,ED_442,ED_443,ED_444,ED_445,ED_446,ED_447,ED_448,ED_449,D_90_NOT,D_91_NOT,N334_NOT,N334_OBF,ED_450,ED_451,ED_452,ED_453,ED_454,ED_455,ED_456,ED_457,ED_458,ED_459,D_92_NOT,D_93_NOT,N407_NOT,N407_OBF,ED_460,ED_461,ED_462,ED_463,ED_464,ED_465,ED_466,ED_467,ED_468,ED_469,D_94_NOT,D_95_NOT,N14_NOT,N14_OBF,ED_470,ED_471,ED_472,ED_473,ED_474,ED_475,ED_476,ED_477,ED_478,ED_479,D_96_NOT,D_97_NOT,N79_NOT,N79_OBF,ED_480,ED_481,ED_482,ED_483,ED_484,ED_485,ED_486,ED_487,ED_488,ED_489,D_98_NOT,D_99_NOT,N296_NOT,N296_OBF,ED_490,ED_491,ED_492,ED_493,ED_494,ED_495,ED_496,ED_497,ED_498,ED_499,D_100_NOT,D_101_NOT,N131_NOT,N131_OBF,ED_500,ED_501,ED_502,ED_503,ED_504,ED_505,ED_506,ED_507,ED_508,ED_509,D_102_NOT,D_103_NOT,N135_NOT,N135_OBF,ED_510,ED_511,ED_512,ED_513,ED_514,ED_515,ED_516,ED_517,ED_518,ED_519,D_104_NOT,D_105_NOT,N360_NOT,N360_OBF,ED_520,ED_521,ED_522,ED_523,ED_524,ED_525,ED_526,ED_527,ED_528,ED_529,D_106_NOT,D_107_NOT,N69_NOT,N69_OBF,ED_530,ED_531,ED_532,ED_533,ED_534,ED_535,ED_536,ED_537,ED_538,ED_539,D_108_NOT,D_109_NOT,N386_NOT,N386_OBF,ED_540,ED_541,ED_542,ED_543,ED_544,ED_545,ED_546,ED_547,ED_548,ED_549,D_110_NOT,D_111_NOT,N330_NOT,N330_OBF,ED_550,ED_551,ED_552,ED_553,ED_554,ED_555,ED_556,ED_557,ED_558,ED_559,D_112_NOT,D_113_NOT,N11_NOT,N11_OBF,ED_560,ED_561,ED_562,ED_563,ED_564,ED_565,ED_566,ED_567,ED_568,ED_569,D_114_NOT,D_115_NOT,N295_NOT,N295_OBF,ED_570,ED_571,ED_572,ED_573,ED_574,ED_575,ED_576,ED_577,ED_578,ED_579,D_116_NOT,D_117_NOT,N4_NOT,N4_OBF,ED_580,ED_581,ED_582,ED_583,ED_584,ED_585,ED_586,ED_587,ED_588,ED_589,D_118_NOT,D_119_NOT,N296_NOT,N296_OBF,ED_590,ED_591,ED_592,ED_593,ED_594,ED_595,ED_596,ED_597,ED_598,ED_599,D_120_NOT,D_121_NOT,N56_NOT,N56_OBF,ED_600,ED_601,ED_602,ED_603,ED_604,ED_605,ED_606,ED_607,ED_608,ED_609,D_122_NOT,D_123_NOT,N404_NOT,N404_OBF,ED_610,ED_611,ED_612,ED_613,ED_614,ED_615,ED_616,ED_617,ED_618,ED_619,D_124_NOT,D_125_NOT,N143_NOT,N143_OBF,ED_620,ED_621,ED_622,ED_623,ED_624,ED_625,ED_626,ED_627,ED_628,ED_629,D_126_NOT,D_127_NOT,N294_NOT,N294_OBF,ED_630,ED_631,ED_632,ED_633,ED_634,ED_635,ED_636,ED_637,ED_638,ED_639,D_128_NOT,D_129_NOT,N8_NOT,N8_OBF,ED_640,ED_641,ED_642,ED_643,ED_644,ED_645,ED_646,ED_647,ED_648,ED_649,D_130_NOT,D_131_NOT,N292_NOT,N292_OBF,ED_650,ED_651,ED_652,ED_653,ED_654,ED_655,ED_656,ED_657,ED_658,ED_659,D_132_NOT,D_133_NOT,N290_NOT,N290_OBF,ED_660,ED_661,ED_662,ED_663,ED_664,ED_665,ED_666,ED_667,ED_668,ED_669,D_134_NOT,D_135_NOT,N50_NOT,N50_OBF,ED_670,ED_671,ED_672,ED_673,ED_674,ED_675,ED_676,ED_677,ED_678,ED_679,D_136_NOT,D_137_NOT,N76_NOT,N76_OBF,ED_680,ED_681,ED_682,ED_683,ED_684,ED_685,ED_686,ED_687,ED_688,ED_689,D_138_NOT,D_139_NOT,N257_NOT,N257_OBF,ED_690,ED_691,ED_692,ED_693,ED_694,ED_695,ED_696,ED_697,ED_698,ED_699,D_140_NOT,D_141_NOT,N247_NOT,N247_OBF,ED_700,ED_701,ED_702,ED_703,ED_704,ED_705,ED_706,ED_707,ED_708,ED_709,D_142_NOT,D_143_NOT,N213_NOT,N213_OBF,ED_710,ED_711,ED_712,ED_713,ED_714,ED_715,ED_716,ED_717,ED_718,ED_719,D_144_NOT,D_145_NOT,N428_NOT,N428_OBF,ED_720,ED_721,ED_722,ED_723,ED_724,ED_725,ED_726,ED_727,ED_728,ED_729,D_146_NOT,D_147_NOT,N338_NOT,N338_OBF,ED_730,ED_731,ED_732,ED_733,ED_734,ED_735,ED_736,ED_737,ED_738,ED_739,D_148_NOT,D_149_NOT,N306_NOT,N306_OBF,ED_740,ED_741,ED_742,ED_743,ED_744,ED_745,ED_746,ED_747,ED_748,ED_749,D_150_NOT,D_151_NOT,N69_NOT,N69_OBF,ED_750,ED_751,ED_752,ED_753,ED_754,ED_755,ED_756,ED_757,ED_758,ED_759,D_152_NOT,D_153_NOT,N263_NOT,N263_OBF,ED_760,ED_761,ED_762,ED_763,ED_764,ED_765,ED_766,ED_767,ED_768,ED_769,D_154_NOT,D_155_NOT,N53_NOT,N53_OBF,ED_770,ED_771,ED_772,ED_773,ED_774,ED_775,ED_776,ED_777,ED_778,ED_779,D_156_NOT,D_157_NOT,N8_NOT,N8_OBF,ED_780,ED_781,ED_782,ED_783,ED_784,ED_785,ED_786,ED_787,ED_788,ED_789,D_158_NOT,D_159_NOT,N37_NOT,N37_OBF,ED_790,ED_791,ED_792,ED_793,ED_794,ED_795,ED_796,ED_797,ED_798,ED_799,D_160_NOT,D_161_NOT,N360_NOT,N360_OBF,ED_800,ED_801,ED_802,ED_803,ED_804,ED_805,ED_806,ED_807,ED_808,ED_809,D_162_NOT,D_163_NOT,N17_NOT,N17_OBF,ED_810,ED_811,ED_812,ED_813,ED_814,ED_815,ED_816,ED_817,ED_818,ED_819,D_164_NOT,D_165_NOT,N112_NOT,N112_OBF,ED_820,ED_821,ED_822,ED_823,ED_824,ED_825,ED_826,ED_827,ED_828,ED_829,D_166_NOT,D_167_NOT,N243_NOT,N243_OBF,ED_830,ED_831,ED_832,ED_833,ED_834,ED_835,ED_836,ED_837,ED_838,ED_839,D_168_NOT,D_169_NOT,N174_NOT,N174_OBF,ED_840,ED_841,ED_842,ED_843,ED_844,ED_845,ED_846,ED_847,ED_848,ED_849,D_170_NOT,D_171_NOT,N213_NOT,N213_OBF,ED_850,ED_851,ED_852,ED_853,ED_854,ED_855,ED_856,ED_857,ED_858,ED_859,D_172_NOT,D_173_NOT,N333_NOT,N333_OBF,ED_860,ED_861,ED_862,ED_863,ED_864,ED_865,ED_866,ED_867,ED_868,ED_869,D_174_NOT,D_175_NOT,N213_NOT,N213_OBF,ED_870,ED_871,ED_872,ED_873,ED_874,ED_875,ED_876,ED_877,ED_878,ED_879,D_176_NOT,D_177_NOT,N76_NOT,N76_OBF,ED_880,ED_881,ED_882,ED_883,ED_884,ED_885,ED_886,ED_887,ED_888,ED_889,D_178_NOT,D_179_NOT,N1_NOT,N1_OBF,ED_890,ED_891,ED_892,ED_893,ED_894,ED_895,ED_896,ED_897,ED_898,ED_899,D_180_NOT,D_181_NOT,N307_NOT,N307_OBF,ED_900,ED_901,ED_902,ED_903,ED_904,ED_905,ED_906,ED_907,ED_908,ED_909,D_182_NOT,D_183_NOT,N190_NOT,N190_OBF,ED_910,ED_911,ED_912,ED_913,ED_914,ED_915,ED_916,ED_917,ED_918,ED_919,D_184_NOT,D_185_NOT,N147_NOT,N147_OBF,ED_920,ED_921,ED_922,ED_923,ED_924,ED_925,ED_926,ED_927,ED_928,ED_929,D_186_NOT,D_187_NOT,N184_NOT,N184_OBF,ED_930,ED_931,ED_932,ED_933,ED_934,ED_935,ED_936,ED_937,ED_938,ED_939,D_188_NOT,D_189_NOT,N319_NOT,N319_OBF,ED_940,ED_941,ED_942,ED_943,ED_944,ED_945,ED_946,ED_947,ED_948,ED_949,D_190_NOT,D_191_NOT,N143_NOT,N143_OBF,ED_950,ED_951,ED_952,ED_953,ED_954,ED_955,ED_956,ED_957,ED_958,ED_959,D_192_NOT,D_193_NOT,N374_NOT,N374_OBF,ED_960,ED_961,ED_962,ED_963,ED_964,ED_965,ED_966,ED_967,ED_968,ED_969,D_194_NOT,D_195_NOT,N194_NOT,N194_OBF,ED_970,ED_971,ED_972,ED_973,ED_974,ED_975,ED_976,ED_977,ED_978,ED_979,D_196_NOT,D_197_NOT,N346_NOT,N346_OBF,ED_980,ED_981,ED_982,ED_983,ED_984,ED_985,ED_986,ED_987,ED_988,ED_989,D_198_NOT,D_199_NOT,N386_NOT,N386_OBF,ED_990,ED_991,ED_992,ED_993,ED_994,ED_995,ED_996,ED_997,ED_998,ED_999,D_200_NOT,D_201_NOT,N349_NOT,N349_OBF,ED_1000,ED_1001,ED_1002,ED_1003,ED_1004,ED_1005,ED_1006,ED_1007,ED_1008,ED_1009,D_202_NOT,D_203_NOT,N411_NOT,N411_OBF,ED_1010,ED_1011,ED_1012,ED_1013,ED_1014,ED_1015,ED_1016,ED_1017,ED_1018,ED_1019,D_204_NOT,D_205_NOT,N185_NOT,N185_OBF,ED_1020,ED_1021,ED_1022,ED_1023,ED_1024,ED_1025,ED_1026,ED_1027,ED_1028,ED_1029,D_206_NOT,D_207_NOT,N60_NOT,N60_OBF,ED_1030,ED_1031,ED_1032,ED_1033,ED_1034,ED_1035,ED_1036,ED_1037,ED_1038,ED_1039,D_208_NOT,D_209_NOT,N289_NOT,N289_OBF,ED_1040,ED_1041,ED_1042,ED_1043,ED_1044,ED_1045,ED_1046,ED_1047,ED_1048,ED_1049,D_210_NOT,D_211_NOT,N21_NOT,N21_OBF,ED_1050,ED_1051,ED_1052,ED_1053,ED_1054,ED_1055,ED_1056,ED_1057,ED_1058,ED_1059,D_212_NOT,D_213_NOT,N360_NOT,N360_OBF,ED_1060,ED_1061,ED_1062,ED_1063,ED_1064,ED_1065,ED_1066,ED_1067,ED_1068,ED_1069,D_214_NOT,D_215_NOT,N372_NOT,N372_OBF,ED_1070,ED_1071,ED_1072,ED_1073,ED_1074,ED_1075,ED_1076,ED_1077,ED_1078,ED_1079,D_216_NOT,D_217_NOT,N213_NOT,N213_OBF,ED_1080,ED_1081,ED_1082,ED_1083,ED_1084,ED_1085,ED_1086,ED_1087,ED_1088,ED_1089,D_218_NOT,D_219_NOT,N115_NOT,N115_OBF,ED_1090,ED_1091,ED_1092,ED_1093,ED_1094,ED_1095,ED_1096,ED_1097,ED_1098,ED_1099,D_220_NOT,D_221_NOT,N267_NOT,N267_OBF,ED_1100,ED_1101,ED_1102,ED_1103,ED_1104,ED_1105,ED_1106,ED_1107,ED_1108,ED_1109,D_222_NOT,D_223_NOT,N158_NOT,N158_OBF,ED_1110,ED_1111,ED_1112,ED_1113,ED_1114,ED_1115,ED_1116,ED_1117,ED_1118,ED_1119,D_224_NOT,D_225_NOT,N239_NOT,N239_OBF,ED_1120,ED_1121,ED_1122,ED_1123,ED_1124,ED_1125,ED_1126,ED_1127,ED_1128,ED_1129,D_226_NOT,D_227_NOT,N1_NOT,N1_OBF,ED_1130,ED_1131,ED_1132,ED_1133,ED_1134,ED_1135,ED_1136,ED_1137,ED_1138,ED_1139,D_228_NOT,D_229_NOT,N187_NOT,N187_OBF,ED_1140,ED_1141,ED_1142,ED_1143,ED_1144,ED_1145,ED_1146,ED_1147,ED_1148,ED_1149,D_230_NOT,D_231_NOT,N63_NOT,N63_OBF,ED_1150,ED_1151,ED_1152,ED_1153,ED_1154,ED_1155,ED_1156,ED_1157,ED_1158,ED_1159,D_232_NOT,D_233_NOT,N381_NOT,N381_OBF,ED_1160,ED_1161,ED_1162,ED_1163,ED_1164,ED_1165,ED_1166,ED_1167,ED_1168,ED_1169,D_234_NOT,D_235_NOT,N199_NOT,N199_OBF,ED_1170,ED_1171,ED_1172,ED_1173,ED_1174,ED_1175,ED_1176,ED_1177,ED_1178,ED_1179,D_236_NOT,D_237_NOT,N102_NOT,N102_OBF,ED_1180,ED_1181,ED_1182,ED_1183,ED_1184,ED_1185,ED_1186,ED_1187,ED_1188,ED_1189,D_238_NOT,D_239_NOT,N108_NOT,N108_OBF,ED_1190,ED_1191,ED_1192,ED_1193,ED_1194,ED_1195,ED_1196,ED_1197,ED_1198,ED_1199,D_240_NOT,D_241_NOT,N360_NOT,N360_OBF,ED_1200,ED_1201,ED_1202,ED_1203,ED_1204,ED_1205,ED_1206,ED_1207,ED_1208,ED_1209,D_242_NOT,D_243_NOT,N95_NOT,N95_OBF,ED_1210,ED_1211,ED_1212,ED_1213,ED_1214,ED_1215,ED_1216,ED_1217,ED_1218,ED_1219,D_244_NOT,D_245_NOT,N43_NOT,N43_OBF,ED_1220,ED_1221,ED_1222,ED_1223,ED_1224,ED_1225,ED_1226,ED_1227,ED_1228,ED_1229,D_246_NOT,D_247_NOT,N24_NOT,N24_OBF,ED_1230,ED_1231,ED_1232,ED_1233,ED_1234,ED_1235,ED_1236,ED_1237,ED_1238,ED_1239,D_248_NOT,D_249_NOT,N259_NOT,N259_OBF,ED_1240,ED_1241,ED_1242,ED_1243,ED_1244,ED_1245,ED_1246,ED_1247,ED_1248,ED_1249,D_250_NOT,D_251_NOT,N319_NOT,N319_OBF,ED_1250,ED_1251,ED_1252,ED_1253,ED_1254,ED_1255,ED_1256,ED_1257,ED_1258,ED_1259,D_252_NOT,D_253_NOT,N105_NOT,N105_OBF,ED_1260,ED_1261,ED_1262,ED_1263,ED_1264,ED_1265,ED_1266,ED_1267,ED_1268,ED_1269,D_254_NOT,D_255_NOT,N343_NOT,N343_OBF,ED_1270,ED_1271,ED_1272,ED_1273,ED_1274,ED_1275,ED_1276,ED_1277,ED_1278,ED_1279,D_256_NOT,D_257_NOT,N89_NOT,N89_OBF,ED_1280,ED_1281,ED_1282,ED_1283,ED_1284,ED_1285,ED_1286,ED_1287,ED_1288,ED_1289,D_258_NOT,D_259_NOT,N380_NOT,N380_OBF,ED_1290,ED_1291,ED_1292,ED_1293,ED_1294,ED_1295,ED_1296,ED_1297,ED_1298,ED_1299,D_260_NOT,D_261_NOT,N224_NOT,N224_OBF,ED_1300,ED_1301,ED_1302,ED_1303,ED_1304,ED_1305,ED_1306,ED_1307,ED_1308,ED_1309,D_262_NOT,D_263_NOT,N255_NOT,N255_OBF,ED_1310,ED_1311,ED_1312,ED_1313,ED_1314,ED_1315,ED_1316,ED_1317,ED_1318,ED_1319,D_264_NOT,D_265_NOT,N198_NOT,N198_OBF,ED_1320,ED_1321,ED_1322,ED_1323,ED_1324,ED_1325,ED_1326,ED_1327,ED_1328,ED_1329,D_266_NOT,D_267_NOT,N34_NOT,N34_OBF,ED_1330,ED_1331,ED_1332,ED_1333,ED_1334,ED_1335,ED_1336,ED_1337,ED_1338,ED_1339,D_268_NOT,D_269_NOT,N337_NOT,N337_OBF,ED_1340,ED_1341,ED_1342,ED_1343,ED_1344,ED_1345,ED_1346,ED_1347,ED_1348,ED_1349,D_270_NOT,D_271_NOT,N142_NOT,N142_OBF,ED_1350,ED_1351,ED_1352,ED_1353,ED_1354,ED_1355,ED_1356,ED_1357,ED_1358,ED_1359,D_272_NOT,D_273_NOT,N393_NOT,N393_OBF,ED_1360,ED_1361,ED_1362,ED_1363,ED_1364,ED_1365,ED_1366,ED_1367,ED_1368,ED_1369,D_274_NOT,D_275_NOT,N82_NOT,N82_OBF,ED_1370,ED_1371,ED_1372,ED_1373,ED_1374,ED_1375,ED_1376,ED_1377,ED_1378,ED_1379,D_276_NOT,D_277_NOT,N319_NOT,N319_OBF,ED_1380,ED_1381,ED_1382,ED_1383,ED_1384,ED_1385,ED_1386,ED_1387,ED_1388,ED_1389,D_278_NOT,D_279_NOT,N30_NOT,N30_OBF,ED_1390,ED_1391,ED_1392,ED_1393,ED_1394,ED_1395,ED_1396,ED_1397,ED_1398,ED_1399,D_280_NOT,D_281_NOT,N357_NOT,N357_OBF,ED_1400,ED_1401,ED_1402,ED_1403,ED_1404,ED_1405,ED_1406,ED_1407,ED_1408,ED_1409,D_282_NOT,D_283_NOT,N126_NOT,N126_OBF,ED_1410,ED_1411,ED_1412,ED_1413,ED_1414,ED_1415,ED_1416,ED_1417,ED_1418,ED_1419;


inv1 gate1( .a(N1_OBF), .O(N118) );
inv1 gate2( .a(N4_OBF), .O(N119) );
inv1 gate3( .a(N11_OBF), .O(N122) );
inv1 gate4( .a(N17_OBF), .O(N123) );
inv1 gate5( .a(N24_OBF), .O(N126) );
inv1 gate6( .a(N30_OBF), .O(N127) );
inv1 gate7( .a(N37_OBF), .O(N130) );
inv1 gate8( .a(N43_OBF), .O(N131) );
inv1 gate9( .a(N50_OBF), .O(N134) );
inv1 gate10( .a(N56_OBF), .O(N135) );
inv1 gate11( .a(N63_OBF), .O(N138) );
inv1 gate12( .a(N69_OBF), .O(N139) );
inv1 gate13( .a(N76_OBF), .O(N142) );
inv1 gate14( .a(N82_OBF), .O(N143) );
inv1 gate15( .a(N89_OBF), .O(N146) );
inv1 gate16( .a(N95_OBF), .O(N147) );
inv1 gate17( .a(N102_OBF), .O(N150) );
inv1 gate18( .a(N108_OBF), .O(N151) );
nand2 gate19( .a(N118), .b(N4_OBF), .O(N154) );
nor2 gate20( .a(N8_OBF), .b(N119), .O(N157) );
nor2 gate21( .a(N14_OBF), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17_OBF), .O(N159) );
nand2 gate23( .a(N126_OBF), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43_OBF), .O(N165) );
nand2 gate25( .a(N134), .b(N56_OBF), .O(N168) );
nand2 gate26( .a(N138), .b(N69_OBF), .O(N171) );
nand2 gate27( .a(N142_OBF), .b(N82), .O(N174) );
nand2 gate28( .a(N146_OBF), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108_OBF), .O(N180) );
nor2 gate30( .a(N21_OBF), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123_OBF), .O(N184) );
nor2 gate32( .a(N34_OBF), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127_OBF), .O(N186) );
nor2 gate34( .a(N47), .b(N131_OBF), .O(N187) );
nor2 gate35( .a(N53_OBF), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135_OBF), .O(N189) );
nor2 gate37( .a(N66), .b(N135_OBF), .O(N190) );
nor2 gate38( .a(N73), .b(N139_OBF), .O(N191) );
nor2 gate39( .a(N79_OBF), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143_OBF), .O(N193) );
nor2 gate41( .a(N92), .b(N143_OBF), .O(N194) );
nor2 gate42( .a(N99), .b(N147_OBF), .O(N195) );
nor2 gate43( .a(N105_OBF), .b(N147), .O(N196) );
nor2 gate44( .a(N112_OBF), .b(N151), .O(N197) );
nor2 gate45( .a(N115_OBF), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174_OBF), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199_OBF), .O(N203) );
inv1 gate48( .a(N199_OBF), .O(N213) );
inv1 gate49( .a(N199_OBF), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1_OBF), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213_OBF), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24_OBF), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213_OBF), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50_OBF), .O(N255) );
nand2 gate64( .a(N213_OBF), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76_OBF), .O(N257) );
nand2 gate66( .a(N213), .b(N89_OBF), .O(N258) );
nand2 gate67( .a(N213_OBF), .b(N102), .O(N259) );
nand2 gate68( .a(N224_OBF), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158_OBF), .O(N263) );
nand2 gate70( .a(N227), .b(N183_OBF), .O(N264) );
nand2 gate71( .a(N230), .b(N185_OBF), .O(N267) );
nand2 gate72( .a(N233), .b(N187_OBF), .O(N270) );
nand2 gate73( .a(N236_OBF), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191_OBF), .O(N276) );
nand2 gate75( .a(N243_OBF), .b(N193), .O(N279) );
nand2 gate76( .a(N247_OBF), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197_OBF), .O(N285) );
nand2 gate78( .a(N227), .b(N184_OBF), .O(N288) );
nand2 gate79( .a(N230), .b(N186_OBF), .O(N289) );
nand2 gate80( .a(N233_OBF), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190_OBF), .O(N291) );
nand2 gate82( .a(N239_OBF), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194_OBF), .O(N293) );
nand2 gate84( .a(N247_OBF), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198_OBF), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267_OBF), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263_OBF), .O(N300) );
inv1 gate88( .a(N288_OBF), .O(N301) );
inv1 gate89( .a(N289_OBF), .O(N302) );
inv1 gate90( .a(N290_OBF), .O(N303) );
inv1 gate91( .a(N291_OBF), .O(N304) );
inv1 gate92( .a(N292_OBF), .O(N305) );
inv1 gate93( .a(N293_OBF), .O(N306) );
inv1 gate94( .a(N294_OBF), .O(N307) );
inv1 gate95( .a(N295_OBF), .O(N308) );
inv1 gate96( .a(N296_OBF), .O(N309) );
inv1 gate97( .a(N296_OBF), .O(N319) );
inv1 gate98( .a(N296_OBF), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8_OBF), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21_OBF), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319_OBF), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319_OBF), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60_OBF), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319_OBF), .b(N73), .O(N344) );
nand2 gate114( .a(N319_OBF), .b(N86), .O(N345) );
nand2 gate115( .a(N319_OBF), .b(N99), .O(N346) );
nand2 gate116( .a(N319_OBF), .b(N112), .O(N347) );
nand2 gate117( .a(N330_OBF), .b(N300), .O(N348) );
nand2 gate118( .a(N331_OBF), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302_OBF), .O(N350) );
nand2 gate120( .a(N333_OBF), .b(N303), .O(N351) );
nand2 gate121( .a(N335_OBF), .b(N304), .O(N352) );
nand2 gate122( .a(N337_OBF), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306_OBF), .O(N354) );
nand2 gate124( .a(N341), .b(N307_OBF), .O(N355) );
nand2 gate125( .a(N343_OBF), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349_OBF), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357_OBF), .O(N360) );
inv1 gate128( .a(N357_OBF), .O(N370) );
nand2 gate129( .a(N14_OBF), .b(N360), .O(N371) );
nand2 gate130( .a(N360_OBF), .b(N27), .O(N372) );
nand2 gate131( .a(N360_OBF), .b(N40), .O(N373) );
nand2 gate132( .a(N360_OBF), .b(N53), .O(N374) );
nand2 gate133( .a(N360_OBF), .b(N66), .O(N375) );
nand2 gate134( .a(N360_OBF), .b(N79), .O(N376) );
nand2 gate135( .a(N360_OBF), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105_OBF), .O(N378) );
nand2 gate137( .a(N360), .b(N115_OBF), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334_OBF), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372_OBF), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338_OBF), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374_OBF), .d(N43), .O(N393) );
nand4 gate142( .a(N255_OBF), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69_OBF), .O(N404) );
nand4 gate144( .a(N257_OBF), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346_OBF), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259_OBF), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380_OBF), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393_OBF), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393_OBF), .O(N417) );
inv1 gate150( .a(N404_OBF), .O(N418) );
inv1 gate151( .a(N407_OBF), .O(N419) );
inv1 gate152( .a(N411_OBF), .O(N420) );
nor2 gate153( .a(N415), .b(N416_OBF), .O(N421) );
nand2 gate154( .a(N386_OBF), .b(N417), .O(N422) );
nand4 gate155( .a(N386_OBF), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393_OBF), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407_OBF), .d(N420), .O(N429) );
nand4 gate158( .a(N381_OBF), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428_OBF), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425_OBF), .d(N429), .O(N432) );
inv1 gate( .a(D_0), .O(D_0_NOT) );
inv1 gate( .a(D_1), .O(D_1_NOT) );
inv1 gate( .a(N199), .O(N199_NOT) );
and2 gate( .a(N199), .b(D_0_NOT), .O(ED_0) );
and2 gate( .a(N199_NOT), .b(D_0_NOT), .O(ED_1) );
and2 gate( .a(CONST1), .b(D_0), .O(ED_2) );
and2 gate( .a(CONST0), .b(D_0), .O(ED_3) );
and2 gate( .a(ED_0), .b(D_1_NOT), .O(ED_9) );
and2 gate( .a(ED_1), .b(D_1), .O(ED_7) );
and2 gate( .a(ED_2), .b(D_1_NOT), .O(ED_5) );
and2 gate( .a(ED_3), .b(D_1), .O(ED_4) );
or2  gate( .a(ED_4), .b(ED_5), .O(ED_6) );
or2  gate( .a(ED_6), .b(ED_7), .O(ED_8) );
or2  gate( .a(ED_9), .b(ED_8), .O(N199_OBF) );
inv1 gate( .a(D_2), .O(D_2_NOT) );
inv1 gate( .a(D_3), .O(D_3_NOT) );
inv1 gate( .a(N319), .O(N319_NOT) );
and2 gate( .a(N319), .b(D_2_NOT), .O(ED_10) );
and2 gate( .a(N319_NOT), .b(D_2_NOT), .O(ED_11) );
and2 gate( .a(CONST1), .b(D_2), .O(ED_12) );
and2 gate( .a(CONST0), .b(D_2), .O(ED_13) );
and2 gate( .a(ED_10), .b(D_3_NOT), .O(ED_19) );
and2 gate( .a(ED_11), .b(D_3), .O(ED_17) );
and2 gate( .a(ED_12), .b(D_3_NOT), .O(ED_15) );
and2 gate( .a(ED_13), .b(D_3), .O(ED_14) );
or2  gate( .a(ED_14), .b(ED_15), .O(ED_16) );
or2  gate( .a(ED_16), .b(ED_17), .O(ED_18) );
or2  gate( .a(ED_19), .b(ED_18), .O(N319_OBF) );
inv1 gate( .a(D_4), .O(D_4_NOT) );
inv1 gate( .a(D_5), .O(D_5_NOT) );
inv1 gate( .a(N89), .O(N89_NOT) );
and2 gate( .a(N89), .b(D_4_NOT), .O(ED_20) );
and2 gate( .a(N89_NOT), .b(D_4_NOT), .O(ED_21) );
and2 gate( .a(CONST1), .b(D_4), .O(ED_22) );
and2 gate( .a(CONST0), .b(D_4), .O(ED_23) );
and2 gate( .a(ED_20), .b(D_5_NOT), .O(ED_29) );
and2 gate( .a(ED_21), .b(D_5), .O(ED_27) );
and2 gate( .a(ED_22), .b(D_5_NOT), .O(ED_25) );
and2 gate( .a(ED_23), .b(D_5), .O(ED_24) );
or2  gate( .a(ED_24), .b(ED_25), .O(ED_26) );
or2  gate( .a(ED_26), .b(ED_27), .O(ED_28) );
or2  gate( .a(ED_29), .b(ED_28), .O(N89_OBF) );
inv1 gate( .a(D_6), .O(D_6_NOT) );
inv1 gate( .a(D_7), .O(D_7_NOT) );
inv1 gate( .a(N105), .O(N105_NOT) );
and2 gate( .a(N105), .b(D_6_NOT), .O(ED_30) );
and2 gate( .a(N105_NOT), .b(D_6_NOT), .O(ED_31) );
and2 gate( .a(CONST1), .b(D_6), .O(ED_32) );
and2 gate( .a(CONST0), .b(D_6), .O(ED_33) );
and2 gate( .a(ED_30), .b(D_7_NOT), .O(ED_39) );
and2 gate( .a(ED_31), .b(D_7), .O(ED_37) );
and2 gate( .a(ED_32), .b(D_7_NOT), .O(ED_35) );
and2 gate( .a(ED_33), .b(D_7), .O(ED_34) );
or2  gate( .a(ED_34), .b(ED_35), .O(ED_36) );
or2  gate( .a(ED_36), .b(ED_37), .O(ED_38) );
or2  gate( .a(ED_39), .b(ED_38), .O(N105_OBF) );
inv1 gate( .a(D_8), .O(D_8_NOT) );
inv1 gate( .a(D_9), .O(D_9_NOT) );
inv1 gate( .a(N393), .O(N393_NOT) );
and2 gate( .a(N393), .b(D_8_NOT), .O(ED_40) );
and2 gate( .a(N393_NOT), .b(D_8_NOT), .O(ED_41) );
and2 gate( .a(CONST1), .b(D_8), .O(ED_42) );
and2 gate( .a(CONST0), .b(D_8), .O(ED_43) );
and2 gate( .a(ED_40), .b(D_9_NOT), .O(ED_49) );
and2 gate( .a(ED_41), .b(D_9), .O(ED_47) );
and2 gate( .a(ED_42), .b(D_9_NOT), .O(ED_45) );
and2 gate( .a(ED_43), .b(D_9), .O(ED_44) );
or2  gate( .a(ED_44), .b(ED_45), .O(ED_46) );
or2  gate( .a(ED_46), .b(ED_47), .O(ED_48) );
or2  gate( .a(ED_49), .b(ED_48), .O(N393_OBF) );
inv1 gate( .a(D_10), .O(D_10_NOT) );
inv1 gate( .a(D_11), .O(D_11_NOT) );
inv1 gate( .a(N357), .O(N357_NOT) );
and2 gate( .a(N357), .b(D_10_NOT), .O(ED_50) );
and2 gate( .a(N357_NOT), .b(D_10_NOT), .O(ED_51) );
and2 gate( .a(CONST1), .b(D_10), .O(ED_52) );
and2 gate( .a(CONST0), .b(D_10), .O(ED_53) );
and2 gate( .a(ED_50), .b(D_11_NOT), .O(ED_59) );
and2 gate( .a(ED_51), .b(D_11), .O(ED_57) );
and2 gate( .a(ED_52), .b(D_11_NOT), .O(ED_55) );
and2 gate( .a(ED_53), .b(D_11), .O(ED_54) );
or2  gate( .a(ED_54), .b(ED_55), .O(ED_56) );
or2  gate( .a(ED_56), .b(ED_57), .O(ED_58) );
or2  gate( .a(ED_59), .b(ED_58), .O(N357_OBF) );
inv1 gate( .a(D_12), .O(D_12_NOT) );
inv1 gate( .a(D_13), .O(D_13_NOT) );
inv1 gate( .a(N425), .O(N425_NOT) );
and2 gate( .a(N425), .b(D_12_NOT), .O(ED_60) );
and2 gate( .a(N425_NOT), .b(D_12_NOT), .O(ED_61) );
and2 gate( .a(CONST1), .b(D_12), .O(ED_62) );
and2 gate( .a(CONST0), .b(D_12), .O(ED_63) );
and2 gate( .a(ED_60), .b(D_13_NOT), .O(ED_69) );
and2 gate( .a(ED_61), .b(D_13), .O(ED_67) );
and2 gate( .a(ED_62), .b(D_13_NOT), .O(ED_65) );
and2 gate( .a(ED_63), .b(D_13), .O(ED_64) );
or2  gate( .a(ED_64), .b(ED_65), .O(ED_66) );
or2  gate( .a(ED_66), .b(ED_67), .O(ED_68) );
or2  gate( .a(ED_69), .b(ED_68), .O(N425_OBF) );
inv1 gate( .a(D_14), .O(D_14_NOT) );
inv1 gate( .a(D_15), .O(D_15_NOT) );
inv1 gate( .a(N115), .O(N115_NOT) );
and2 gate( .a(N115), .b(D_14_NOT), .O(ED_70) );
and2 gate( .a(N115_NOT), .b(D_14_NOT), .O(ED_71) );
and2 gate( .a(CONST1), .b(D_14), .O(ED_72) );
and2 gate( .a(CONST0), .b(D_14), .O(ED_73) );
and2 gate( .a(ED_70), .b(D_15_NOT), .O(ED_79) );
and2 gate( .a(ED_71), .b(D_15), .O(ED_77) );
and2 gate( .a(ED_72), .b(D_15_NOT), .O(ED_75) );
and2 gate( .a(ED_73), .b(D_15), .O(ED_74) );
or2  gate( .a(ED_74), .b(ED_75), .O(ED_76) );
or2  gate( .a(ED_76), .b(ED_77), .O(ED_78) );
or2  gate( .a(ED_79), .b(ED_78), .O(N115_OBF) );
inv1 gate( .a(D_16), .O(D_16_NOT) );
inv1 gate( .a(D_17), .O(D_17_NOT) );
inv1 gate( .a(N233), .O(N233_NOT) );
and2 gate( .a(N233), .b(D_16_NOT), .O(ED_80) );
and2 gate( .a(N233_NOT), .b(D_16_NOT), .O(ED_81) );
and2 gate( .a(CONST1), .b(D_16), .O(ED_82) );
and2 gate( .a(CONST0), .b(D_16), .O(ED_83) );
and2 gate( .a(ED_80), .b(D_17_NOT), .O(ED_89) );
and2 gate( .a(ED_81), .b(D_17), .O(ED_87) );
and2 gate( .a(ED_82), .b(D_17_NOT), .O(ED_85) );
and2 gate( .a(ED_83), .b(D_17), .O(ED_84) );
or2  gate( .a(ED_84), .b(ED_85), .O(ED_86) );
or2  gate( .a(ED_86), .b(ED_87), .O(ED_88) );
or2  gate( .a(ED_89), .b(ED_88), .O(N233_OBF) );
inv1 gate( .a(D_18), .O(D_18_NOT) );
inv1 gate( .a(D_19), .O(D_19_NOT) );
inv1 gate( .a(N4), .O(N4_NOT) );
and2 gate( .a(N4), .b(D_18_NOT), .O(ED_90) );
and2 gate( .a(N4_NOT), .b(D_18_NOT), .O(ED_91) );
and2 gate( .a(CONST1), .b(D_18), .O(ED_92) );
and2 gate( .a(CONST0), .b(D_18), .O(ED_93) );
and2 gate( .a(ED_90), .b(D_19_NOT), .O(ED_99) );
and2 gate( .a(ED_91), .b(D_19), .O(ED_97) );
and2 gate( .a(ED_92), .b(D_19_NOT), .O(ED_95) );
and2 gate( .a(ED_93), .b(D_19), .O(ED_94) );
or2  gate( .a(ED_94), .b(ED_95), .O(ED_96) );
or2  gate( .a(ED_96), .b(ED_97), .O(ED_98) );
or2  gate( .a(ED_99), .b(ED_98), .O(N4_OBF) );
inv1 gate( .a(D_20), .O(D_20_NOT) );
inv1 gate( .a(D_21), .O(D_21_NOT) );
inv1 gate( .a(N335), .O(N335_NOT) );
and2 gate( .a(N335), .b(D_20_NOT), .O(ED_100) );
and2 gate( .a(N335_NOT), .b(D_20_NOT), .O(ED_101) );
and2 gate( .a(CONST1), .b(D_20), .O(ED_102) );
and2 gate( .a(CONST0), .b(D_20), .O(ED_103) );
and2 gate( .a(ED_100), .b(D_21_NOT), .O(ED_109) );
and2 gate( .a(ED_101), .b(D_21), .O(ED_107) );
and2 gate( .a(ED_102), .b(D_21_NOT), .O(ED_105) );
and2 gate( .a(ED_103), .b(D_21), .O(ED_104) );
or2  gate( .a(ED_104), .b(ED_105), .O(ED_106) );
or2  gate( .a(ED_106), .b(ED_107), .O(ED_108) );
or2  gate( .a(ED_109), .b(ED_108), .O(N335_OBF) );
inv1 gate( .a(D_22), .O(D_22_NOT) );
inv1 gate( .a(D_23), .O(D_23_NOT) );
inv1 gate( .a(N191), .O(N191_NOT) );
and2 gate( .a(N191), .b(D_22_NOT), .O(ED_110) );
and2 gate( .a(N191_NOT), .b(D_22_NOT), .O(ED_111) );
and2 gate( .a(CONST1), .b(D_22), .O(ED_112) );
and2 gate( .a(CONST0), .b(D_22), .O(ED_113) );
and2 gate( .a(ED_110), .b(D_23_NOT), .O(ED_119) );
and2 gate( .a(ED_111), .b(D_23), .O(ED_117) );
and2 gate( .a(ED_112), .b(D_23_NOT), .O(ED_115) );
and2 gate( .a(ED_113), .b(D_23), .O(ED_114) );
or2  gate( .a(ED_114), .b(ED_115), .O(ED_116) );
or2  gate( .a(ED_116), .b(ED_117), .O(ED_118) );
or2  gate( .a(ED_119), .b(ED_118), .O(N191_OBF) );
inv1 gate( .a(D_24), .O(D_24_NOT) );
inv1 gate( .a(D_25), .O(D_25_NOT) );
inv1 gate( .a(N50), .O(N50_NOT) );
and2 gate( .a(N50), .b(D_24_NOT), .O(ED_120) );
and2 gate( .a(N50_NOT), .b(D_24_NOT), .O(ED_121) );
and2 gate( .a(CONST1), .b(D_24), .O(ED_122) );
and2 gate( .a(CONST0), .b(D_24), .O(ED_123) );
and2 gate( .a(ED_120), .b(D_25_NOT), .O(ED_129) );
and2 gate( .a(ED_121), .b(D_25), .O(ED_127) );
and2 gate( .a(ED_122), .b(D_25_NOT), .O(ED_125) );
and2 gate( .a(ED_123), .b(D_25), .O(ED_124) );
or2  gate( .a(ED_124), .b(ED_125), .O(ED_126) );
or2  gate( .a(ED_126), .b(ED_127), .O(ED_128) );
or2  gate( .a(ED_129), .b(ED_128), .O(N50_OBF) );
inv1 gate( .a(D_26), .O(D_26_NOT) );
inv1 gate( .a(D_27), .O(D_27_NOT) );
inv1 gate( .a(N199), .O(N199_NOT) );
and2 gate( .a(N199), .b(D_26_NOT), .O(ED_130) );
and2 gate( .a(N199_NOT), .b(D_26_NOT), .O(ED_131) );
and2 gate( .a(CONST1), .b(D_26), .O(ED_132) );
and2 gate( .a(CONST0), .b(D_26), .O(ED_133) );
and2 gate( .a(ED_130), .b(D_27_NOT), .O(ED_139) );
and2 gate( .a(ED_131), .b(D_27), .O(ED_137) );
and2 gate( .a(ED_132), .b(D_27_NOT), .O(ED_135) );
and2 gate( .a(ED_133), .b(D_27), .O(ED_134) );
or2  gate( .a(ED_134), .b(ED_135), .O(ED_136) );
or2  gate( .a(ED_136), .b(ED_137), .O(ED_138) );
or2  gate( .a(ED_139), .b(ED_138), .O(N199_OBF) );
inv1 gate( .a(D_28), .O(D_28_NOT) );
inv1 gate( .a(D_29), .O(D_29_NOT) );
inv1 gate( .a(N135), .O(N135_NOT) );
and2 gate( .a(N135), .b(D_28_NOT), .O(ED_140) );
and2 gate( .a(N135_NOT), .b(D_28_NOT), .O(ED_141) );
and2 gate( .a(CONST1), .b(D_28), .O(ED_142) );
and2 gate( .a(CONST0), .b(D_28), .O(ED_143) );
and2 gate( .a(ED_140), .b(D_29_NOT), .O(ED_149) );
and2 gate( .a(ED_141), .b(D_29), .O(ED_147) );
and2 gate( .a(ED_142), .b(D_29_NOT), .O(ED_145) );
and2 gate( .a(ED_143), .b(D_29), .O(ED_144) );
or2  gate( .a(ED_144), .b(ED_145), .O(ED_146) );
or2  gate( .a(ED_146), .b(ED_147), .O(ED_148) );
or2  gate( .a(ED_149), .b(ED_148), .O(N135_OBF) );
inv1 gate( .a(D_30), .O(D_30_NOT) );
inv1 gate( .a(D_31), .O(D_31_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_30_NOT), .O(ED_150) );
and2 gate( .a(N360_NOT), .b(D_30_NOT), .O(ED_151) );
and2 gate( .a(CONST1), .b(D_30), .O(ED_152) );
and2 gate( .a(CONST0), .b(D_30), .O(ED_153) );
and2 gate( .a(ED_150), .b(D_31_NOT), .O(ED_159) );
and2 gate( .a(ED_151), .b(D_31), .O(ED_157) );
and2 gate( .a(ED_152), .b(D_31_NOT), .O(ED_155) );
and2 gate( .a(ED_153), .b(D_31), .O(ED_154) );
or2  gate( .a(ED_154), .b(ED_155), .O(ED_156) );
or2  gate( .a(ED_156), .b(ED_157), .O(ED_158) );
or2  gate( .a(ED_159), .b(ED_158), .O(N360_OBF) );
inv1 gate( .a(D_32), .O(D_32_NOT) );
inv1 gate( .a(D_33), .O(D_33_NOT) );
inv1 gate( .a(N319), .O(N319_NOT) );
and2 gate( .a(N319), .b(D_32_NOT), .O(ED_160) );
and2 gate( .a(N319_NOT), .b(D_32_NOT), .O(ED_161) );
and2 gate( .a(CONST1), .b(D_32), .O(ED_162) );
and2 gate( .a(CONST0), .b(D_32), .O(ED_163) );
and2 gate( .a(ED_160), .b(D_33_NOT), .O(ED_169) );
and2 gate( .a(ED_161), .b(D_33), .O(ED_167) );
and2 gate( .a(ED_162), .b(D_33_NOT), .O(ED_165) );
and2 gate( .a(ED_163), .b(D_33), .O(ED_164) );
or2  gate( .a(ED_164), .b(ED_165), .O(ED_166) );
or2  gate( .a(ED_166), .b(ED_167), .O(ED_168) );
or2  gate( .a(ED_169), .b(ED_168), .O(N319_OBF) );
inv1 gate( .a(D_34), .O(D_34_NOT) );
inv1 gate( .a(D_35), .O(D_35_NOT) );
inv1 gate( .a(N186), .O(N186_NOT) );
and2 gate( .a(N186), .b(D_34_NOT), .O(ED_170) );
and2 gate( .a(N186_NOT), .b(D_34_NOT), .O(ED_171) );
and2 gate( .a(CONST1), .b(D_34), .O(ED_172) );
and2 gate( .a(CONST0), .b(D_34), .O(ED_173) );
and2 gate( .a(ED_170), .b(D_35_NOT), .O(ED_179) );
and2 gate( .a(ED_171), .b(D_35), .O(ED_177) );
and2 gate( .a(ED_172), .b(D_35_NOT), .O(ED_175) );
and2 gate( .a(ED_173), .b(D_35), .O(ED_174) );
or2  gate( .a(ED_174), .b(ED_175), .O(ED_176) );
or2  gate( .a(ED_176), .b(ED_177), .O(ED_178) );
or2  gate( .a(ED_179), .b(ED_178), .O(N186_OBF) );
inv1 gate( .a(D_36), .O(D_36_NOT) );
inv1 gate( .a(D_37), .O(D_37_NOT) );
inv1 gate( .a(N331), .O(N331_NOT) );
and2 gate( .a(N331), .b(D_36_NOT), .O(ED_180) );
and2 gate( .a(N331_NOT), .b(D_36_NOT), .O(ED_181) );
and2 gate( .a(CONST1), .b(D_36), .O(ED_182) );
and2 gate( .a(CONST0), .b(D_36), .O(ED_183) );
and2 gate( .a(ED_180), .b(D_37_NOT), .O(ED_189) );
and2 gate( .a(ED_181), .b(D_37), .O(ED_187) );
and2 gate( .a(ED_182), .b(D_37_NOT), .O(ED_185) );
and2 gate( .a(ED_183), .b(D_37), .O(ED_184) );
or2  gate( .a(ED_184), .b(ED_185), .O(ED_186) );
or2  gate( .a(ED_186), .b(ED_187), .O(ED_188) );
or2  gate( .a(ED_189), .b(ED_188), .O(N331_OBF) );
inv1 gate( .a(D_38), .O(D_38_NOT) );
inv1 gate( .a(D_39), .O(D_39_NOT) );
inv1 gate( .a(N247), .O(N247_NOT) );
and2 gate( .a(N247), .b(D_38_NOT), .O(ED_190) );
and2 gate( .a(N247_NOT), .b(D_38_NOT), .O(ED_191) );
and2 gate( .a(CONST1), .b(D_38), .O(ED_192) );
and2 gate( .a(CONST0), .b(D_38), .O(ED_193) );
and2 gate( .a(ED_190), .b(D_39_NOT), .O(ED_199) );
and2 gate( .a(ED_191), .b(D_39), .O(ED_197) );
and2 gate( .a(ED_192), .b(D_39_NOT), .O(ED_195) );
and2 gate( .a(ED_193), .b(D_39), .O(ED_194) );
or2  gate( .a(ED_194), .b(ED_195), .O(ED_196) );
or2  gate( .a(ED_196), .b(ED_197), .O(ED_198) );
or2  gate( .a(ED_199), .b(ED_198), .O(N247_OBF) );
inv1 gate( .a(D_40), .O(D_40_NOT) );
inv1 gate( .a(D_41), .O(D_41_NOT) );
inv1 gate( .a(N17), .O(N17_NOT) );
and2 gate( .a(N17), .b(D_40_NOT), .O(ED_200) );
and2 gate( .a(N17_NOT), .b(D_40_NOT), .O(ED_201) );
and2 gate( .a(CONST1), .b(D_40), .O(ED_202) );
and2 gate( .a(CONST0), .b(D_40), .O(ED_203) );
and2 gate( .a(ED_200), .b(D_41_NOT), .O(ED_209) );
and2 gate( .a(ED_201), .b(D_41), .O(ED_207) );
and2 gate( .a(ED_202), .b(D_41_NOT), .O(ED_205) );
and2 gate( .a(ED_203), .b(D_41), .O(ED_204) );
or2  gate( .a(ED_204), .b(ED_205), .O(ED_206) );
or2  gate( .a(ED_206), .b(ED_207), .O(ED_208) );
or2  gate( .a(ED_209), .b(ED_208), .O(N17_OBF) );
inv1 gate( .a(D_42), .O(D_42_NOT) );
inv1 gate( .a(D_43), .O(D_43_NOT) );
inv1 gate( .a(N43), .O(N43_NOT) );
and2 gate( .a(N43), .b(D_42_NOT), .O(ED_210) );
and2 gate( .a(N43_NOT), .b(D_42_NOT), .O(ED_211) );
and2 gate( .a(CONST1), .b(D_42), .O(ED_212) );
and2 gate( .a(CONST0), .b(D_42), .O(ED_213) );
and2 gate( .a(ED_210), .b(D_43_NOT), .O(ED_219) );
and2 gate( .a(ED_211), .b(D_43), .O(ED_217) );
and2 gate( .a(ED_212), .b(D_43_NOT), .O(ED_215) );
and2 gate( .a(ED_213), .b(D_43), .O(ED_214) );
or2  gate( .a(ED_214), .b(ED_215), .O(ED_216) );
or2  gate( .a(ED_216), .b(ED_217), .O(ED_218) );
or2  gate( .a(ED_219), .b(ED_218), .O(N43_OBF) );
inv1 gate( .a(D_44), .O(D_44_NOT) );
inv1 gate( .a(D_45), .O(D_45_NOT) );
inv1 gate( .a(N293), .O(N293_NOT) );
and2 gate( .a(N293), .b(D_44_NOT), .O(ED_220) );
and2 gate( .a(N293_NOT), .b(D_44_NOT), .O(ED_221) );
and2 gate( .a(CONST1), .b(D_44), .O(ED_222) );
and2 gate( .a(CONST0), .b(D_44), .O(ED_223) );
and2 gate( .a(ED_220), .b(D_45_NOT), .O(ED_229) );
and2 gate( .a(ED_221), .b(D_45), .O(ED_227) );
and2 gate( .a(ED_222), .b(D_45_NOT), .O(ED_225) );
and2 gate( .a(ED_223), .b(D_45), .O(ED_224) );
or2  gate( .a(ED_224), .b(ED_225), .O(ED_226) );
or2  gate( .a(ED_226), .b(ED_227), .O(ED_228) );
or2  gate( .a(ED_229), .b(ED_228), .O(N293_OBF) );
inv1 gate( .a(D_46), .O(D_46_NOT) );
inv1 gate( .a(D_47), .O(D_47_NOT) );
inv1 gate( .a(N127), .O(N127_NOT) );
and2 gate( .a(N127), .b(D_46_NOT), .O(ED_230) );
and2 gate( .a(N127_NOT), .b(D_46_NOT), .O(ED_231) );
and2 gate( .a(CONST1), .b(D_46), .O(ED_232) );
and2 gate( .a(CONST0), .b(D_46), .O(ED_233) );
and2 gate( .a(ED_230), .b(D_47_NOT), .O(ED_239) );
and2 gate( .a(ED_231), .b(D_47), .O(ED_237) );
and2 gate( .a(ED_232), .b(D_47_NOT), .O(ED_235) );
and2 gate( .a(ED_233), .b(D_47), .O(ED_234) );
or2  gate( .a(ED_234), .b(ED_235), .O(ED_236) );
or2  gate( .a(ED_236), .b(ED_237), .O(ED_238) );
or2  gate( .a(ED_239), .b(ED_238), .O(N127_OBF) );
inv1 gate( .a(D_48), .O(D_48_NOT) );
inv1 gate( .a(D_49), .O(D_49_NOT) );
inv1 gate( .a(N407), .O(N407_NOT) );
and2 gate( .a(N407), .b(D_48_NOT), .O(ED_240) );
and2 gate( .a(N407_NOT), .b(D_48_NOT), .O(ED_241) );
and2 gate( .a(CONST1), .b(D_48), .O(ED_242) );
and2 gate( .a(CONST0), .b(D_48), .O(ED_243) );
and2 gate( .a(ED_240), .b(D_49_NOT), .O(ED_249) );
and2 gate( .a(ED_241), .b(D_49), .O(ED_247) );
and2 gate( .a(ED_242), .b(D_49_NOT), .O(ED_245) );
and2 gate( .a(ED_243), .b(D_49), .O(ED_244) );
or2  gate( .a(ED_244), .b(ED_245), .O(ED_246) );
or2  gate( .a(ED_246), .b(ED_247), .O(ED_248) );
or2  gate( .a(ED_249), .b(ED_248), .O(N407_OBF) );
inv1 gate( .a(D_50), .O(D_50_NOT) );
inv1 gate( .a(D_51), .O(D_51_NOT) );
inv1 gate( .a(N21), .O(N21_NOT) );
and2 gate( .a(N21), .b(D_50_NOT), .O(ED_250) );
and2 gate( .a(N21_NOT), .b(D_50_NOT), .O(ED_251) );
and2 gate( .a(CONST1), .b(D_50), .O(ED_252) );
and2 gate( .a(CONST0), .b(D_50), .O(ED_253) );
and2 gate( .a(ED_250), .b(D_51_NOT), .O(ED_259) );
and2 gate( .a(ED_251), .b(D_51), .O(ED_257) );
and2 gate( .a(ED_252), .b(D_51_NOT), .O(ED_255) );
and2 gate( .a(ED_253), .b(D_51), .O(ED_254) );
or2  gate( .a(ED_254), .b(ED_255), .O(ED_256) );
or2  gate( .a(ED_256), .b(ED_257), .O(ED_258) );
or2  gate( .a(ED_259), .b(ED_258), .O(N21_OBF) );
inv1 gate( .a(D_52), .O(D_52_NOT) );
inv1 gate( .a(D_53), .O(D_53_NOT) );
inv1 gate( .a(N288), .O(N288_NOT) );
and2 gate( .a(N288), .b(D_52_NOT), .O(ED_260) );
and2 gate( .a(N288_NOT), .b(D_52_NOT), .O(ED_261) );
and2 gate( .a(CONST1), .b(D_52), .O(ED_262) );
and2 gate( .a(CONST0), .b(D_52), .O(ED_263) );
and2 gate( .a(ED_260), .b(D_53_NOT), .O(ED_269) );
and2 gate( .a(ED_261), .b(D_53), .O(ED_267) );
and2 gate( .a(ED_262), .b(D_53_NOT), .O(ED_265) );
and2 gate( .a(ED_263), .b(D_53), .O(ED_264) );
or2  gate( .a(ED_264), .b(ED_265), .O(ED_266) );
or2  gate( .a(ED_266), .b(ED_267), .O(ED_268) );
or2  gate( .a(ED_269), .b(ED_268), .O(N288_OBF) );
inv1 gate( .a(D_54), .O(D_54_NOT) );
inv1 gate( .a(D_55), .O(D_55_NOT) );
inv1 gate( .a(N139), .O(N139_NOT) );
and2 gate( .a(N139), .b(D_54_NOT), .O(ED_270) );
and2 gate( .a(N139_NOT), .b(D_54_NOT), .O(ED_271) );
and2 gate( .a(CONST1), .b(D_54), .O(ED_272) );
and2 gate( .a(CONST0), .b(D_54), .O(ED_273) );
and2 gate( .a(ED_270), .b(D_55_NOT), .O(ED_279) );
and2 gate( .a(ED_271), .b(D_55), .O(ED_277) );
and2 gate( .a(ED_272), .b(D_55_NOT), .O(ED_275) );
and2 gate( .a(ED_273), .b(D_55), .O(ED_274) );
or2  gate( .a(ED_274), .b(ED_275), .O(ED_276) );
or2  gate( .a(ED_276), .b(ED_277), .O(ED_278) );
or2  gate( .a(ED_279), .b(ED_278), .O(N139_OBF) );
inv1 gate( .a(D_56), .O(D_56_NOT) );
inv1 gate( .a(D_57), .O(D_57_NOT) );
inv1 gate( .a(N296), .O(N296_NOT) );
and2 gate( .a(N296), .b(D_56_NOT), .O(ED_280) );
and2 gate( .a(N296_NOT), .b(D_56_NOT), .O(ED_281) );
and2 gate( .a(CONST1), .b(D_56), .O(ED_282) );
and2 gate( .a(CONST0), .b(D_56), .O(ED_283) );
and2 gate( .a(ED_280), .b(D_57_NOT), .O(ED_289) );
and2 gate( .a(ED_281), .b(D_57), .O(ED_287) );
and2 gate( .a(ED_282), .b(D_57_NOT), .O(ED_285) );
and2 gate( .a(ED_283), .b(D_57), .O(ED_284) );
or2  gate( .a(ED_284), .b(ED_285), .O(ED_286) );
or2  gate( .a(ED_286), .b(ED_287), .O(ED_288) );
or2  gate( .a(ED_289), .b(ED_288), .O(N296_OBF) );
inv1 gate( .a(D_58), .O(D_58_NOT) );
inv1 gate( .a(D_59), .O(D_59_NOT) );
inv1 gate( .a(N123), .O(N123_NOT) );
and2 gate( .a(N123), .b(D_58_NOT), .O(ED_290) );
and2 gate( .a(N123_NOT), .b(D_58_NOT), .O(ED_291) );
and2 gate( .a(CONST1), .b(D_58), .O(ED_292) );
and2 gate( .a(CONST0), .b(D_58), .O(ED_293) );
and2 gate( .a(ED_290), .b(D_59_NOT), .O(ED_299) );
and2 gate( .a(ED_291), .b(D_59), .O(ED_297) );
and2 gate( .a(ED_292), .b(D_59_NOT), .O(ED_295) );
and2 gate( .a(ED_293), .b(D_59), .O(ED_294) );
or2  gate( .a(ED_294), .b(ED_295), .O(ED_296) );
or2  gate( .a(ED_296), .b(ED_297), .O(ED_298) );
or2  gate( .a(ED_299), .b(ED_298), .O(N123_OBF) );
inv1 gate( .a(D_60), .O(D_60_NOT) );
inv1 gate( .a(D_61), .O(D_61_NOT) );
inv1 gate( .a(N197), .O(N197_NOT) );
and2 gate( .a(N197), .b(D_60_NOT), .O(ED_300) );
and2 gate( .a(N197_NOT), .b(D_60_NOT), .O(ED_301) );
and2 gate( .a(CONST1), .b(D_60), .O(ED_302) );
and2 gate( .a(CONST0), .b(D_60), .O(ED_303) );
and2 gate( .a(ED_300), .b(D_61_NOT), .O(ED_309) );
and2 gate( .a(ED_301), .b(D_61), .O(ED_307) );
and2 gate( .a(ED_302), .b(D_61_NOT), .O(ED_305) );
and2 gate( .a(ED_303), .b(D_61), .O(ED_304) );
or2  gate( .a(ED_304), .b(ED_305), .O(ED_306) );
or2  gate( .a(ED_306), .b(ED_307), .O(ED_308) );
or2  gate( .a(ED_309), .b(ED_308), .O(N197_OBF) );
inv1 gate( .a(D_62), .O(D_62_NOT) );
inv1 gate( .a(D_63), .O(D_63_NOT) );
inv1 gate( .a(N393), .O(N393_NOT) );
and2 gate( .a(N393), .b(D_62_NOT), .O(ED_310) );
and2 gate( .a(N393_NOT), .b(D_62_NOT), .O(ED_311) );
and2 gate( .a(CONST1), .b(D_62), .O(ED_312) );
and2 gate( .a(CONST0), .b(D_62), .O(ED_313) );
and2 gate( .a(ED_310), .b(D_63_NOT), .O(ED_319) );
and2 gate( .a(ED_311), .b(D_63), .O(ED_317) );
and2 gate( .a(ED_312), .b(D_63_NOT), .O(ED_315) );
and2 gate( .a(ED_313), .b(D_63), .O(ED_314) );
or2  gate( .a(ED_314), .b(ED_315), .O(ED_316) );
or2  gate( .a(ED_316), .b(ED_317), .O(ED_318) );
or2  gate( .a(ED_319), .b(ED_318), .O(N393_OBF) );
inv1 gate( .a(D_64), .O(D_64_NOT) );
inv1 gate( .a(D_65), .O(D_65_NOT) );
inv1 gate( .a(N416), .O(N416_NOT) );
and2 gate( .a(N416), .b(D_64_NOT), .O(ED_320) );
and2 gate( .a(N416_NOT), .b(D_64_NOT), .O(ED_321) );
and2 gate( .a(CONST1), .b(D_64), .O(ED_322) );
and2 gate( .a(CONST0), .b(D_64), .O(ED_323) );
and2 gate( .a(ED_320), .b(D_65_NOT), .O(ED_329) );
and2 gate( .a(ED_321), .b(D_65), .O(ED_327) );
and2 gate( .a(ED_322), .b(D_65_NOT), .O(ED_325) );
and2 gate( .a(ED_323), .b(D_65), .O(ED_324) );
or2  gate( .a(ED_324), .b(ED_325), .O(ED_326) );
or2  gate( .a(ED_326), .b(ED_327), .O(ED_328) );
or2  gate( .a(ED_329), .b(ED_328), .O(N416_OBF) );
inv1 gate( .a(D_66), .O(D_66_NOT) );
inv1 gate( .a(D_67), .O(D_67_NOT) );
inv1 gate( .a(N319), .O(N319_NOT) );
and2 gate( .a(N319), .b(D_66_NOT), .O(ED_330) );
and2 gate( .a(N319_NOT), .b(D_66_NOT), .O(ED_331) );
and2 gate( .a(CONST1), .b(D_66), .O(ED_332) );
and2 gate( .a(CONST0), .b(D_66), .O(ED_333) );
and2 gate( .a(ED_330), .b(D_67_NOT), .O(ED_339) );
and2 gate( .a(ED_331), .b(D_67), .O(ED_337) );
and2 gate( .a(ED_332), .b(D_67_NOT), .O(ED_335) );
and2 gate( .a(ED_333), .b(D_67), .O(ED_334) );
or2  gate( .a(ED_334), .b(ED_335), .O(ED_336) );
or2  gate( .a(ED_336), .b(ED_337), .O(ED_338) );
or2  gate( .a(ED_339), .b(ED_338), .O(N319_OBF) );
inv1 gate( .a(D_68), .O(D_68_NOT) );
inv1 gate( .a(D_69), .O(D_69_NOT) );
inv1 gate( .a(N14), .O(N14_NOT) );
and2 gate( .a(N14), .b(D_68_NOT), .O(ED_340) );
and2 gate( .a(N14_NOT), .b(D_68_NOT), .O(ED_341) );
and2 gate( .a(CONST1), .b(D_68), .O(ED_342) );
and2 gate( .a(CONST0), .b(D_68), .O(ED_343) );
and2 gate( .a(ED_340), .b(D_69_NOT), .O(ED_349) );
and2 gate( .a(ED_341), .b(D_69), .O(ED_347) );
and2 gate( .a(ED_342), .b(D_69_NOT), .O(ED_345) );
and2 gate( .a(ED_343), .b(D_69), .O(ED_344) );
or2  gate( .a(ED_344), .b(ED_345), .O(ED_346) );
or2  gate( .a(ED_346), .b(ED_347), .O(ED_348) );
or2  gate( .a(ED_349), .b(ED_348), .O(N14_OBF) );
inv1 gate( .a(D_70), .O(D_70_NOT) );
inv1 gate( .a(D_71), .O(D_71_NOT) );
inv1 gate( .a(N69), .O(N69_NOT) );
and2 gate( .a(N69), .b(D_70_NOT), .O(ED_350) );
and2 gate( .a(N69_NOT), .b(D_70_NOT), .O(ED_351) );
and2 gate( .a(CONST1), .b(D_70), .O(ED_352) );
and2 gate( .a(CONST0), .b(D_70), .O(ED_353) );
and2 gate( .a(ED_350), .b(D_71_NOT), .O(ED_359) );
and2 gate( .a(ED_351), .b(D_71), .O(ED_357) );
and2 gate( .a(ED_352), .b(D_71_NOT), .O(ED_355) );
and2 gate( .a(ED_353), .b(D_71), .O(ED_354) );
or2  gate( .a(ED_354), .b(ED_355), .O(ED_356) );
or2  gate( .a(ED_356), .b(ED_357), .O(ED_358) );
or2  gate( .a(ED_359), .b(ED_358), .O(N69_OBF) );
inv1 gate( .a(D_72), .O(D_72_NOT) );
inv1 gate( .a(D_73), .O(D_73_NOT) );
inv1 gate( .a(N236), .O(N236_NOT) );
and2 gate( .a(N236), .b(D_72_NOT), .O(ED_360) );
and2 gate( .a(N236_NOT), .b(D_72_NOT), .O(ED_361) );
and2 gate( .a(CONST1), .b(D_72), .O(ED_362) );
and2 gate( .a(CONST0), .b(D_72), .O(ED_363) );
and2 gate( .a(ED_360), .b(D_73_NOT), .O(ED_369) );
and2 gate( .a(ED_361), .b(D_73), .O(ED_367) );
and2 gate( .a(ED_362), .b(D_73_NOT), .O(ED_365) );
and2 gate( .a(ED_363), .b(D_73), .O(ED_364) );
or2  gate( .a(ED_364), .b(ED_365), .O(ED_366) );
or2  gate( .a(ED_366), .b(ED_367), .O(ED_368) );
or2  gate( .a(ED_369), .b(ED_368), .O(N236_OBF) );
inv1 gate( .a(D_74), .O(D_74_NOT) );
inv1 gate( .a(D_75), .O(D_75_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_74_NOT), .O(ED_370) );
and2 gate( .a(N360_NOT), .b(D_74_NOT), .O(ED_371) );
and2 gate( .a(CONST1), .b(D_74), .O(ED_372) );
and2 gate( .a(CONST0), .b(D_74), .O(ED_373) );
and2 gate( .a(ED_370), .b(D_75_NOT), .O(ED_379) );
and2 gate( .a(ED_371), .b(D_75), .O(ED_377) );
and2 gate( .a(ED_372), .b(D_75_NOT), .O(ED_375) );
and2 gate( .a(ED_373), .b(D_75), .O(ED_374) );
or2  gate( .a(ED_374), .b(ED_375), .O(ED_376) );
or2  gate( .a(ED_376), .b(ED_377), .O(ED_378) );
or2  gate( .a(ED_379), .b(ED_378), .O(N360_OBF) );
inv1 gate( .a(D_76), .O(D_76_NOT) );
inv1 gate( .a(D_77), .O(D_77_NOT) );
inv1 gate( .a(N56), .O(N56_NOT) );
and2 gate( .a(N56), .b(D_76_NOT), .O(ED_380) );
and2 gate( .a(N56_NOT), .b(D_76_NOT), .O(ED_381) );
and2 gate( .a(CONST1), .b(D_76), .O(ED_382) );
and2 gate( .a(CONST0), .b(D_76), .O(ED_383) );
and2 gate( .a(ED_380), .b(D_77_NOT), .O(ED_389) );
and2 gate( .a(ED_381), .b(D_77), .O(ED_387) );
and2 gate( .a(ED_382), .b(D_77_NOT), .O(ED_385) );
and2 gate( .a(ED_383), .b(D_77), .O(ED_384) );
or2  gate( .a(ED_384), .b(ED_385), .O(ED_386) );
or2  gate( .a(ED_386), .b(ED_387), .O(ED_388) );
or2  gate( .a(ED_389), .b(ED_388), .O(N56_OBF) );
inv1 gate( .a(D_78), .O(D_78_NOT) );
inv1 gate( .a(D_79), .O(D_79_NOT) );
inv1 gate( .a(N24), .O(N24_NOT) );
and2 gate( .a(N24), .b(D_78_NOT), .O(ED_390) );
and2 gate( .a(N24_NOT), .b(D_78_NOT), .O(ED_391) );
and2 gate( .a(CONST1), .b(D_78), .O(ED_392) );
and2 gate( .a(CONST0), .b(D_78), .O(ED_393) );
and2 gate( .a(ED_390), .b(D_79_NOT), .O(ED_399) );
and2 gate( .a(ED_391), .b(D_79), .O(ED_397) );
and2 gate( .a(ED_392), .b(D_79_NOT), .O(ED_395) );
and2 gate( .a(ED_393), .b(D_79), .O(ED_394) );
or2  gate( .a(ED_394), .b(ED_395), .O(ED_396) );
or2  gate( .a(ED_396), .b(ED_397), .O(ED_398) );
or2  gate( .a(ED_399), .b(ED_398), .O(N24_OBF) );
inv1 gate( .a(D_80), .O(D_80_NOT) );
inv1 gate( .a(D_81), .O(D_81_NOT) );
inv1 gate( .a(N302), .O(N302_NOT) );
and2 gate( .a(N302), .b(D_80_NOT), .O(ED_400) );
and2 gate( .a(N302_NOT), .b(D_80_NOT), .O(ED_401) );
and2 gate( .a(CONST1), .b(D_80), .O(ED_402) );
and2 gate( .a(CONST0), .b(D_80), .O(ED_403) );
and2 gate( .a(ED_400), .b(D_81_NOT), .O(ED_409) );
and2 gate( .a(ED_401), .b(D_81), .O(ED_407) );
and2 gate( .a(ED_402), .b(D_81_NOT), .O(ED_405) );
and2 gate( .a(ED_403), .b(D_81), .O(ED_404) );
or2  gate( .a(ED_404), .b(ED_405), .O(ED_406) );
or2  gate( .a(ED_406), .b(ED_407), .O(ED_408) );
or2  gate( .a(ED_409), .b(ED_408), .O(N302_OBF) );
inv1 gate( .a(D_82), .O(D_82_NOT) );
inv1 gate( .a(D_83), .O(D_83_NOT) );
inv1 gate( .a(N183), .O(N183_NOT) );
and2 gate( .a(N183), .b(D_82_NOT), .O(ED_410) );
and2 gate( .a(N183_NOT), .b(D_82_NOT), .O(ED_411) );
and2 gate( .a(CONST1), .b(D_82), .O(ED_412) );
and2 gate( .a(CONST0), .b(D_82), .O(ED_413) );
and2 gate( .a(ED_410), .b(D_83_NOT), .O(ED_419) );
and2 gate( .a(ED_411), .b(D_83), .O(ED_417) );
and2 gate( .a(ED_412), .b(D_83_NOT), .O(ED_415) );
and2 gate( .a(ED_413), .b(D_83), .O(ED_414) );
or2  gate( .a(ED_414), .b(ED_415), .O(ED_416) );
or2  gate( .a(ED_416), .b(ED_417), .O(ED_418) );
or2  gate( .a(ED_419), .b(ED_418), .O(N183_OBF) );
inv1 gate( .a(D_84), .O(D_84_NOT) );
inv1 gate( .a(D_85), .O(D_85_NOT) );
inv1 gate( .a(N108), .O(N108_NOT) );
and2 gate( .a(N108), .b(D_84_NOT), .O(ED_420) );
and2 gate( .a(N108_NOT), .b(D_84_NOT), .O(ED_421) );
and2 gate( .a(CONST1), .b(D_84), .O(ED_422) );
and2 gate( .a(CONST0), .b(D_84), .O(ED_423) );
and2 gate( .a(ED_420), .b(D_85_NOT), .O(ED_429) );
and2 gate( .a(ED_421), .b(D_85), .O(ED_427) );
and2 gate( .a(ED_422), .b(D_85_NOT), .O(ED_425) );
and2 gate( .a(ED_423), .b(D_85), .O(ED_424) );
or2  gate( .a(ED_424), .b(ED_425), .O(ED_426) );
or2  gate( .a(ED_426), .b(ED_427), .O(ED_428) );
or2  gate( .a(ED_429), .b(ED_428), .O(N108_OBF) );
inv1 gate( .a(D_86), .O(D_86_NOT) );
inv1 gate( .a(D_87), .O(D_87_NOT) );
inv1 gate( .a(N146), .O(N146_NOT) );
and2 gate( .a(N146), .b(D_86_NOT), .O(ED_430) );
and2 gate( .a(N146_NOT), .b(D_86_NOT), .O(ED_431) );
and2 gate( .a(CONST1), .b(D_86), .O(ED_432) );
and2 gate( .a(CONST0), .b(D_86), .O(ED_433) );
and2 gate( .a(ED_430), .b(D_87_NOT), .O(ED_439) );
and2 gate( .a(ED_431), .b(D_87), .O(ED_437) );
and2 gate( .a(ED_432), .b(D_87_NOT), .O(ED_435) );
and2 gate( .a(ED_433), .b(D_87), .O(ED_434) );
or2  gate( .a(ED_434), .b(ED_435), .O(ED_436) );
or2  gate( .a(ED_436), .b(ED_437), .O(ED_438) );
or2  gate( .a(ED_439), .b(ED_438), .O(N146_OBF) );
inv1 gate( .a(D_88), .O(D_88_NOT) );
inv1 gate( .a(D_89), .O(D_89_NOT) );
inv1 gate( .a(N291), .O(N291_NOT) );
and2 gate( .a(N291), .b(D_88_NOT), .O(ED_440) );
and2 gate( .a(N291_NOT), .b(D_88_NOT), .O(ED_441) );
and2 gate( .a(CONST1), .b(D_88), .O(ED_442) );
and2 gate( .a(CONST0), .b(D_88), .O(ED_443) );
and2 gate( .a(ED_440), .b(D_89_NOT), .O(ED_449) );
and2 gate( .a(ED_441), .b(D_89), .O(ED_447) );
and2 gate( .a(ED_442), .b(D_89_NOT), .O(ED_445) );
and2 gate( .a(ED_443), .b(D_89), .O(ED_444) );
or2  gate( .a(ED_444), .b(ED_445), .O(ED_446) );
or2  gate( .a(ED_446), .b(ED_447), .O(ED_448) );
or2  gate( .a(ED_449), .b(ED_448), .O(N291_OBF) );
inv1 gate( .a(D_90), .O(D_90_NOT) );
inv1 gate( .a(D_91), .O(D_91_NOT) );
inv1 gate( .a(N334), .O(N334_NOT) );
and2 gate( .a(N334), .b(D_90_NOT), .O(ED_450) );
and2 gate( .a(N334_NOT), .b(D_90_NOT), .O(ED_451) );
and2 gate( .a(CONST1), .b(D_90), .O(ED_452) );
and2 gate( .a(CONST0), .b(D_90), .O(ED_453) );
and2 gate( .a(ED_450), .b(D_91_NOT), .O(ED_459) );
and2 gate( .a(ED_451), .b(D_91), .O(ED_457) );
and2 gate( .a(ED_452), .b(D_91_NOT), .O(ED_455) );
and2 gate( .a(ED_453), .b(D_91), .O(ED_454) );
or2  gate( .a(ED_454), .b(ED_455), .O(ED_456) );
or2  gate( .a(ED_456), .b(ED_457), .O(ED_458) );
or2  gate( .a(ED_459), .b(ED_458), .O(N334_OBF) );
inv1 gate( .a(D_92), .O(D_92_NOT) );
inv1 gate( .a(D_93), .O(D_93_NOT) );
inv1 gate( .a(N407), .O(N407_NOT) );
and2 gate( .a(N407), .b(D_92_NOT), .O(ED_460) );
and2 gate( .a(N407_NOT), .b(D_92_NOT), .O(ED_461) );
and2 gate( .a(CONST1), .b(D_92), .O(ED_462) );
and2 gate( .a(CONST0), .b(D_92), .O(ED_463) );
and2 gate( .a(ED_460), .b(D_93_NOT), .O(ED_469) );
and2 gate( .a(ED_461), .b(D_93), .O(ED_467) );
and2 gate( .a(ED_462), .b(D_93_NOT), .O(ED_465) );
and2 gate( .a(ED_463), .b(D_93), .O(ED_464) );
or2  gate( .a(ED_464), .b(ED_465), .O(ED_466) );
or2  gate( .a(ED_466), .b(ED_467), .O(ED_468) );
or2  gate( .a(ED_469), .b(ED_468), .O(N407_OBF) );
inv1 gate( .a(D_94), .O(D_94_NOT) );
inv1 gate( .a(D_95), .O(D_95_NOT) );
inv1 gate( .a(N14), .O(N14_NOT) );
and2 gate( .a(N14), .b(D_94_NOT), .O(ED_470) );
and2 gate( .a(N14_NOT), .b(D_94_NOT), .O(ED_471) );
and2 gate( .a(CONST1), .b(D_94), .O(ED_472) );
and2 gate( .a(CONST0), .b(D_94), .O(ED_473) );
and2 gate( .a(ED_470), .b(D_95_NOT), .O(ED_479) );
and2 gate( .a(ED_471), .b(D_95), .O(ED_477) );
and2 gate( .a(ED_472), .b(D_95_NOT), .O(ED_475) );
and2 gate( .a(ED_473), .b(D_95), .O(ED_474) );
or2  gate( .a(ED_474), .b(ED_475), .O(ED_476) );
or2  gate( .a(ED_476), .b(ED_477), .O(ED_478) );
or2  gate( .a(ED_479), .b(ED_478), .O(N14_OBF) );
inv1 gate( .a(D_96), .O(D_96_NOT) );
inv1 gate( .a(D_97), .O(D_97_NOT) );
inv1 gate( .a(N79), .O(N79_NOT) );
and2 gate( .a(N79), .b(D_96_NOT), .O(ED_480) );
and2 gate( .a(N79_NOT), .b(D_96_NOT), .O(ED_481) );
and2 gate( .a(CONST1), .b(D_96), .O(ED_482) );
and2 gate( .a(CONST0), .b(D_96), .O(ED_483) );
and2 gate( .a(ED_480), .b(D_97_NOT), .O(ED_489) );
and2 gate( .a(ED_481), .b(D_97), .O(ED_487) );
and2 gate( .a(ED_482), .b(D_97_NOT), .O(ED_485) );
and2 gate( .a(ED_483), .b(D_97), .O(ED_484) );
or2  gate( .a(ED_484), .b(ED_485), .O(ED_486) );
or2  gate( .a(ED_486), .b(ED_487), .O(ED_488) );
or2  gate( .a(ED_489), .b(ED_488), .O(N79_OBF) );
inv1 gate( .a(D_98), .O(D_98_NOT) );
inv1 gate( .a(D_99), .O(D_99_NOT) );
inv1 gate( .a(N296), .O(N296_NOT) );
and2 gate( .a(N296), .b(D_98_NOT), .O(ED_490) );
and2 gate( .a(N296_NOT), .b(D_98_NOT), .O(ED_491) );
and2 gate( .a(CONST1), .b(D_98), .O(ED_492) );
and2 gate( .a(CONST0), .b(D_98), .O(ED_493) );
and2 gate( .a(ED_490), .b(D_99_NOT), .O(ED_499) );
and2 gate( .a(ED_491), .b(D_99), .O(ED_497) );
and2 gate( .a(ED_492), .b(D_99_NOT), .O(ED_495) );
and2 gate( .a(ED_493), .b(D_99), .O(ED_494) );
or2  gate( .a(ED_494), .b(ED_495), .O(ED_496) );
or2  gate( .a(ED_496), .b(ED_497), .O(ED_498) );
or2  gate( .a(ED_499), .b(ED_498), .O(N296_OBF) );
inv1 gate( .a(D_100), .O(D_100_NOT) );
inv1 gate( .a(D_101), .O(D_101_NOT) );
inv1 gate( .a(N131), .O(N131_NOT) );
and2 gate( .a(N131), .b(D_100_NOT), .O(ED_500) );
and2 gate( .a(N131_NOT), .b(D_100_NOT), .O(ED_501) );
and2 gate( .a(CONST1), .b(D_100), .O(ED_502) );
and2 gate( .a(CONST0), .b(D_100), .O(ED_503) );
and2 gate( .a(ED_500), .b(D_101_NOT), .O(ED_509) );
and2 gate( .a(ED_501), .b(D_101), .O(ED_507) );
and2 gate( .a(ED_502), .b(D_101_NOT), .O(ED_505) );
and2 gate( .a(ED_503), .b(D_101), .O(ED_504) );
or2  gate( .a(ED_504), .b(ED_505), .O(ED_506) );
or2  gate( .a(ED_506), .b(ED_507), .O(ED_508) );
or2  gate( .a(ED_509), .b(ED_508), .O(N131_OBF) );
inv1 gate( .a(D_102), .O(D_102_NOT) );
inv1 gate( .a(D_103), .O(D_103_NOT) );
inv1 gate( .a(N135), .O(N135_NOT) );
and2 gate( .a(N135), .b(D_102_NOT), .O(ED_510) );
and2 gate( .a(N135_NOT), .b(D_102_NOT), .O(ED_511) );
and2 gate( .a(CONST1), .b(D_102), .O(ED_512) );
and2 gate( .a(CONST0), .b(D_102), .O(ED_513) );
and2 gate( .a(ED_510), .b(D_103_NOT), .O(ED_519) );
and2 gate( .a(ED_511), .b(D_103), .O(ED_517) );
and2 gate( .a(ED_512), .b(D_103_NOT), .O(ED_515) );
and2 gate( .a(ED_513), .b(D_103), .O(ED_514) );
or2  gate( .a(ED_514), .b(ED_515), .O(ED_516) );
or2  gate( .a(ED_516), .b(ED_517), .O(ED_518) );
or2  gate( .a(ED_519), .b(ED_518), .O(N135_OBF) );
inv1 gate( .a(D_104), .O(D_104_NOT) );
inv1 gate( .a(D_105), .O(D_105_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_104_NOT), .O(ED_520) );
and2 gate( .a(N360_NOT), .b(D_104_NOT), .O(ED_521) );
and2 gate( .a(CONST1), .b(D_104), .O(ED_522) );
and2 gate( .a(CONST0), .b(D_104), .O(ED_523) );
and2 gate( .a(ED_520), .b(D_105_NOT), .O(ED_529) );
and2 gate( .a(ED_521), .b(D_105), .O(ED_527) );
and2 gate( .a(ED_522), .b(D_105_NOT), .O(ED_525) );
and2 gate( .a(ED_523), .b(D_105), .O(ED_524) );
or2  gate( .a(ED_524), .b(ED_525), .O(ED_526) );
or2  gate( .a(ED_526), .b(ED_527), .O(ED_528) );
or2  gate( .a(ED_529), .b(ED_528), .O(N360_OBF) );
inv1 gate( .a(D_106), .O(D_106_NOT) );
inv1 gate( .a(D_107), .O(D_107_NOT) );
inv1 gate( .a(N69), .O(N69_NOT) );
and2 gate( .a(N69), .b(D_106_NOT), .O(ED_530) );
and2 gate( .a(N69_NOT), .b(D_106_NOT), .O(ED_531) );
and2 gate( .a(CONST1), .b(D_106), .O(ED_532) );
and2 gate( .a(CONST0), .b(D_106), .O(ED_533) );
and2 gate( .a(ED_530), .b(D_107_NOT), .O(ED_539) );
and2 gate( .a(ED_531), .b(D_107), .O(ED_537) );
and2 gate( .a(ED_532), .b(D_107_NOT), .O(ED_535) );
and2 gate( .a(ED_533), .b(D_107), .O(ED_534) );
or2  gate( .a(ED_534), .b(ED_535), .O(ED_536) );
or2  gate( .a(ED_536), .b(ED_537), .O(ED_538) );
or2  gate( .a(ED_539), .b(ED_538), .O(N69_OBF) );
inv1 gate( .a(D_108), .O(D_108_NOT) );
inv1 gate( .a(D_109), .O(D_109_NOT) );
inv1 gate( .a(N386), .O(N386_NOT) );
and2 gate( .a(N386), .b(D_108_NOT), .O(ED_540) );
and2 gate( .a(N386_NOT), .b(D_108_NOT), .O(ED_541) );
and2 gate( .a(CONST1), .b(D_108), .O(ED_542) );
and2 gate( .a(CONST0), .b(D_108), .O(ED_543) );
and2 gate( .a(ED_540), .b(D_109_NOT), .O(ED_549) );
and2 gate( .a(ED_541), .b(D_109), .O(ED_547) );
and2 gate( .a(ED_542), .b(D_109_NOT), .O(ED_545) );
and2 gate( .a(ED_543), .b(D_109), .O(ED_544) );
or2  gate( .a(ED_544), .b(ED_545), .O(ED_546) );
or2  gate( .a(ED_546), .b(ED_547), .O(ED_548) );
or2  gate( .a(ED_549), .b(ED_548), .O(N386_OBF) );
inv1 gate( .a(D_110), .O(D_110_NOT) );
inv1 gate( .a(D_111), .O(D_111_NOT) );
inv1 gate( .a(N330), .O(N330_NOT) );
and2 gate( .a(N330), .b(D_110_NOT), .O(ED_550) );
and2 gate( .a(N330_NOT), .b(D_110_NOT), .O(ED_551) );
and2 gate( .a(CONST1), .b(D_110), .O(ED_552) );
and2 gate( .a(CONST0), .b(D_110), .O(ED_553) );
and2 gate( .a(ED_550), .b(D_111_NOT), .O(ED_559) );
and2 gate( .a(ED_551), .b(D_111), .O(ED_557) );
and2 gate( .a(ED_552), .b(D_111_NOT), .O(ED_555) );
and2 gate( .a(ED_553), .b(D_111), .O(ED_554) );
or2  gate( .a(ED_554), .b(ED_555), .O(ED_556) );
or2  gate( .a(ED_556), .b(ED_557), .O(ED_558) );
or2  gate( .a(ED_559), .b(ED_558), .O(N330_OBF) );
inv1 gate( .a(D_112), .O(D_112_NOT) );
inv1 gate( .a(D_113), .O(D_113_NOT) );
inv1 gate( .a(N11), .O(N11_NOT) );
and2 gate( .a(N11), .b(D_112_NOT), .O(ED_560) );
and2 gate( .a(N11_NOT), .b(D_112_NOT), .O(ED_561) );
and2 gate( .a(CONST1), .b(D_112), .O(ED_562) );
and2 gate( .a(CONST0), .b(D_112), .O(ED_563) );
and2 gate( .a(ED_560), .b(D_113_NOT), .O(ED_569) );
and2 gate( .a(ED_561), .b(D_113), .O(ED_567) );
and2 gate( .a(ED_562), .b(D_113_NOT), .O(ED_565) );
and2 gate( .a(ED_563), .b(D_113), .O(ED_564) );
or2  gate( .a(ED_564), .b(ED_565), .O(ED_566) );
or2  gate( .a(ED_566), .b(ED_567), .O(ED_568) );
or2  gate( .a(ED_569), .b(ED_568), .O(N11_OBF) );
inv1 gate( .a(D_114), .O(D_114_NOT) );
inv1 gate( .a(D_115), .O(D_115_NOT) );
inv1 gate( .a(N295), .O(N295_NOT) );
and2 gate( .a(N295), .b(D_114_NOT), .O(ED_570) );
and2 gate( .a(N295_NOT), .b(D_114_NOT), .O(ED_571) );
and2 gate( .a(CONST1), .b(D_114), .O(ED_572) );
and2 gate( .a(CONST0), .b(D_114), .O(ED_573) );
and2 gate( .a(ED_570), .b(D_115_NOT), .O(ED_579) );
and2 gate( .a(ED_571), .b(D_115), .O(ED_577) );
and2 gate( .a(ED_572), .b(D_115_NOT), .O(ED_575) );
and2 gate( .a(ED_573), .b(D_115), .O(ED_574) );
or2  gate( .a(ED_574), .b(ED_575), .O(ED_576) );
or2  gate( .a(ED_576), .b(ED_577), .O(ED_578) );
or2  gate( .a(ED_579), .b(ED_578), .O(N295_OBF) );
inv1 gate( .a(D_116), .O(D_116_NOT) );
inv1 gate( .a(D_117), .O(D_117_NOT) );
inv1 gate( .a(N4), .O(N4_NOT) );
and2 gate( .a(N4), .b(D_116_NOT), .O(ED_580) );
and2 gate( .a(N4_NOT), .b(D_116_NOT), .O(ED_581) );
and2 gate( .a(CONST1), .b(D_116), .O(ED_582) );
and2 gate( .a(CONST0), .b(D_116), .O(ED_583) );
and2 gate( .a(ED_580), .b(D_117_NOT), .O(ED_589) );
and2 gate( .a(ED_581), .b(D_117), .O(ED_587) );
and2 gate( .a(ED_582), .b(D_117_NOT), .O(ED_585) );
and2 gate( .a(ED_583), .b(D_117), .O(ED_584) );
or2  gate( .a(ED_584), .b(ED_585), .O(ED_586) );
or2  gate( .a(ED_586), .b(ED_587), .O(ED_588) );
or2  gate( .a(ED_589), .b(ED_588), .O(N4_OBF) );
inv1 gate( .a(D_118), .O(D_118_NOT) );
inv1 gate( .a(D_119), .O(D_119_NOT) );
inv1 gate( .a(N296), .O(N296_NOT) );
and2 gate( .a(N296), .b(D_118_NOT), .O(ED_590) );
and2 gate( .a(N296_NOT), .b(D_118_NOT), .O(ED_591) );
and2 gate( .a(CONST1), .b(D_118), .O(ED_592) );
and2 gate( .a(CONST0), .b(D_118), .O(ED_593) );
and2 gate( .a(ED_590), .b(D_119_NOT), .O(ED_599) );
and2 gate( .a(ED_591), .b(D_119), .O(ED_597) );
and2 gate( .a(ED_592), .b(D_119_NOT), .O(ED_595) );
and2 gate( .a(ED_593), .b(D_119), .O(ED_594) );
or2  gate( .a(ED_594), .b(ED_595), .O(ED_596) );
or2  gate( .a(ED_596), .b(ED_597), .O(ED_598) );
or2  gate( .a(ED_599), .b(ED_598), .O(N296_OBF) );
inv1 gate( .a(D_120), .O(D_120_NOT) );
inv1 gate( .a(D_121), .O(D_121_NOT) );
inv1 gate( .a(N56), .O(N56_NOT) );
and2 gate( .a(N56), .b(D_120_NOT), .O(ED_600) );
and2 gate( .a(N56_NOT), .b(D_120_NOT), .O(ED_601) );
and2 gate( .a(CONST1), .b(D_120), .O(ED_602) );
and2 gate( .a(CONST0), .b(D_120), .O(ED_603) );
and2 gate( .a(ED_600), .b(D_121_NOT), .O(ED_609) );
and2 gate( .a(ED_601), .b(D_121), .O(ED_607) );
and2 gate( .a(ED_602), .b(D_121_NOT), .O(ED_605) );
and2 gate( .a(ED_603), .b(D_121), .O(ED_604) );
or2  gate( .a(ED_604), .b(ED_605), .O(ED_606) );
or2  gate( .a(ED_606), .b(ED_607), .O(ED_608) );
or2  gate( .a(ED_609), .b(ED_608), .O(N56_OBF) );
inv1 gate( .a(D_122), .O(D_122_NOT) );
inv1 gate( .a(D_123), .O(D_123_NOT) );
inv1 gate( .a(N404), .O(N404_NOT) );
and2 gate( .a(N404), .b(D_122_NOT), .O(ED_610) );
and2 gate( .a(N404_NOT), .b(D_122_NOT), .O(ED_611) );
and2 gate( .a(CONST1), .b(D_122), .O(ED_612) );
and2 gate( .a(CONST0), .b(D_122), .O(ED_613) );
and2 gate( .a(ED_610), .b(D_123_NOT), .O(ED_619) );
and2 gate( .a(ED_611), .b(D_123), .O(ED_617) );
and2 gate( .a(ED_612), .b(D_123_NOT), .O(ED_615) );
and2 gate( .a(ED_613), .b(D_123), .O(ED_614) );
or2  gate( .a(ED_614), .b(ED_615), .O(ED_616) );
or2  gate( .a(ED_616), .b(ED_617), .O(ED_618) );
or2  gate( .a(ED_619), .b(ED_618), .O(N404_OBF) );
inv1 gate( .a(D_124), .O(D_124_NOT) );
inv1 gate( .a(D_125), .O(D_125_NOT) );
inv1 gate( .a(N143), .O(N143_NOT) );
and2 gate( .a(N143), .b(D_124_NOT), .O(ED_620) );
and2 gate( .a(N143_NOT), .b(D_124_NOT), .O(ED_621) );
and2 gate( .a(CONST1), .b(D_124), .O(ED_622) );
and2 gate( .a(CONST0), .b(D_124), .O(ED_623) );
and2 gate( .a(ED_620), .b(D_125_NOT), .O(ED_629) );
and2 gate( .a(ED_621), .b(D_125), .O(ED_627) );
and2 gate( .a(ED_622), .b(D_125_NOT), .O(ED_625) );
and2 gate( .a(ED_623), .b(D_125), .O(ED_624) );
or2  gate( .a(ED_624), .b(ED_625), .O(ED_626) );
or2  gate( .a(ED_626), .b(ED_627), .O(ED_628) );
or2  gate( .a(ED_629), .b(ED_628), .O(N143_OBF) );
inv1 gate( .a(D_126), .O(D_126_NOT) );
inv1 gate( .a(D_127), .O(D_127_NOT) );
inv1 gate( .a(N294), .O(N294_NOT) );
and2 gate( .a(N294), .b(D_126_NOT), .O(ED_630) );
and2 gate( .a(N294_NOT), .b(D_126_NOT), .O(ED_631) );
and2 gate( .a(CONST1), .b(D_126), .O(ED_632) );
and2 gate( .a(CONST0), .b(D_126), .O(ED_633) );
and2 gate( .a(ED_630), .b(D_127_NOT), .O(ED_639) );
and2 gate( .a(ED_631), .b(D_127), .O(ED_637) );
and2 gate( .a(ED_632), .b(D_127_NOT), .O(ED_635) );
and2 gate( .a(ED_633), .b(D_127), .O(ED_634) );
or2  gate( .a(ED_634), .b(ED_635), .O(ED_636) );
or2  gate( .a(ED_636), .b(ED_637), .O(ED_638) );
or2  gate( .a(ED_639), .b(ED_638), .O(N294_OBF) );
inv1 gate( .a(D_128), .O(D_128_NOT) );
inv1 gate( .a(D_129), .O(D_129_NOT) );
inv1 gate( .a(N8), .O(N8_NOT) );
and2 gate( .a(N8), .b(D_128_NOT), .O(ED_640) );
and2 gate( .a(N8_NOT), .b(D_128_NOT), .O(ED_641) );
and2 gate( .a(CONST1), .b(D_128), .O(ED_642) );
and2 gate( .a(CONST0), .b(D_128), .O(ED_643) );
and2 gate( .a(ED_640), .b(D_129_NOT), .O(ED_649) );
and2 gate( .a(ED_641), .b(D_129), .O(ED_647) );
and2 gate( .a(ED_642), .b(D_129_NOT), .O(ED_645) );
and2 gate( .a(ED_643), .b(D_129), .O(ED_644) );
or2  gate( .a(ED_644), .b(ED_645), .O(ED_646) );
or2  gate( .a(ED_646), .b(ED_647), .O(ED_648) );
or2  gate( .a(ED_649), .b(ED_648), .O(N8_OBF) );
inv1 gate( .a(D_130), .O(D_130_NOT) );
inv1 gate( .a(D_131), .O(D_131_NOT) );
inv1 gate( .a(N292), .O(N292_NOT) );
and2 gate( .a(N292), .b(D_130_NOT), .O(ED_650) );
and2 gate( .a(N292_NOT), .b(D_130_NOT), .O(ED_651) );
and2 gate( .a(CONST1), .b(D_130), .O(ED_652) );
and2 gate( .a(CONST0), .b(D_130), .O(ED_653) );
and2 gate( .a(ED_650), .b(D_131_NOT), .O(ED_659) );
and2 gate( .a(ED_651), .b(D_131), .O(ED_657) );
and2 gate( .a(ED_652), .b(D_131_NOT), .O(ED_655) );
and2 gate( .a(ED_653), .b(D_131), .O(ED_654) );
or2  gate( .a(ED_654), .b(ED_655), .O(ED_656) );
or2  gate( .a(ED_656), .b(ED_657), .O(ED_658) );
or2  gate( .a(ED_659), .b(ED_658), .O(N292_OBF) );
inv1 gate( .a(D_132), .O(D_132_NOT) );
inv1 gate( .a(D_133), .O(D_133_NOT) );
inv1 gate( .a(N290), .O(N290_NOT) );
and2 gate( .a(N290), .b(D_132_NOT), .O(ED_660) );
and2 gate( .a(N290_NOT), .b(D_132_NOT), .O(ED_661) );
and2 gate( .a(CONST1), .b(D_132), .O(ED_662) );
and2 gate( .a(CONST0), .b(D_132), .O(ED_663) );
and2 gate( .a(ED_660), .b(D_133_NOT), .O(ED_669) );
and2 gate( .a(ED_661), .b(D_133), .O(ED_667) );
and2 gate( .a(ED_662), .b(D_133_NOT), .O(ED_665) );
and2 gate( .a(ED_663), .b(D_133), .O(ED_664) );
or2  gate( .a(ED_664), .b(ED_665), .O(ED_666) );
or2  gate( .a(ED_666), .b(ED_667), .O(ED_668) );
or2  gate( .a(ED_669), .b(ED_668), .O(N290_OBF) );
inv1 gate( .a(D_134), .O(D_134_NOT) );
inv1 gate( .a(D_135), .O(D_135_NOT) );
inv1 gate( .a(N50), .O(N50_NOT) );
and2 gate( .a(N50), .b(D_134_NOT), .O(ED_670) );
and2 gate( .a(N50_NOT), .b(D_134_NOT), .O(ED_671) );
and2 gate( .a(CONST1), .b(D_134), .O(ED_672) );
and2 gate( .a(CONST0), .b(D_134), .O(ED_673) );
and2 gate( .a(ED_670), .b(D_135_NOT), .O(ED_679) );
and2 gate( .a(ED_671), .b(D_135), .O(ED_677) );
and2 gate( .a(ED_672), .b(D_135_NOT), .O(ED_675) );
and2 gate( .a(ED_673), .b(D_135), .O(ED_674) );
or2  gate( .a(ED_674), .b(ED_675), .O(ED_676) );
or2  gate( .a(ED_676), .b(ED_677), .O(ED_678) );
or2  gate( .a(ED_679), .b(ED_678), .O(N50_OBF) );
inv1 gate( .a(D_136), .O(D_136_NOT) );
inv1 gate( .a(D_137), .O(D_137_NOT) );
inv1 gate( .a(N76), .O(N76_NOT) );
and2 gate( .a(N76), .b(D_136_NOT), .O(ED_680) );
and2 gate( .a(N76_NOT), .b(D_136_NOT), .O(ED_681) );
and2 gate( .a(CONST1), .b(D_136), .O(ED_682) );
and2 gate( .a(CONST0), .b(D_136), .O(ED_683) );
and2 gate( .a(ED_680), .b(D_137_NOT), .O(ED_689) );
and2 gate( .a(ED_681), .b(D_137), .O(ED_687) );
and2 gate( .a(ED_682), .b(D_137_NOT), .O(ED_685) );
and2 gate( .a(ED_683), .b(D_137), .O(ED_684) );
or2  gate( .a(ED_684), .b(ED_685), .O(ED_686) );
or2  gate( .a(ED_686), .b(ED_687), .O(ED_688) );
or2  gate( .a(ED_689), .b(ED_688), .O(N76_OBF) );
inv1 gate( .a(D_138), .O(D_138_NOT) );
inv1 gate( .a(D_139), .O(D_139_NOT) );
inv1 gate( .a(N257), .O(N257_NOT) );
and2 gate( .a(N257), .b(D_138_NOT), .O(ED_690) );
and2 gate( .a(N257_NOT), .b(D_138_NOT), .O(ED_691) );
and2 gate( .a(CONST1), .b(D_138), .O(ED_692) );
and2 gate( .a(CONST0), .b(D_138), .O(ED_693) );
and2 gate( .a(ED_690), .b(D_139_NOT), .O(ED_699) );
and2 gate( .a(ED_691), .b(D_139), .O(ED_697) );
and2 gate( .a(ED_692), .b(D_139_NOT), .O(ED_695) );
and2 gate( .a(ED_693), .b(D_139), .O(ED_694) );
or2  gate( .a(ED_694), .b(ED_695), .O(ED_696) );
or2  gate( .a(ED_696), .b(ED_697), .O(ED_698) );
or2  gate( .a(ED_699), .b(ED_698), .O(N257_OBF) );
inv1 gate( .a(D_140), .O(D_140_NOT) );
inv1 gate( .a(D_141), .O(D_141_NOT) );
inv1 gate( .a(N247), .O(N247_NOT) );
and2 gate( .a(N247), .b(D_140_NOT), .O(ED_700) );
and2 gate( .a(N247_NOT), .b(D_140_NOT), .O(ED_701) );
and2 gate( .a(CONST1), .b(D_140), .O(ED_702) );
and2 gate( .a(CONST0), .b(D_140), .O(ED_703) );
and2 gate( .a(ED_700), .b(D_141_NOT), .O(ED_709) );
and2 gate( .a(ED_701), .b(D_141), .O(ED_707) );
and2 gate( .a(ED_702), .b(D_141_NOT), .O(ED_705) );
and2 gate( .a(ED_703), .b(D_141), .O(ED_704) );
or2  gate( .a(ED_704), .b(ED_705), .O(ED_706) );
or2  gate( .a(ED_706), .b(ED_707), .O(ED_708) );
or2  gate( .a(ED_709), .b(ED_708), .O(N247_OBF) );
inv1 gate( .a(D_142), .O(D_142_NOT) );
inv1 gate( .a(D_143), .O(D_143_NOT) );
inv1 gate( .a(N213), .O(N213_NOT) );
and2 gate( .a(N213), .b(D_142_NOT), .O(ED_710) );
and2 gate( .a(N213_NOT), .b(D_142_NOT), .O(ED_711) );
and2 gate( .a(CONST1), .b(D_142), .O(ED_712) );
and2 gate( .a(CONST0), .b(D_142), .O(ED_713) );
and2 gate( .a(ED_710), .b(D_143_NOT), .O(ED_719) );
and2 gate( .a(ED_711), .b(D_143), .O(ED_717) );
and2 gate( .a(ED_712), .b(D_143_NOT), .O(ED_715) );
and2 gate( .a(ED_713), .b(D_143), .O(ED_714) );
or2  gate( .a(ED_714), .b(ED_715), .O(ED_716) );
or2  gate( .a(ED_716), .b(ED_717), .O(ED_718) );
or2  gate( .a(ED_719), .b(ED_718), .O(N213_OBF) );
inv1 gate( .a(D_144), .O(D_144_NOT) );
inv1 gate( .a(D_145), .O(D_145_NOT) );
inv1 gate( .a(N428), .O(N428_NOT) );
and2 gate( .a(N428), .b(D_144_NOT), .O(ED_720) );
and2 gate( .a(N428_NOT), .b(D_144_NOT), .O(ED_721) );
and2 gate( .a(CONST1), .b(D_144), .O(ED_722) );
and2 gate( .a(CONST0), .b(D_144), .O(ED_723) );
and2 gate( .a(ED_720), .b(D_145_NOT), .O(ED_729) );
and2 gate( .a(ED_721), .b(D_145), .O(ED_727) );
and2 gate( .a(ED_722), .b(D_145_NOT), .O(ED_725) );
and2 gate( .a(ED_723), .b(D_145), .O(ED_724) );
or2  gate( .a(ED_724), .b(ED_725), .O(ED_726) );
or2  gate( .a(ED_726), .b(ED_727), .O(ED_728) );
or2  gate( .a(ED_729), .b(ED_728), .O(N428_OBF) );
inv1 gate( .a(D_146), .O(D_146_NOT) );
inv1 gate( .a(D_147), .O(D_147_NOT) );
inv1 gate( .a(N338), .O(N338_NOT) );
and2 gate( .a(N338), .b(D_146_NOT), .O(ED_730) );
and2 gate( .a(N338_NOT), .b(D_146_NOT), .O(ED_731) );
and2 gate( .a(CONST1), .b(D_146), .O(ED_732) );
and2 gate( .a(CONST0), .b(D_146), .O(ED_733) );
and2 gate( .a(ED_730), .b(D_147_NOT), .O(ED_739) );
and2 gate( .a(ED_731), .b(D_147), .O(ED_737) );
and2 gate( .a(ED_732), .b(D_147_NOT), .O(ED_735) );
and2 gate( .a(ED_733), .b(D_147), .O(ED_734) );
or2  gate( .a(ED_734), .b(ED_735), .O(ED_736) );
or2  gate( .a(ED_736), .b(ED_737), .O(ED_738) );
or2  gate( .a(ED_739), .b(ED_738), .O(N338_OBF) );
inv1 gate( .a(D_148), .O(D_148_NOT) );
inv1 gate( .a(D_149), .O(D_149_NOT) );
inv1 gate( .a(N306), .O(N306_NOT) );
and2 gate( .a(N306), .b(D_148_NOT), .O(ED_740) );
and2 gate( .a(N306_NOT), .b(D_148_NOT), .O(ED_741) );
and2 gate( .a(CONST1), .b(D_148), .O(ED_742) );
and2 gate( .a(CONST0), .b(D_148), .O(ED_743) );
and2 gate( .a(ED_740), .b(D_149_NOT), .O(ED_749) );
and2 gate( .a(ED_741), .b(D_149), .O(ED_747) );
and2 gate( .a(ED_742), .b(D_149_NOT), .O(ED_745) );
and2 gate( .a(ED_743), .b(D_149), .O(ED_744) );
or2  gate( .a(ED_744), .b(ED_745), .O(ED_746) );
or2  gate( .a(ED_746), .b(ED_747), .O(ED_748) );
or2  gate( .a(ED_749), .b(ED_748), .O(N306_OBF) );
inv1 gate( .a(D_150), .O(D_150_NOT) );
inv1 gate( .a(D_151), .O(D_151_NOT) );
inv1 gate( .a(N69), .O(N69_NOT) );
and2 gate( .a(N69), .b(D_150_NOT), .O(ED_750) );
and2 gate( .a(N69_NOT), .b(D_150_NOT), .O(ED_751) );
and2 gate( .a(CONST1), .b(D_150), .O(ED_752) );
and2 gate( .a(CONST0), .b(D_150), .O(ED_753) );
and2 gate( .a(ED_750), .b(D_151_NOT), .O(ED_759) );
and2 gate( .a(ED_751), .b(D_151), .O(ED_757) );
and2 gate( .a(ED_752), .b(D_151_NOT), .O(ED_755) );
and2 gate( .a(ED_753), .b(D_151), .O(ED_754) );
or2  gate( .a(ED_754), .b(ED_755), .O(ED_756) );
or2  gate( .a(ED_756), .b(ED_757), .O(ED_758) );
or2  gate( .a(ED_759), .b(ED_758), .O(N69_OBF) );
inv1 gate( .a(D_152), .O(D_152_NOT) );
inv1 gate( .a(D_153), .O(D_153_NOT) );
inv1 gate( .a(N263), .O(N263_NOT) );
and2 gate( .a(N263), .b(D_152_NOT), .O(ED_760) );
and2 gate( .a(N263_NOT), .b(D_152_NOT), .O(ED_761) );
and2 gate( .a(CONST1), .b(D_152), .O(ED_762) );
and2 gate( .a(CONST0), .b(D_152), .O(ED_763) );
and2 gate( .a(ED_760), .b(D_153_NOT), .O(ED_769) );
and2 gate( .a(ED_761), .b(D_153), .O(ED_767) );
and2 gate( .a(ED_762), .b(D_153_NOT), .O(ED_765) );
and2 gate( .a(ED_763), .b(D_153), .O(ED_764) );
or2  gate( .a(ED_764), .b(ED_765), .O(ED_766) );
or2  gate( .a(ED_766), .b(ED_767), .O(ED_768) );
or2  gate( .a(ED_769), .b(ED_768), .O(N263_OBF) );
inv1 gate( .a(D_154), .O(D_154_NOT) );
inv1 gate( .a(D_155), .O(D_155_NOT) );
inv1 gate( .a(N53), .O(N53_NOT) );
and2 gate( .a(N53), .b(D_154_NOT), .O(ED_770) );
and2 gate( .a(N53_NOT), .b(D_154_NOT), .O(ED_771) );
and2 gate( .a(CONST1), .b(D_154), .O(ED_772) );
and2 gate( .a(CONST0), .b(D_154), .O(ED_773) );
and2 gate( .a(ED_770), .b(D_155_NOT), .O(ED_779) );
and2 gate( .a(ED_771), .b(D_155), .O(ED_777) );
and2 gate( .a(ED_772), .b(D_155_NOT), .O(ED_775) );
and2 gate( .a(ED_773), .b(D_155), .O(ED_774) );
or2  gate( .a(ED_774), .b(ED_775), .O(ED_776) );
or2  gate( .a(ED_776), .b(ED_777), .O(ED_778) );
or2  gate( .a(ED_779), .b(ED_778), .O(N53_OBF) );
inv1 gate( .a(D_156), .O(D_156_NOT) );
inv1 gate( .a(D_157), .O(D_157_NOT) );
inv1 gate( .a(N8), .O(N8_NOT) );
and2 gate( .a(N8), .b(D_156_NOT), .O(ED_780) );
and2 gate( .a(N8_NOT), .b(D_156_NOT), .O(ED_781) );
and2 gate( .a(CONST1), .b(D_156), .O(ED_782) );
and2 gate( .a(CONST0), .b(D_156), .O(ED_783) );
and2 gate( .a(ED_780), .b(D_157_NOT), .O(ED_789) );
and2 gate( .a(ED_781), .b(D_157), .O(ED_787) );
and2 gate( .a(ED_782), .b(D_157_NOT), .O(ED_785) );
and2 gate( .a(ED_783), .b(D_157), .O(ED_784) );
or2  gate( .a(ED_784), .b(ED_785), .O(ED_786) );
or2  gate( .a(ED_786), .b(ED_787), .O(ED_788) );
or2  gate( .a(ED_789), .b(ED_788), .O(N8_OBF) );
inv1 gate( .a(D_158), .O(D_158_NOT) );
inv1 gate( .a(D_159), .O(D_159_NOT) );
inv1 gate( .a(N37), .O(N37_NOT) );
and2 gate( .a(N37), .b(D_158_NOT), .O(ED_790) );
and2 gate( .a(N37_NOT), .b(D_158_NOT), .O(ED_791) );
and2 gate( .a(CONST1), .b(D_158), .O(ED_792) );
and2 gate( .a(CONST0), .b(D_158), .O(ED_793) );
and2 gate( .a(ED_790), .b(D_159_NOT), .O(ED_799) );
and2 gate( .a(ED_791), .b(D_159), .O(ED_797) );
and2 gate( .a(ED_792), .b(D_159_NOT), .O(ED_795) );
and2 gate( .a(ED_793), .b(D_159), .O(ED_794) );
or2  gate( .a(ED_794), .b(ED_795), .O(ED_796) );
or2  gate( .a(ED_796), .b(ED_797), .O(ED_798) );
or2  gate( .a(ED_799), .b(ED_798), .O(N37_OBF) );
inv1 gate( .a(D_160), .O(D_160_NOT) );
inv1 gate( .a(D_161), .O(D_161_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_160_NOT), .O(ED_800) );
and2 gate( .a(N360_NOT), .b(D_160_NOT), .O(ED_801) );
and2 gate( .a(CONST1), .b(D_160), .O(ED_802) );
and2 gate( .a(CONST0), .b(D_160), .O(ED_803) );
and2 gate( .a(ED_800), .b(D_161_NOT), .O(ED_809) );
and2 gate( .a(ED_801), .b(D_161), .O(ED_807) );
and2 gate( .a(ED_802), .b(D_161_NOT), .O(ED_805) );
and2 gate( .a(ED_803), .b(D_161), .O(ED_804) );
or2  gate( .a(ED_804), .b(ED_805), .O(ED_806) );
or2  gate( .a(ED_806), .b(ED_807), .O(ED_808) );
or2  gate( .a(ED_809), .b(ED_808), .O(N360_OBF) );
inv1 gate( .a(D_162), .O(D_162_NOT) );
inv1 gate( .a(D_163), .O(D_163_NOT) );
inv1 gate( .a(N17), .O(N17_NOT) );
and2 gate( .a(N17), .b(D_162_NOT), .O(ED_810) );
and2 gate( .a(N17_NOT), .b(D_162_NOT), .O(ED_811) );
and2 gate( .a(CONST1), .b(D_162), .O(ED_812) );
and2 gate( .a(CONST0), .b(D_162), .O(ED_813) );
and2 gate( .a(ED_810), .b(D_163_NOT), .O(ED_819) );
and2 gate( .a(ED_811), .b(D_163), .O(ED_817) );
and2 gate( .a(ED_812), .b(D_163_NOT), .O(ED_815) );
and2 gate( .a(ED_813), .b(D_163), .O(ED_814) );
or2  gate( .a(ED_814), .b(ED_815), .O(ED_816) );
or2  gate( .a(ED_816), .b(ED_817), .O(ED_818) );
or2  gate( .a(ED_819), .b(ED_818), .O(N17_OBF) );
inv1 gate( .a(D_164), .O(D_164_NOT) );
inv1 gate( .a(D_165), .O(D_165_NOT) );
inv1 gate( .a(N112), .O(N112_NOT) );
and2 gate( .a(N112), .b(D_164_NOT), .O(ED_820) );
and2 gate( .a(N112_NOT), .b(D_164_NOT), .O(ED_821) );
and2 gate( .a(CONST1), .b(D_164), .O(ED_822) );
and2 gate( .a(CONST0), .b(D_164), .O(ED_823) );
and2 gate( .a(ED_820), .b(D_165_NOT), .O(ED_829) );
and2 gate( .a(ED_821), .b(D_165), .O(ED_827) );
and2 gate( .a(ED_822), .b(D_165_NOT), .O(ED_825) );
and2 gate( .a(ED_823), .b(D_165), .O(ED_824) );
or2  gate( .a(ED_824), .b(ED_825), .O(ED_826) );
or2  gate( .a(ED_826), .b(ED_827), .O(ED_828) );
or2  gate( .a(ED_829), .b(ED_828), .O(N112_OBF) );
inv1 gate( .a(D_166), .O(D_166_NOT) );
inv1 gate( .a(D_167), .O(D_167_NOT) );
inv1 gate( .a(N243), .O(N243_NOT) );
and2 gate( .a(N243), .b(D_166_NOT), .O(ED_830) );
and2 gate( .a(N243_NOT), .b(D_166_NOT), .O(ED_831) );
and2 gate( .a(CONST1), .b(D_166), .O(ED_832) );
and2 gate( .a(CONST0), .b(D_166), .O(ED_833) );
and2 gate( .a(ED_830), .b(D_167_NOT), .O(ED_839) );
and2 gate( .a(ED_831), .b(D_167), .O(ED_837) );
and2 gate( .a(ED_832), .b(D_167_NOT), .O(ED_835) );
and2 gate( .a(ED_833), .b(D_167), .O(ED_834) );
or2  gate( .a(ED_834), .b(ED_835), .O(ED_836) );
or2  gate( .a(ED_836), .b(ED_837), .O(ED_838) );
or2  gate( .a(ED_839), .b(ED_838), .O(N243_OBF) );
inv1 gate( .a(D_168), .O(D_168_NOT) );
inv1 gate( .a(D_169), .O(D_169_NOT) );
inv1 gate( .a(N174), .O(N174_NOT) );
and2 gate( .a(N174), .b(D_168_NOT), .O(ED_840) );
and2 gate( .a(N174_NOT), .b(D_168_NOT), .O(ED_841) );
and2 gate( .a(CONST1), .b(D_168), .O(ED_842) );
and2 gate( .a(CONST0), .b(D_168), .O(ED_843) );
and2 gate( .a(ED_840), .b(D_169_NOT), .O(ED_849) );
and2 gate( .a(ED_841), .b(D_169), .O(ED_847) );
and2 gate( .a(ED_842), .b(D_169_NOT), .O(ED_845) );
and2 gate( .a(ED_843), .b(D_169), .O(ED_844) );
or2  gate( .a(ED_844), .b(ED_845), .O(ED_846) );
or2  gate( .a(ED_846), .b(ED_847), .O(ED_848) );
or2  gate( .a(ED_849), .b(ED_848), .O(N174_OBF) );
inv1 gate( .a(D_170), .O(D_170_NOT) );
inv1 gate( .a(D_171), .O(D_171_NOT) );
inv1 gate( .a(N213), .O(N213_NOT) );
and2 gate( .a(N213), .b(D_170_NOT), .O(ED_850) );
and2 gate( .a(N213_NOT), .b(D_170_NOT), .O(ED_851) );
and2 gate( .a(CONST1), .b(D_170), .O(ED_852) );
and2 gate( .a(CONST0), .b(D_170), .O(ED_853) );
and2 gate( .a(ED_850), .b(D_171_NOT), .O(ED_859) );
and2 gate( .a(ED_851), .b(D_171), .O(ED_857) );
and2 gate( .a(ED_852), .b(D_171_NOT), .O(ED_855) );
and2 gate( .a(ED_853), .b(D_171), .O(ED_854) );
or2  gate( .a(ED_854), .b(ED_855), .O(ED_856) );
or2  gate( .a(ED_856), .b(ED_857), .O(ED_858) );
or2  gate( .a(ED_859), .b(ED_858), .O(N213_OBF) );
inv1 gate( .a(D_172), .O(D_172_NOT) );
inv1 gate( .a(D_173), .O(D_173_NOT) );
inv1 gate( .a(N333), .O(N333_NOT) );
and2 gate( .a(N333), .b(D_172_NOT), .O(ED_860) );
and2 gate( .a(N333_NOT), .b(D_172_NOT), .O(ED_861) );
and2 gate( .a(CONST1), .b(D_172), .O(ED_862) );
and2 gate( .a(CONST0), .b(D_172), .O(ED_863) );
and2 gate( .a(ED_860), .b(D_173_NOT), .O(ED_869) );
and2 gate( .a(ED_861), .b(D_173), .O(ED_867) );
and2 gate( .a(ED_862), .b(D_173_NOT), .O(ED_865) );
and2 gate( .a(ED_863), .b(D_173), .O(ED_864) );
or2  gate( .a(ED_864), .b(ED_865), .O(ED_866) );
or2  gate( .a(ED_866), .b(ED_867), .O(ED_868) );
or2  gate( .a(ED_869), .b(ED_868), .O(N333_OBF) );
inv1 gate( .a(D_174), .O(D_174_NOT) );
inv1 gate( .a(D_175), .O(D_175_NOT) );
inv1 gate( .a(N213), .O(N213_NOT) );
and2 gate( .a(N213), .b(D_174_NOT), .O(ED_870) );
and2 gate( .a(N213_NOT), .b(D_174_NOT), .O(ED_871) );
and2 gate( .a(CONST1), .b(D_174), .O(ED_872) );
and2 gate( .a(CONST0), .b(D_174), .O(ED_873) );
and2 gate( .a(ED_870), .b(D_175_NOT), .O(ED_879) );
and2 gate( .a(ED_871), .b(D_175), .O(ED_877) );
and2 gate( .a(ED_872), .b(D_175_NOT), .O(ED_875) );
and2 gate( .a(ED_873), .b(D_175), .O(ED_874) );
or2  gate( .a(ED_874), .b(ED_875), .O(ED_876) );
or2  gate( .a(ED_876), .b(ED_877), .O(ED_878) );
or2  gate( .a(ED_879), .b(ED_878), .O(N213_OBF) );
inv1 gate( .a(D_176), .O(D_176_NOT) );
inv1 gate( .a(D_177), .O(D_177_NOT) );
inv1 gate( .a(N76), .O(N76_NOT) );
and2 gate( .a(N76), .b(D_176_NOT), .O(ED_880) );
and2 gate( .a(N76_NOT), .b(D_176_NOT), .O(ED_881) );
and2 gate( .a(CONST1), .b(D_176), .O(ED_882) );
and2 gate( .a(CONST0), .b(D_176), .O(ED_883) );
and2 gate( .a(ED_880), .b(D_177_NOT), .O(ED_889) );
and2 gate( .a(ED_881), .b(D_177), .O(ED_887) );
and2 gate( .a(ED_882), .b(D_177_NOT), .O(ED_885) );
and2 gate( .a(ED_883), .b(D_177), .O(ED_884) );
or2  gate( .a(ED_884), .b(ED_885), .O(ED_886) );
or2  gate( .a(ED_886), .b(ED_887), .O(ED_888) );
or2  gate( .a(ED_889), .b(ED_888), .O(N76_OBF) );
inv1 gate( .a(D_178), .O(D_178_NOT) );
inv1 gate( .a(D_179), .O(D_179_NOT) );
inv1 gate( .a(N1), .O(N1_NOT) );
and2 gate( .a(N1), .b(D_178_NOT), .O(ED_890) );
and2 gate( .a(N1_NOT), .b(D_178_NOT), .O(ED_891) );
and2 gate( .a(CONST1), .b(D_178), .O(ED_892) );
and2 gate( .a(CONST0), .b(D_178), .O(ED_893) );
and2 gate( .a(ED_890), .b(D_179_NOT), .O(ED_899) );
and2 gate( .a(ED_891), .b(D_179), .O(ED_897) );
and2 gate( .a(ED_892), .b(D_179_NOT), .O(ED_895) );
and2 gate( .a(ED_893), .b(D_179), .O(ED_894) );
or2  gate( .a(ED_894), .b(ED_895), .O(ED_896) );
or2  gate( .a(ED_896), .b(ED_897), .O(ED_898) );
or2  gate( .a(ED_899), .b(ED_898), .O(N1_OBF) );
inv1 gate( .a(D_180), .O(D_180_NOT) );
inv1 gate( .a(D_181), .O(D_181_NOT) );
inv1 gate( .a(N307), .O(N307_NOT) );
and2 gate( .a(N307), .b(D_180_NOT), .O(ED_900) );
and2 gate( .a(N307_NOT), .b(D_180_NOT), .O(ED_901) );
and2 gate( .a(CONST1), .b(D_180), .O(ED_902) );
and2 gate( .a(CONST0), .b(D_180), .O(ED_903) );
and2 gate( .a(ED_900), .b(D_181_NOT), .O(ED_909) );
and2 gate( .a(ED_901), .b(D_181), .O(ED_907) );
and2 gate( .a(ED_902), .b(D_181_NOT), .O(ED_905) );
and2 gate( .a(ED_903), .b(D_181), .O(ED_904) );
or2  gate( .a(ED_904), .b(ED_905), .O(ED_906) );
or2  gate( .a(ED_906), .b(ED_907), .O(ED_908) );
or2  gate( .a(ED_909), .b(ED_908), .O(N307_OBF) );
inv1 gate( .a(D_182), .O(D_182_NOT) );
inv1 gate( .a(D_183), .O(D_183_NOT) );
inv1 gate( .a(N190), .O(N190_NOT) );
and2 gate( .a(N190), .b(D_182_NOT), .O(ED_910) );
and2 gate( .a(N190_NOT), .b(D_182_NOT), .O(ED_911) );
and2 gate( .a(CONST1), .b(D_182), .O(ED_912) );
and2 gate( .a(CONST0), .b(D_182), .O(ED_913) );
and2 gate( .a(ED_910), .b(D_183_NOT), .O(ED_919) );
and2 gate( .a(ED_911), .b(D_183), .O(ED_917) );
and2 gate( .a(ED_912), .b(D_183_NOT), .O(ED_915) );
and2 gate( .a(ED_913), .b(D_183), .O(ED_914) );
or2  gate( .a(ED_914), .b(ED_915), .O(ED_916) );
or2  gate( .a(ED_916), .b(ED_917), .O(ED_918) );
or2  gate( .a(ED_919), .b(ED_918), .O(N190_OBF) );
inv1 gate( .a(D_184), .O(D_184_NOT) );
inv1 gate( .a(D_185), .O(D_185_NOT) );
inv1 gate( .a(N147), .O(N147_NOT) );
and2 gate( .a(N147), .b(D_184_NOT), .O(ED_920) );
and2 gate( .a(N147_NOT), .b(D_184_NOT), .O(ED_921) );
and2 gate( .a(CONST1), .b(D_184), .O(ED_922) );
and2 gate( .a(CONST0), .b(D_184), .O(ED_923) );
and2 gate( .a(ED_920), .b(D_185_NOT), .O(ED_929) );
and2 gate( .a(ED_921), .b(D_185), .O(ED_927) );
and2 gate( .a(ED_922), .b(D_185_NOT), .O(ED_925) );
and2 gate( .a(ED_923), .b(D_185), .O(ED_924) );
or2  gate( .a(ED_924), .b(ED_925), .O(ED_926) );
or2  gate( .a(ED_926), .b(ED_927), .O(ED_928) );
or2  gate( .a(ED_929), .b(ED_928), .O(N147_OBF) );
inv1 gate( .a(D_186), .O(D_186_NOT) );
inv1 gate( .a(D_187), .O(D_187_NOT) );
inv1 gate( .a(N184), .O(N184_NOT) );
and2 gate( .a(N184), .b(D_186_NOT), .O(ED_930) );
and2 gate( .a(N184_NOT), .b(D_186_NOT), .O(ED_931) );
and2 gate( .a(CONST1), .b(D_186), .O(ED_932) );
and2 gate( .a(CONST0), .b(D_186), .O(ED_933) );
and2 gate( .a(ED_930), .b(D_187_NOT), .O(ED_939) );
and2 gate( .a(ED_931), .b(D_187), .O(ED_937) );
and2 gate( .a(ED_932), .b(D_187_NOT), .O(ED_935) );
and2 gate( .a(ED_933), .b(D_187), .O(ED_934) );
or2  gate( .a(ED_934), .b(ED_935), .O(ED_936) );
or2  gate( .a(ED_936), .b(ED_937), .O(ED_938) );
or2  gate( .a(ED_939), .b(ED_938), .O(N184_OBF) );
inv1 gate( .a(D_188), .O(D_188_NOT) );
inv1 gate( .a(D_189), .O(D_189_NOT) );
inv1 gate( .a(N319), .O(N319_NOT) );
and2 gate( .a(N319), .b(D_188_NOT), .O(ED_940) );
and2 gate( .a(N319_NOT), .b(D_188_NOT), .O(ED_941) );
and2 gate( .a(CONST1), .b(D_188), .O(ED_942) );
and2 gate( .a(CONST0), .b(D_188), .O(ED_943) );
and2 gate( .a(ED_940), .b(D_189_NOT), .O(ED_949) );
and2 gate( .a(ED_941), .b(D_189), .O(ED_947) );
and2 gate( .a(ED_942), .b(D_189_NOT), .O(ED_945) );
and2 gate( .a(ED_943), .b(D_189), .O(ED_944) );
or2  gate( .a(ED_944), .b(ED_945), .O(ED_946) );
or2  gate( .a(ED_946), .b(ED_947), .O(ED_948) );
or2  gate( .a(ED_949), .b(ED_948), .O(N319_OBF) );
inv1 gate( .a(D_190), .O(D_190_NOT) );
inv1 gate( .a(D_191), .O(D_191_NOT) );
inv1 gate( .a(N143), .O(N143_NOT) );
and2 gate( .a(N143), .b(D_190_NOT), .O(ED_950) );
and2 gate( .a(N143_NOT), .b(D_190_NOT), .O(ED_951) );
and2 gate( .a(CONST1), .b(D_190), .O(ED_952) );
and2 gate( .a(CONST0), .b(D_190), .O(ED_953) );
and2 gate( .a(ED_950), .b(D_191_NOT), .O(ED_959) );
and2 gate( .a(ED_951), .b(D_191), .O(ED_957) );
and2 gate( .a(ED_952), .b(D_191_NOT), .O(ED_955) );
and2 gate( .a(ED_953), .b(D_191), .O(ED_954) );
or2  gate( .a(ED_954), .b(ED_955), .O(ED_956) );
or2  gate( .a(ED_956), .b(ED_957), .O(ED_958) );
or2  gate( .a(ED_959), .b(ED_958), .O(N143_OBF) );
inv1 gate( .a(D_192), .O(D_192_NOT) );
inv1 gate( .a(D_193), .O(D_193_NOT) );
inv1 gate( .a(N374), .O(N374_NOT) );
and2 gate( .a(N374), .b(D_192_NOT), .O(ED_960) );
and2 gate( .a(N374_NOT), .b(D_192_NOT), .O(ED_961) );
and2 gate( .a(CONST1), .b(D_192), .O(ED_962) );
and2 gate( .a(CONST0), .b(D_192), .O(ED_963) );
and2 gate( .a(ED_960), .b(D_193_NOT), .O(ED_969) );
and2 gate( .a(ED_961), .b(D_193), .O(ED_967) );
and2 gate( .a(ED_962), .b(D_193_NOT), .O(ED_965) );
and2 gate( .a(ED_963), .b(D_193), .O(ED_964) );
or2  gate( .a(ED_964), .b(ED_965), .O(ED_966) );
or2  gate( .a(ED_966), .b(ED_967), .O(ED_968) );
or2  gate( .a(ED_969), .b(ED_968), .O(N374_OBF) );
inv1 gate( .a(D_194), .O(D_194_NOT) );
inv1 gate( .a(D_195), .O(D_195_NOT) );
inv1 gate( .a(N194), .O(N194_NOT) );
and2 gate( .a(N194), .b(D_194_NOT), .O(ED_970) );
and2 gate( .a(N194_NOT), .b(D_194_NOT), .O(ED_971) );
and2 gate( .a(CONST1), .b(D_194), .O(ED_972) );
and2 gate( .a(CONST0), .b(D_194), .O(ED_973) );
and2 gate( .a(ED_970), .b(D_195_NOT), .O(ED_979) );
and2 gate( .a(ED_971), .b(D_195), .O(ED_977) );
and2 gate( .a(ED_972), .b(D_195_NOT), .O(ED_975) );
and2 gate( .a(ED_973), .b(D_195), .O(ED_974) );
or2  gate( .a(ED_974), .b(ED_975), .O(ED_976) );
or2  gate( .a(ED_976), .b(ED_977), .O(ED_978) );
or2  gate( .a(ED_979), .b(ED_978), .O(N194_OBF) );
inv1 gate( .a(D_196), .O(D_196_NOT) );
inv1 gate( .a(D_197), .O(D_197_NOT) );
inv1 gate( .a(N346), .O(N346_NOT) );
and2 gate( .a(N346), .b(D_196_NOT), .O(ED_980) );
and2 gate( .a(N346_NOT), .b(D_196_NOT), .O(ED_981) );
and2 gate( .a(CONST1), .b(D_196), .O(ED_982) );
and2 gate( .a(CONST0), .b(D_196), .O(ED_983) );
and2 gate( .a(ED_980), .b(D_197_NOT), .O(ED_989) );
and2 gate( .a(ED_981), .b(D_197), .O(ED_987) );
and2 gate( .a(ED_982), .b(D_197_NOT), .O(ED_985) );
and2 gate( .a(ED_983), .b(D_197), .O(ED_984) );
or2  gate( .a(ED_984), .b(ED_985), .O(ED_986) );
or2  gate( .a(ED_986), .b(ED_987), .O(ED_988) );
or2  gate( .a(ED_989), .b(ED_988), .O(N346_OBF) );
inv1 gate( .a(D_198), .O(D_198_NOT) );
inv1 gate( .a(D_199), .O(D_199_NOT) );
inv1 gate( .a(N386), .O(N386_NOT) );
and2 gate( .a(N386), .b(D_198_NOT), .O(ED_990) );
and2 gate( .a(N386_NOT), .b(D_198_NOT), .O(ED_991) );
and2 gate( .a(CONST1), .b(D_198), .O(ED_992) );
and2 gate( .a(CONST0), .b(D_198), .O(ED_993) );
and2 gate( .a(ED_990), .b(D_199_NOT), .O(ED_999) );
and2 gate( .a(ED_991), .b(D_199), .O(ED_997) );
and2 gate( .a(ED_992), .b(D_199_NOT), .O(ED_995) );
and2 gate( .a(ED_993), .b(D_199), .O(ED_994) );
or2  gate( .a(ED_994), .b(ED_995), .O(ED_996) );
or2  gate( .a(ED_996), .b(ED_997), .O(ED_998) );
or2  gate( .a(ED_999), .b(ED_998), .O(N386_OBF) );
inv1 gate( .a(D_200), .O(D_200_NOT) );
inv1 gate( .a(D_201), .O(D_201_NOT) );
inv1 gate( .a(N349), .O(N349_NOT) );
and2 gate( .a(N349), .b(D_200_NOT), .O(ED_1000) );
and2 gate( .a(N349_NOT), .b(D_200_NOT), .O(ED_1001) );
and2 gate( .a(CONST1), .b(D_200), .O(ED_1002) );
and2 gate( .a(CONST0), .b(D_200), .O(ED_1003) );
and2 gate( .a(ED_1000), .b(D_201_NOT), .O(ED_1009) );
and2 gate( .a(ED_1001), .b(D_201), .O(ED_1007) );
and2 gate( .a(ED_1002), .b(D_201_NOT), .O(ED_1005) );
and2 gate( .a(ED_1003), .b(D_201), .O(ED_1004) );
or2  gate( .a(ED_1004), .b(ED_1005), .O(ED_1006) );
or2  gate( .a(ED_1006), .b(ED_1007), .O(ED_1008) );
or2  gate( .a(ED_1009), .b(ED_1008), .O(N349_OBF) );
inv1 gate( .a(D_202), .O(D_202_NOT) );
inv1 gate( .a(D_203), .O(D_203_NOT) );
inv1 gate( .a(N411), .O(N411_NOT) );
and2 gate( .a(N411), .b(D_202_NOT), .O(ED_1010) );
and2 gate( .a(N411_NOT), .b(D_202_NOT), .O(ED_1011) );
and2 gate( .a(CONST1), .b(D_202), .O(ED_1012) );
and2 gate( .a(CONST0), .b(D_202), .O(ED_1013) );
and2 gate( .a(ED_1010), .b(D_203_NOT), .O(ED_1019) );
and2 gate( .a(ED_1011), .b(D_203), .O(ED_1017) );
and2 gate( .a(ED_1012), .b(D_203_NOT), .O(ED_1015) );
and2 gate( .a(ED_1013), .b(D_203), .O(ED_1014) );
or2  gate( .a(ED_1014), .b(ED_1015), .O(ED_1016) );
or2  gate( .a(ED_1016), .b(ED_1017), .O(ED_1018) );
or2  gate( .a(ED_1019), .b(ED_1018), .O(N411_OBF) );
inv1 gate( .a(D_204), .O(D_204_NOT) );
inv1 gate( .a(D_205), .O(D_205_NOT) );
inv1 gate( .a(N185), .O(N185_NOT) );
and2 gate( .a(N185), .b(D_204_NOT), .O(ED_1020) );
and2 gate( .a(N185_NOT), .b(D_204_NOT), .O(ED_1021) );
and2 gate( .a(CONST1), .b(D_204), .O(ED_1022) );
and2 gate( .a(CONST0), .b(D_204), .O(ED_1023) );
and2 gate( .a(ED_1020), .b(D_205_NOT), .O(ED_1029) );
and2 gate( .a(ED_1021), .b(D_205), .O(ED_1027) );
and2 gate( .a(ED_1022), .b(D_205_NOT), .O(ED_1025) );
and2 gate( .a(ED_1023), .b(D_205), .O(ED_1024) );
or2  gate( .a(ED_1024), .b(ED_1025), .O(ED_1026) );
or2  gate( .a(ED_1026), .b(ED_1027), .O(ED_1028) );
or2  gate( .a(ED_1029), .b(ED_1028), .O(N185_OBF) );
inv1 gate( .a(D_206), .O(D_206_NOT) );
inv1 gate( .a(D_207), .O(D_207_NOT) );
inv1 gate( .a(N60), .O(N60_NOT) );
and2 gate( .a(N60), .b(D_206_NOT), .O(ED_1030) );
and2 gate( .a(N60_NOT), .b(D_206_NOT), .O(ED_1031) );
and2 gate( .a(CONST1), .b(D_206), .O(ED_1032) );
and2 gate( .a(CONST0), .b(D_206), .O(ED_1033) );
and2 gate( .a(ED_1030), .b(D_207_NOT), .O(ED_1039) );
and2 gate( .a(ED_1031), .b(D_207), .O(ED_1037) );
and2 gate( .a(ED_1032), .b(D_207_NOT), .O(ED_1035) );
and2 gate( .a(ED_1033), .b(D_207), .O(ED_1034) );
or2  gate( .a(ED_1034), .b(ED_1035), .O(ED_1036) );
or2  gate( .a(ED_1036), .b(ED_1037), .O(ED_1038) );
or2  gate( .a(ED_1039), .b(ED_1038), .O(N60_OBF) );
inv1 gate( .a(D_208), .O(D_208_NOT) );
inv1 gate( .a(D_209), .O(D_209_NOT) );
inv1 gate( .a(N289), .O(N289_NOT) );
and2 gate( .a(N289), .b(D_208_NOT), .O(ED_1040) );
and2 gate( .a(N289_NOT), .b(D_208_NOT), .O(ED_1041) );
and2 gate( .a(CONST1), .b(D_208), .O(ED_1042) );
and2 gate( .a(CONST0), .b(D_208), .O(ED_1043) );
and2 gate( .a(ED_1040), .b(D_209_NOT), .O(ED_1049) );
and2 gate( .a(ED_1041), .b(D_209), .O(ED_1047) );
and2 gate( .a(ED_1042), .b(D_209_NOT), .O(ED_1045) );
and2 gate( .a(ED_1043), .b(D_209), .O(ED_1044) );
or2  gate( .a(ED_1044), .b(ED_1045), .O(ED_1046) );
or2  gate( .a(ED_1046), .b(ED_1047), .O(ED_1048) );
or2  gate( .a(ED_1049), .b(ED_1048), .O(N289_OBF) );
inv1 gate( .a(D_210), .O(D_210_NOT) );
inv1 gate( .a(D_211), .O(D_211_NOT) );
inv1 gate( .a(N21), .O(N21_NOT) );
and2 gate( .a(N21), .b(D_210_NOT), .O(ED_1050) );
and2 gate( .a(N21_NOT), .b(D_210_NOT), .O(ED_1051) );
and2 gate( .a(CONST1), .b(D_210), .O(ED_1052) );
and2 gate( .a(CONST0), .b(D_210), .O(ED_1053) );
and2 gate( .a(ED_1050), .b(D_211_NOT), .O(ED_1059) );
and2 gate( .a(ED_1051), .b(D_211), .O(ED_1057) );
and2 gate( .a(ED_1052), .b(D_211_NOT), .O(ED_1055) );
and2 gate( .a(ED_1053), .b(D_211), .O(ED_1054) );
or2  gate( .a(ED_1054), .b(ED_1055), .O(ED_1056) );
or2  gate( .a(ED_1056), .b(ED_1057), .O(ED_1058) );
or2  gate( .a(ED_1059), .b(ED_1058), .O(N21_OBF) );
inv1 gate( .a(D_212), .O(D_212_NOT) );
inv1 gate( .a(D_213), .O(D_213_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_212_NOT), .O(ED_1060) );
and2 gate( .a(N360_NOT), .b(D_212_NOT), .O(ED_1061) );
and2 gate( .a(CONST1), .b(D_212), .O(ED_1062) );
and2 gate( .a(CONST0), .b(D_212), .O(ED_1063) );
and2 gate( .a(ED_1060), .b(D_213_NOT), .O(ED_1069) );
and2 gate( .a(ED_1061), .b(D_213), .O(ED_1067) );
and2 gate( .a(ED_1062), .b(D_213_NOT), .O(ED_1065) );
and2 gate( .a(ED_1063), .b(D_213), .O(ED_1064) );
or2  gate( .a(ED_1064), .b(ED_1065), .O(ED_1066) );
or2  gate( .a(ED_1066), .b(ED_1067), .O(ED_1068) );
or2  gate( .a(ED_1069), .b(ED_1068), .O(N360_OBF) );
inv1 gate( .a(D_214), .O(D_214_NOT) );
inv1 gate( .a(D_215), .O(D_215_NOT) );
inv1 gate( .a(N372), .O(N372_NOT) );
and2 gate( .a(N372), .b(D_214_NOT), .O(ED_1070) );
and2 gate( .a(N372_NOT), .b(D_214_NOT), .O(ED_1071) );
and2 gate( .a(CONST1), .b(D_214), .O(ED_1072) );
and2 gate( .a(CONST0), .b(D_214), .O(ED_1073) );
and2 gate( .a(ED_1070), .b(D_215_NOT), .O(ED_1079) );
and2 gate( .a(ED_1071), .b(D_215), .O(ED_1077) );
and2 gate( .a(ED_1072), .b(D_215_NOT), .O(ED_1075) );
and2 gate( .a(ED_1073), .b(D_215), .O(ED_1074) );
or2  gate( .a(ED_1074), .b(ED_1075), .O(ED_1076) );
or2  gate( .a(ED_1076), .b(ED_1077), .O(ED_1078) );
or2  gate( .a(ED_1079), .b(ED_1078), .O(N372_OBF) );
inv1 gate( .a(D_216), .O(D_216_NOT) );
inv1 gate( .a(D_217), .O(D_217_NOT) );
inv1 gate( .a(N213), .O(N213_NOT) );
and2 gate( .a(N213), .b(D_216_NOT), .O(ED_1080) );
and2 gate( .a(N213_NOT), .b(D_216_NOT), .O(ED_1081) );
and2 gate( .a(CONST1), .b(D_216), .O(ED_1082) );
and2 gate( .a(CONST0), .b(D_216), .O(ED_1083) );
and2 gate( .a(ED_1080), .b(D_217_NOT), .O(ED_1089) );
and2 gate( .a(ED_1081), .b(D_217), .O(ED_1087) );
and2 gate( .a(ED_1082), .b(D_217_NOT), .O(ED_1085) );
and2 gate( .a(ED_1083), .b(D_217), .O(ED_1084) );
or2  gate( .a(ED_1084), .b(ED_1085), .O(ED_1086) );
or2  gate( .a(ED_1086), .b(ED_1087), .O(ED_1088) );
or2  gate( .a(ED_1089), .b(ED_1088), .O(N213_OBF) );
inv1 gate( .a(D_218), .O(D_218_NOT) );
inv1 gate( .a(D_219), .O(D_219_NOT) );
inv1 gate( .a(N115), .O(N115_NOT) );
and2 gate( .a(N115), .b(D_218_NOT), .O(ED_1090) );
and2 gate( .a(N115_NOT), .b(D_218_NOT), .O(ED_1091) );
and2 gate( .a(CONST1), .b(D_218), .O(ED_1092) );
and2 gate( .a(CONST0), .b(D_218), .O(ED_1093) );
and2 gate( .a(ED_1090), .b(D_219_NOT), .O(ED_1099) );
and2 gate( .a(ED_1091), .b(D_219), .O(ED_1097) );
and2 gate( .a(ED_1092), .b(D_219_NOT), .O(ED_1095) );
and2 gate( .a(ED_1093), .b(D_219), .O(ED_1094) );
or2  gate( .a(ED_1094), .b(ED_1095), .O(ED_1096) );
or2  gate( .a(ED_1096), .b(ED_1097), .O(ED_1098) );
or2  gate( .a(ED_1099), .b(ED_1098), .O(N115_OBF) );
inv1 gate( .a(D_220), .O(D_220_NOT) );
inv1 gate( .a(D_221), .O(D_221_NOT) );
inv1 gate( .a(N267), .O(N267_NOT) );
and2 gate( .a(N267), .b(D_220_NOT), .O(ED_1100) );
and2 gate( .a(N267_NOT), .b(D_220_NOT), .O(ED_1101) );
and2 gate( .a(CONST1), .b(D_220), .O(ED_1102) );
and2 gate( .a(CONST0), .b(D_220), .O(ED_1103) );
and2 gate( .a(ED_1100), .b(D_221_NOT), .O(ED_1109) );
and2 gate( .a(ED_1101), .b(D_221), .O(ED_1107) );
and2 gate( .a(ED_1102), .b(D_221_NOT), .O(ED_1105) );
and2 gate( .a(ED_1103), .b(D_221), .O(ED_1104) );
or2  gate( .a(ED_1104), .b(ED_1105), .O(ED_1106) );
or2  gate( .a(ED_1106), .b(ED_1107), .O(ED_1108) );
or2  gate( .a(ED_1109), .b(ED_1108), .O(N267_OBF) );
inv1 gate( .a(D_222), .O(D_222_NOT) );
inv1 gate( .a(D_223), .O(D_223_NOT) );
inv1 gate( .a(N158), .O(N158_NOT) );
and2 gate( .a(N158), .b(D_222_NOT), .O(ED_1110) );
and2 gate( .a(N158_NOT), .b(D_222_NOT), .O(ED_1111) );
and2 gate( .a(CONST1), .b(D_222), .O(ED_1112) );
and2 gate( .a(CONST0), .b(D_222), .O(ED_1113) );
and2 gate( .a(ED_1110), .b(D_223_NOT), .O(ED_1119) );
and2 gate( .a(ED_1111), .b(D_223), .O(ED_1117) );
and2 gate( .a(ED_1112), .b(D_223_NOT), .O(ED_1115) );
and2 gate( .a(ED_1113), .b(D_223), .O(ED_1114) );
or2  gate( .a(ED_1114), .b(ED_1115), .O(ED_1116) );
or2  gate( .a(ED_1116), .b(ED_1117), .O(ED_1118) );
or2  gate( .a(ED_1119), .b(ED_1118), .O(N158_OBF) );
inv1 gate( .a(D_224), .O(D_224_NOT) );
inv1 gate( .a(D_225), .O(D_225_NOT) );
inv1 gate( .a(N239), .O(N239_NOT) );
and2 gate( .a(N239), .b(D_224_NOT), .O(ED_1120) );
and2 gate( .a(N239_NOT), .b(D_224_NOT), .O(ED_1121) );
and2 gate( .a(CONST1), .b(D_224), .O(ED_1122) );
and2 gate( .a(CONST0), .b(D_224), .O(ED_1123) );
and2 gate( .a(ED_1120), .b(D_225_NOT), .O(ED_1129) );
and2 gate( .a(ED_1121), .b(D_225), .O(ED_1127) );
and2 gate( .a(ED_1122), .b(D_225_NOT), .O(ED_1125) );
and2 gate( .a(ED_1123), .b(D_225), .O(ED_1124) );
or2  gate( .a(ED_1124), .b(ED_1125), .O(ED_1126) );
or2  gate( .a(ED_1126), .b(ED_1127), .O(ED_1128) );
or2  gate( .a(ED_1129), .b(ED_1128), .O(N239_OBF) );
inv1 gate( .a(D_226), .O(D_226_NOT) );
inv1 gate( .a(D_227), .O(D_227_NOT) );
inv1 gate( .a(N1), .O(N1_NOT) );
and2 gate( .a(N1), .b(D_226_NOT), .O(ED_1130) );
and2 gate( .a(N1_NOT), .b(D_226_NOT), .O(ED_1131) );
and2 gate( .a(CONST1), .b(D_226), .O(ED_1132) );
and2 gate( .a(CONST0), .b(D_226), .O(ED_1133) );
and2 gate( .a(ED_1130), .b(D_227_NOT), .O(ED_1139) );
and2 gate( .a(ED_1131), .b(D_227), .O(ED_1137) );
and2 gate( .a(ED_1132), .b(D_227_NOT), .O(ED_1135) );
and2 gate( .a(ED_1133), .b(D_227), .O(ED_1134) );
or2  gate( .a(ED_1134), .b(ED_1135), .O(ED_1136) );
or2  gate( .a(ED_1136), .b(ED_1137), .O(ED_1138) );
or2  gate( .a(ED_1139), .b(ED_1138), .O(N1_OBF) );
inv1 gate( .a(D_228), .O(D_228_NOT) );
inv1 gate( .a(D_229), .O(D_229_NOT) );
inv1 gate( .a(N187), .O(N187_NOT) );
and2 gate( .a(N187), .b(D_228_NOT), .O(ED_1140) );
and2 gate( .a(N187_NOT), .b(D_228_NOT), .O(ED_1141) );
and2 gate( .a(CONST1), .b(D_228), .O(ED_1142) );
and2 gate( .a(CONST0), .b(D_228), .O(ED_1143) );
and2 gate( .a(ED_1140), .b(D_229_NOT), .O(ED_1149) );
and2 gate( .a(ED_1141), .b(D_229), .O(ED_1147) );
and2 gate( .a(ED_1142), .b(D_229_NOT), .O(ED_1145) );
and2 gate( .a(ED_1143), .b(D_229), .O(ED_1144) );
or2  gate( .a(ED_1144), .b(ED_1145), .O(ED_1146) );
or2  gate( .a(ED_1146), .b(ED_1147), .O(ED_1148) );
or2  gate( .a(ED_1149), .b(ED_1148), .O(N187_OBF) );
inv1 gate( .a(D_230), .O(D_230_NOT) );
inv1 gate( .a(D_231), .O(D_231_NOT) );
inv1 gate( .a(N63), .O(N63_NOT) );
and2 gate( .a(N63), .b(D_230_NOT), .O(ED_1150) );
and2 gate( .a(N63_NOT), .b(D_230_NOT), .O(ED_1151) );
and2 gate( .a(CONST1), .b(D_230), .O(ED_1152) );
and2 gate( .a(CONST0), .b(D_230), .O(ED_1153) );
and2 gate( .a(ED_1150), .b(D_231_NOT), .O(ED_1159) );
and2 gate( .a(ED_1151), .b(D_231), .O(ED_1157) );
and2 gate( .a(ED_1152), .b(D_231_NOT), .O(ED_1155) );
and2 gate( .a(ED_1153), .b(D_231), .O(ED_1154) );
or2  gate( .a(ED_1154), .b(ED_1155), .O(ED_1156) );
or2  gate( .a(ED_1156), .b(ED_1157), .O(ED_1158) );
or2  gate( .a(ED_1159), .b(ED_1158), .O(N63_OBF) );
inv1 gate( .a(D_232), .O(D_232_NOT) );
inv1 gate( .a(D_233), .O(D_233_NOT) );
inv1 gate( .a(N381), .O(N381_NOT) );
and2 gate( .a(N381), .b(D_232_NOT), .O(ED_1160) );
and2 gate( .a(N381_NOT), .b(D_232_NOT), .O(ED_1161) );
and2 gate( .a(CONST1), .b(D_232), .O(ED_1162) );
and2 gate( .a(CONST0), .b(D_232), .O(ED_1163) );
and2 gate( .a(ED_1160), .b(D_233_NOT), .O(ED_1169) );
and2 gate( .a(ED_1161), .b(D_233), .O(ED_1167) );
and2 gate( .a(ED_1162), .b(D_233_NOT), .O(ED_1165) );
and2 gate( .a(ED_1163), .b(D_233), .O(ED_1164) );
or2  gate( .a(ED_1164), .b(ED_1165), .O(ED_1166) );
or2  gate( .a(ED_1166), .b(ED_1167), .O(ED_1168) );
or2  gate( .a(ED_1169), .b(ED_1168), .O(N381_OBF) );
inv1 gate( .a(D_234), .O(D_234_NOT) );
inv1 gate( .a(D_235), .O(D_235_NOT) );
inv1 gate( .a(N199), .O(N199_NOT) );
and2 gate( .a(N199), .b(D_234_NOT), .O(ED_1170) );
and2 gate( .a(N199_NOT), .b(D_234_NOT), .O(ED_1171) );
and2 gate( .a(CONST1), .b(D_234), .O(ED_1172) );
and2 gate( .a(CONST0), .b(D_234), .O(ED_1173) );
and2 gate( .a(ED_1170), .b(D_235_NOT), .O(ED_1179) );
and2 gate( .a(ED_1171), .b(D_235), .O(ED_1177) );
and2 gate( .a(ED_1172), .b(D_235_NOT), .O(ED_1175) );
and2 gate( .a(ED_1173), .b(D_235), .O(ED_1174) );
or2  gate( .a(ED_1174), .b(ED_1175), .O(ED_1176) );
or2  gate( .a(ED_1176), .b(ED_1177), .O(ED_1178) );
or2  gate( .a(ED_1179), .b(ED_1178), .O(N199_OBF) );
inv1 gate( .a(D_236), .O(D_236_NOT) );
inv1 gate( .a(D_237), .O(D_237_NOT) );
inv1 gate( .a(N102), .O(N102_NOT) );
and2 gate( .a(N102), .b(D_236_NOT), .O(ED_1180) );
and2 gate( .a(N102_NOT), .b(D_236_NOT), .O(ED_1181) );
and2 gate( .a(CONST1), .b(D_236), .O(ED_1182) );
and2 gate( .a(CONST0), .b(D_236), .O(ED_1183) );
and2 gate( .a(ED_1180), .b(D_237_NOT), .O(ED_1189) );
and2 gate( .a(ED_1181), .b(D_237), .O(ED_1187) );
and2 gate( .a(ED_1182), .b(D_237_NOT), .O(ED_1185) );
and2 gate( .a(ED_1183), .b(D_237), .O(ED_1184) );
or2  gate( .a(ED_1184), .b(ED_1185), .O(ED_1186) );
or2  gate( .a(ED_1186), .b(ED_1187), .O(ED_1188) );
or2  gate( .a(ED_1189), .b(ED_1188), .O(N102_OBF) );
inv1 gate( .a(D_238), .O(D_238_NOT) );
inv1 gate( .a(D_239), .O(D_239_NOT) );
inv1 gate( .a(N108), .O(N108_NOT) );
and2 gate( .a(N108), .b(D_238_NOT), .O(ED_1190) );
and2 gate( .a(N108_NOT), .b(D_238_NOT), .O(ED_1191) );
and2 gate( .a(CONST1), .b(D_238), .O(ED_1192) );
and2 gate( .a(CONST0), .b(D_238), .O(ED_1193) );
and2 gate( .a(ED_1190), .b(D_239_NOT), .O(ED_1199) );
and2 gate( .a(ED_1191), .b(D_239), .O(ED_1197) );
and2 gate( .a(ED_1192), .b(D_239_NOT), .O(ED_1195) );
and2 gate( .a(ED_1193), .b(D_239), .O(ED_1194) );
or2  gate( .a(ED_1194), .b(ED_1195), .O(ED_1196) );
or2  gate( .a(ED_1196), .b(ED_1197), .O(ED_1198) );
or2  gate( .a(ED_1199), .b(ED_1198), .O(N108_OBF) );
inv1 gate( .a(D_240), .O(D_240_NOT) );
inv1 gate( .a(D_241), .O(D_241_NOT) );
inv1 gate( .a(N360), .O(N360_NOT) );
and2 gate( .a(N360), .b(D_240_NOT), .O(ED_1200) );
and2 gate( .a(N360_NOT), .b(D_240_NOT), .O(ED_1201) );
and2 gate( .a(CONST1), .b(D_240), .O(ED_1202) );
and2 gate( .a(CONST0), .b(D_240), .O(ED_1203) );
and2 gate( .a(ED_1200), .b(D_241_NOT), .O(ED_1209) );
and2 gate( .a(ED_1201), .b(D_241), .O(ED_1207) );
and2 gate( .a(ED_1202), .b(D_241_NOT), .O(ED_1205) );
and2 gate( .a(ED_1203), .b(D_241), .O(ED_1204) );
or2  gate( .a(ED_1204), .b(ED_1205), .O(ED_1206) );
or2  gate( .a(ED_1206), .b(ED_1207), .O(ED_1208) );
or2  gate( .a(ED_1209), .b(ED_1208), .O(N360_OBF) );
inv1 gate( .a(D_242), .O(D_242_NOT) );
inv1 gate( .a(D_243), .O(D_243_NOT) );
inv1 gate( .a(N95), .O(N95_NOT) );
and2 gate( .a(N95), .b(D_242_NOT), .O(ED_1210) );
and2 gate( .a(N95_NOT), .b(D_242_NOT), .O(ED_1211) );
and2 gate( .a(CONST1), .b(D_242), .O(ED_1212) );
and2 gate( .a(CONST0), .b(D_242), .O(ED_1213) );
and2 gate( .a(ED_1210), .b(D_243_NOT), .O(ED_1219) );
and2 gate( .a(ED_1211), .b(D_243), .O(ED_1217) );
and2 gate( .a(ED_1212), .b(D_243_NOT), .O(ED_1215) );
and2 gate( .a(ED_1213), .b(D_243), .O(ED_1214) );
or2  gate( .a(ED_1214), .b(ED_1215), .O(ED_1216) );
or2  gate( .a(ED_1216), .b(ED_1217), .O(ED_1218) );
or2  gate( .a(ED_1219), .b(ED_1218), .O(N95_OBF) );
inv1 gate( .a(D_244), .O(D_244_NOT) );
inv1 gate( .a(D_245), .O(D_245_NOT) );
inv1 gate( .a(N43), .O(N43_NOT) );
and2 gate( .a(N43), .b(D_244_NOT), .O(ED_1220) );
and2 gate( .a(N43_NOT), .b(D_244_NOT), .O(ED_1221) );
and2 gate( .a(CONST1), .b(D_244), .O(ED_1222) );
and2 gate( .a(CONST0), .b(D_244), .O(ED_1223) );
and2 gate( .a(ED_1220), .b(D_245_NOT), .O(ED_1229) );
and2 gate( .a(ED_1221), .b(D_245), .O(ED_1227) );
and2 gate( .a(ED_1222), .b(D_245_NOT), .O(ED_1225) );
and2 gate( .a(ED_1223), .b(D_245), .O(ED_1224) );
or2  gate( .a(ED_1224), .b(ED_1225), .O(ED_1226) );
or2  gate( .a(ED_1226), .b(ED_1227), .O(ED_1228) );
or2  gate( .a(ED_1229), .b(ED_1228), .O(N43_OBF) );
inv1 gate( .a(D_246), .O(D_246_NOT) );
inv1 gate( .a(D_247), .O(D_247_NOT) );
inv1 gate( .a(N24), .O(N24_NOT) );
and2 gate( .a(N24), .b(D_246_NOT), .O(ED_1230) );
and2 gate( .a(N24_NOT), .b(D_246_NOT), .O(ED_1231) );
and2 gate( .a(CONST1), .b(D_246), .O(ED_1232) );
and2 gate( .a(CONST0), .b(D_246), .O(ED_1233) );
and2 gate( .a(ED_1230), .b(D_247_NOT), .O(ED_1239) );
and2 gate( .a(ED_1231), .b(D_247), .O(ED_1237) );
and2 gate( .a(ED_1232), .b(D_247_NOT), .O(ED_1235) );
and2 gate( .a(ED_1233), .b(D_247), .O(ED_1234) );
or2  gate( .a(ED_1234), .b(ED_1235), .O(ED_1236) );
or2  gate( .a(ED_1236), .b(ED_1237), .O(ED_1238) );
or2  gate( .a(ED_1239), .b(ED_1238), .O(N24_OBF) );
inv1 gate( .a(D_248), .O(D_248_NOT) );
inv1 gate( .a(D_249), .O(D_249_NOT) );
inv1 gate( .a(N259), .O(N259_NOT) );
and2 gate( .a(N259), .b(D_248_NOT), .O(ED_1240) );
and2 gate( .a(N259_NOT), .b(D_248_NOT), .O(ED_1241) );
and2 gate( .a(CONST1), .b(D_248), .O(ED_1242) );
and2 gate( .a(CONST0), .b(D_248), .O(ED_1243) );
and2 gate( .a(ED_1240), .b(D_249_NOT), .O(ED_1249) );
and2 gate( .a(ED_1241), .b(D_249), .O(ED_1247) );
and2 gate( .a(ED_1242), .b(D_249_NOT), .O(ED_1245) );
and2 gate( .a(ED_1243), .b(D_249), .O(ED_1244) );
or2  gate( .a(ED_1244), .b(ED_1245), .O(ED_1246) );
or2  gate( .a(ED_1246), .b(ED_1247), .O(ED_1248) );
or2  gate( .a(ED_1249), .b(ED_1248), .O(N259_OBF) );
inv1 gate( .a(D_250), .O(D_250_NOT) );
inv1 gate( .a(D_251), .O(D_251_NOT) );
inv1 gate( .a(N319), .O(N319_NOT) );
and2 gate( .a(N319), .b(D_250_NOT), .O(ED_1250) );
and2 gate( .a(N319_NOT), .b(D_250_NOT), .O(ED_1251) );
and2 gate( .a(CONST1), .b(D_250), .O(ED_1252) );
and2 gate( .a(CONST0), .b(D_250), .O(ED_1253) );
and2 gate( .a(ED_1250), .b(D_251_NOT), .O(ED_1259) );
and2 gate( .a(ED_1251), .b(D_251), .O(ED_1257) );
and2 gate( .a(ED_1252), .b(D_251_NOT), .O(ED_1255) );
and2 gate( .a(ED_1253), .b(D_251), .O(ED_1254) );
or2  gate( .a(ED_1254), .b(ED_1255), .O(ED_1256) );
or2  gate( .a(ED_1256), .b(ED_1257), .O(ED_1258) );
or2  gate( .a(ED_1259), .b(ED_1258), .O(N319_OBF) );
inv1 gate( .a(D_252), .O(D_252_NOT) );
inv1 gate( .a(D_253), .O(D_253_NOT) );
inv1 gate( .a(N105), .O(N105_NOT) );
and2 gate( .a(N105), .b(D_252_NOT), .O(ED_1260) );
and2 gate( .a(N105_NOT), .b(D_252_NOT), .O(ED_1261) );
and2 gate( .a(CONST1), .b(D_252), .O(ED_1262) );
and2 gate( .a(CONST0), .b(D_252), .O(ED_1263) );
and2 gate( .a(ED_1260), .b(D_253_NOT), .O(ED_1269) );
and2 gate( .a(ED_1261), .b(D_253), .O(ED_1267) );
and2 gate( .a(ED_1262), .b(D_253_NOT), .O(ED_1265) );
and2 gate( .a(ED_1263), .b(D_253), .O(ED_1264) );
or2  gate( .a(ED_1264), .b(ED_1265), .O(ED_1266) );
or2  gate( .a(ED_1266), .b(ED_1267), .O(ED_1268) );
or2  gate( .a(ED_1269), .b(ED_1268), .O(N105_OBF) );
inv1 gate( .a(D_254), .O(D_254_NOT) );
inv1 gate( .a(D_255), .O(D_255_NOT) );
inv1 gate( .a(N343), .O(N343_NOT) );
and2 gate( .a(N343), .b(D_254_NOT), .O(ED_1270) );
and2 gate( .a(N343_NOT), .b(D_254_NOT), .O(ED_1271) );
and2 gate( .a(CONST1), .b(D_254), .O(ED_1272) );
and2 gate( .a(CONST0), .b(D_254), .O(ED_1273) );
and2 gate( .a(ED_1270), .b(D_255_NOT), .O(ED_1279) );
and2 gate( .a(ED_1271), .b(D_255), .O(ED_1277) );
and2 gate( .a(ED_1272), .b(D_255_NOT), .O(ED_1275) );
and2 gate( .a(ED_1273), .b(D_255), .O(ED_1274) );
or2  gate( .a(ED_1274), .b(ED_1275), .O(ED_1276) );
or2  gate( .a(ED_1276), .b(ED_1277), .O(ED_1278) );
or2  gate( .a(ED_1279), .b(ED_1278), .O(N343_OBF) );
inv1 gate( .a(D_256), .O(D_256_NOT) );
inv1 gate( .a(D_257), .O(D_257_NOT) );
inv1 gate( .a(N89), .O(N89_NOT) );
and2 gate( .a(N89), .b(D_256_NOT), .O(ED_1280) );
and2 gate( .a(N89_NOT), .b(D_256_NOT), .O(ED_1281) );
and2 gate( .a(CONST1), .b(D_256), .O(ED_1282) );
and2 gate( .a(CONST0), .b(D_256), .O(ED_1283) );
and2 gate( .a(ED_1280), .b(D_257_NOT), .O(ED_1289) );
and2 gate( .a(ED_1281), .b(D_257), .O(ED_1287) );
and2 gate( .a(ED_1282), .b(D_257_NOT), .O(ED_1285) );
and2 gate( .a(ED_1283), .b(D_257), .O(ED_1284) );
or2  gate( .a(ED_1284), .b(ED_1285), .O(ED_1286) );
or2  gate( .a(ED_1286), .b(ED_1287), .O(ED_1288) );
or2  gate( .a(ED_1289), .b(ED_1288), .O(N89_OBF) );
inv1 gate( .a(D_258), .O(D_258_NOT) );
inv1 gate( .a(D_259), .O(D_259_NOT) );
inv1 gate( .a(N380), .O(N380_NOT) );
and2 gate( .a(N380), .b(D_258_NOT), .O(ED_1290) );
and2 gate( .a(N380_NOT), .b(D_258_NOT), .O(ED_1291) );
and2 gate( .a(CONST1), .b(D_258), .O(ED_1292) );
and2 gate( .a(CONST0), .b(D_258), .O(ED_1293) );
and2 gate( .a(ED_1290), .b(D_259_NOT), .O(ED_1299) );
and2 gate( .a(ED_1291), .b(D_259), .O(ED_1297) );
and2 gate( .a(ED_1292), .b(D_259_NOT), .O(ED_1295) );
and2 gate( .a(ED_1293), .b(D_259), .O(ED_1294) );
or2  gate( .a(ED_1294), .b(ED_1295), .O(ED_1296) );
or2  gate( .a(ED_1296), .b(ED_1297), .O(ED_1298) );
or2  gate( .a(ED_1299), .b(ED_1298), .O(N380_OBF) );
inv1 gate( .a(D_260), .O(D_260_NOT) );
inv1 gate( .a(D_261), .O(D_261_NOT) );
inv1 gate( .a(N224), .O(N224_NOT) );
and2 gate( .a(N224), .b(D_260_NOT), .O(ED_1300) );
and2 gate( .a(N224_NOT), .b(D_260_NOT), .O(ED_1301) );
and2 gate( .a(CONST1), .b(D_260), .O(ED_1302) );
and2 gate( .a(CONST0), .b(D_260), .O(ED_1303) );
and2 gate( .a(ED_1300), .b(D_261_NOT), .O(ED_1309) );
and2 gate( .a(ED_1301), .b(D_261), .O(ED_1307) );
and2 gate( .a(ED_1302), .b(D_261_NOT), .O(ED_1305) );
and2 gate( .a(ED_1303), .b(D_261), .O(ED_1304) );
or2  gate( .a(ED_1304), .b(ED_1305), .O(ED_1306) );
or2  gate( .a(ED_1306), .b(ED_1307), .O(ED_1308) );
or2  gate( .a(ED_1309), .b(ED_1308), .O(N224_OBF) );
inv1 gate( .a(D_262), .O(D_262_NOT) );
inv1 gate( .a(D_263), .O(D_263_NOT) );
inv1 gate( .a(N255), .O(N255_NOT) );
and2 gate( .a(N255), .b(D_262_NOT), .O(ED_1310) );
and2 gate( .a(N255_NOT), .b(D_262_NOT), .O(ED_1311) );
and2 gate( .a(CONST1), .b(D_262), .O(ED_1312) );
and2 gate( .a(CONST0), .b(D_262), .O(ED_1313) );
and2 gate( .a(ED_1310), .b(D_263_NOT), .O(ED_1319) );
and2 gate( .a(ED_1311), .b(D_263), .O(ED_1317) );
and2 gate( .a(ED_1312), .b(D_263_NOT), .O(ED_1315) );
and2 gate( .a(ED_1313), .b(D_263), .O(ED_1314) );
or2  gate( .a(ED_1314), .b(ED_1315), .O(ED_1316) );
or2  gate( .a(ED_1316), .b(ED_1317), .O(ED_1318) );
or2  gate( .a(ED_1319), .b(ED_1318), .O(N255_OBF) );
inv1 gate( .a(D_264), .O(D_264_NOT) );
inv1 gate( .a(D_265), .O(D_265_NOT) );
inv1 gate( .a(N198), .O(N198_NOT) );
and2 gate( .a(N198), .b(D_264_NOT), .O(ED_1320) );
and2 gate( .a(N198_NOT), .b(D_264_NOT), .O(ED_1321) );
and2 gate( .a(CONST1), .b(D_264), .O(ED_1322) );
and2 gate( .a(CONST0), .b(D_264), .O(ED_1323) );
and2 gate( .a(ED_1320), .b(D_265_NOT), .O(ED_1329) );
and2 gate( .a(ED_1321), .b(D_265), .O(ED_1327) );
and2 gate( .a(ED_1322), .b(D_265_NOT), .O(ED_1325) );
and2 gate( .a(ED_1323), .b(D_265), .O(ED_1324) );
or2  gate( .a(ED_1324), .b(ED_1325), .O(ED_1326) );
or2  gate( .a(ED_1326), .b(ED_1327), .O(ED_1328) );
or2  gate( .a(ED_1329), .b(ED_1328), .O(N198_OBF) );
inv1 gate( .a(D_266), .O(D_266_NOT) );
inv1 gate( .a(D_267), .O(D_267_NOT) );
inv1 gate( .a(N34), .O(N34_NOT) );
and2 gate( .a(N34), .b(D_266_NOT), .O(ED_1330) );
and2 gate( .a(N34_NOT), .b(D_266_NOT), .O(ED_1331) );
and2 gate( .a(CONST1), .b(D_266), .O(ED_1332) );
and2 gate( .a(CONST0), .b(D_266), .O(ED_1333) );
and2 gate( .a(ED_1330), .b(D_267_NOT), .O(ED_1339) );
and2 gate( .a(ED_1331), .b(D_267), .O(ED_1337) );
and2 gate( .a(ED_1332), .b(D_267_NOT), .O(ED_1335) );
and2 gate( .a(ED_1333), .b(D_267), .O(ED_1334) );
or2  gate( .a(ED_1334), .b(ED_1335), .O(ED_1336) );
or2  gate( .a(ED_1336), .b(ED_1337), .O(ED_1338) );
or2  gate( .a(ED_1339), .b(ED_1338), .O(N34_OBF) );
inv1 gate( .a(D_268), .O(D_268_NOT) );
inv1 gate( .a(D_269), .O(D_269_NOT) );
inv1 gate( .a(N337), .O(N337_NOT) );
and2 gate( .a(N337), .b(D_268_NOT), .O(ED_1340) );
and2 gate( .a(N337_NOT), .b(D_268_NOT), .O(ED_1341) );
and2 gate( .a(CONST1), .b(D_268), .O(ED_1342) );
and2 gate( .a(CONST0), .b(D_268), .O(ED_1343) );
and2 gate( .a(ED_1340), .b(D_269_NOT), .O(ED_1349) );
and2 gate( .a(ED_1341), .b(D_269), .O(ED_1347) );
and2 gate( .a(ED_1342), .b(D_269_NOT), .O(ED_1345) );
and2 gate( .a(ED_1343), .b(D_269), .O(ED_1344) );
or2  gate( .a(ED_1344), .b(ED_1345), .O(ED_1346) );
or2  gate( .a(ED_1346), .b(ED_1347), .O(ED_1348) );
or2  gate( .a(ED_1349), .b(ED_1348), .O(N337_OBF) );
inv1 gate( .a(D_270), .O(D_270_NOT) );
inv1 gate( .a(D_271), .O(D_271_NOT) );
inv1 gate( .a(N142), .O(N142_NOT) );
and2 gate( .a(N142), .b(D_270_NOT), .O(ED_1350) );
and2 gate( .a(N142_NOT), .b(D_270_NOT), .O(ED_1351) );
and2 gate( .a(CONST1), .b(D_270), .O(ED_1352) );
and2 gate( .a(CONST0), .b(D_270), .O(ED_1353) );
and2 gate( .a(ED_1350), .b(D_271_NOT), .O(ED_1359) );
and2 gate( .a(ED_1351), .b(D_271), .O(ED_1357) );
and2 gate( .a(ED_1352), .b(D_271_NOT), .O(ED_1355) );
and2 gate( .a(ED_1353), .b(D_271), .O(ED_1354) );
or2  gate( .a(ED_1354), .b(ED_1355), .O(ED_1356) );
or2  gate( .a(ED_1356), .b(ED_1357), .O(ED_1358) );
or2  gate( .a(ED_1359), .b(ED_1358), .O(N142_OBF) );
inv1 gate( .a(D_272), .O(D_272_NOT) );
inv1 gate( .a(D_273), .O(D_273_NOT) );
inv1 gate( .a(N393), .O(N393_NOT) );
and2 gate( .a(N393), .b(D_272_NOT), .O(ED_1360) );
and2 gate( .a(N393_NOT), .b(D_272_NOT), .O(ED_1361) );
and2 gate( .a(CONST1), .b(D_272), .O(ED_1362) );
and2 gate( .a(CONST0), .b(D_272), .O(ED_1363) );
and2 gate( .a(ED_1360), .b(D_273_NOT), .O(ED_1369) );
and2 gate( .a(ED_1361), .b(D_273), .O(ED_1367) );
and2 gate( .a(ED_1362), .b(D_273_NOT), .O(ED_1365) );
and2 gate( .a(ED_1363), .b(D_273), .O(ED_1364) );
or2  gate( .a(ED_1364), .b(ED_1365), .O(ED_1366) );
or2  gate( .a(ED_1366), .b(ED_1367), .O(ED_1368) );
or2  gate( .a(ED_1369), .b(ED_1368), .O(N393_OBF) );
inv1 gate( .a(D_274), .O(D_274_NOT) );
inv1 gate( .a(D_275), .O(D_275_NOT) );
inv1 gate( .a(N82), .O(N82_NOT) );
and2 gate( .a(N82), .b(D_274_NOT), .O(ED_1370) );
and2 gate( .a(N82_NOT), .b(D_274_NOT), .O(ED_1371) );
and2 gate( .a(CONST1), .b(D_274), .O(ED_1372) );
and2 gate( .a(CONST0), .b(D_274), .O(ED_1373) );
and2 gate( .a(ED_1370), .b(D_275_NOT), .O(ED_1379) );
and2 gate( .a(ED_1371), .b(D_275), .O(ED_1377) );
and2 gate( .a(ED_1372), .b(D_275_NOT), .O(ED_1375) );
and2 gate( .a(ED_1373), .b(D_275), .O(ED_1374) );
or2  gate( .a(ED_1374), .b(ED_1375), .O(ED_1376) );
or2  gate( .a(ED_1376), .b(ED_1377), .O(ED_1378) );
or2  gate( .a(ED_1379), .b(ED_1378), .O(N82_OBF) );
inv1 gate( .a(D_276), .O(D_276_NOT) );
inv1 gate( .a(D_277), .O(D_277_NOT) );
inv1 gate( .a(N319), .O(N319_NOT) );
and2 gate( .a(N319), .b(D_276_NOT), .O(ED_1380) );
and2 gate( .a(N319_NOT), .b(D_276_NOT), .O(ED_1381) );
and2 gate( .a(CONST1), .b(D_276), .O(ED_1382) );
and2 gate( .a(CONST0), .b(D_276), .O(ED_1383) );
and2 gate( .a(ED_1380), .b(D_277_NOT), .O(ED_1389) );
and2 gate( .a(ED_1381), .b(D_277), .O(ED_1387) );
and2 gate( .a(ED_1382), .b(D_277_NOT), .O(ED_1385) );
and2 gate( .a(ED_1383), .b(D_277), .O(ED_1384) );
or2  gate( .a(ED_1384), .b(ED_1385), .O(ED_1386) );
or2  gate( .a(ED_1386), .b(ED_1387), .O(ED_1388) );
or2  gate( .a(ED_1389), .b(ED_1388), .O(N319_OBF) );
inv1 gate( .a(D_278), .O(D_278_NOT) );
inv1 gate( .a(D_279), .O(D_279_NOT) );
inv1 gate( .a(N30), .O(N30_NOT) );
and2 gate( .a(N30), .b(D_278_NOT), .O(ED_1390) );
and2 gate( .a(N30_NOT), .b(D_278_NOT), .O(ED_1391) );
and2 gate( .a(CONST1), .b(D_278), .O(ED_1392) );
and2 gate( .a(CONST0), .b(D_278), .O(ED_1393) );
and2 gate( .a(ED_1390), .b(D_279_NOT), .O(ED_1399) );
and2 gate( .a(ED_1391), .b(D_279), .O(ED_1397) );
and2 gate( .a(ED_1392), .b(D_279_NOT), .O(ED_1395) );
and2 gate( .a(ED_1393), .b(D_279), .O(ED_1394) );
or2  gate( .a(ED_1394), .b(ED_1395), .O(ED_1396) );
or2  gate( .a(ED_1396), .b(ED_1397), .O(ED_1398) );
or2  gate( .a(ED_1399), .b(ED_1398), .O(N30_OBF) );
inv1 gate( .a(D_280), .O(D_280_NOT) );
inv1 gate( .a(D_281), .O(D_281_NOT) );
inv1 gate( .a(N357), .O(N357_NOT) );
and2 gate( .a(N357), .b(D_280_NOT), .O(ED_1400) );
and2 gate( .a(N357_NOT), .b(D_280_NOT), .O(ED_1401) );
and2 gate( .a(CONST1), .b(D_280), .O(ED_1402) );
and2 gate( .a(CONST0), .b(D_280), .O(ED_1403) );
and2 gate( .a(ED_1400), .b(D_281_NOT), .O(ED_1409) );
and2 gate( .a(ED_1401), .b(D_281), .O(ED_1407) );
and2 gate( .a(ED_1402), .b(D_281_NOT), .O(ED_1405) );
and2 gate( .a(ED_1403), .b(D_281), .O(ED_1404) );
or2  gate( .a(ED_1404), .b(ED_1405), .O(ED_1406) );
or2  gate( .a(ED_1406), .b(ED_1407), .O(ED_1408) );
or2  gate( .a(ED_1409), .b(ED_1408), .O(N357_OBF) );
inv1 gate( .a(D_282), .O(D_282_NOT) );
inv1 gate( .a(D_283), .O(D_283_NOT) );
inv1 gate( .a(N126), .O(N126_NOT) );
and2 gate( .a(N126), .b(D_282_NOT), .O(ED_1410) );
and2 gate( .a(N126_NOT), .b(D_282_NOT), .O(ED_1411) );
and2 gate( .a(CONST1), .b(D_282), .O(ED_1412) );
and2 gate( .a(CONST0), .b(D_282), .O(ED_1413) );
and2 gate( .a(ED_1410), .b(D_283_NOT), .O(ED_1419) );
and2 gate( .a(ED_1411), .b(D_283), .O(ED_1417) );
and2 gate( .a(ED_1412), .b(D_283_NOT), .O(ED_1415) );
and2 gate( .a(ED_1413), .b(D_283), .O(ED_1414) );
or2  gate( .a(ED_1414), .b(ED_1415), .O(ED_1416) );
or2  gate( .a(ED_1416), .b(ED_1417), .O(ED_1418) );
or2  gate( .a(ED_1419), .b(ED_1418), .O(N126_OBF) );

endmodule
