module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate581(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate582(.a(gate19inter0), .b(s_60), .O(gate19inter1));
  and2  gate583(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate584(.a(s_60), .O(gate19inter3));
  inv1  gate585(.a(s_61), .O(gate19inter4));
  nand2 gate586(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate587(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate588(.a(N118), .O(gate19inter7));
  inv1  gate589(.a(N4), .O(gate19inter8));
  nand2 gate590(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate591(.a(s_61), .b(gate19inter3), .O(gate19inter10));
  nor2  gate592(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate593(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate594(.a(gate19inter12), .b(gate19inter1), .O(N154));
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );

  xor2  gate413(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate414(.a(gate25inter0), .b(s_36), .O(gate25inter1));
  and2  gate415(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate416(.a(s_36), .O(gate25inter3));
  inv1  gate417(.a(s_37), .O(gate25inter4));
  nand2 gate418(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate419(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate420(.a(N134), .O(gate25inter7));
  inv1  gate421(.a(N56), .O(gate25inter8));
  nand2 gate422(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate423(.a(s_37), .b(gate25inter3), .O(gate25inter10));
  nor2  gate424(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate425(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate426(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate231(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate232(.a(gate29inter0), .b(s_10), .O(gate29inter1));
  and2  gate233(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate234(.a(s_10), .O(gate29inter3));
  inv1  gate235(.a(s_11), .O(gate29inter4));
  nand2 gate236(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate237(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate238(.a(N150), .O(gate29inter7));
  inv1  gate239(.a(N108), .O(gate29inter8));
  nand2 gate240(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate241(.a(s_11), .b(gate29inter3), .O(gate29inter10));
  nor2  gate242(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate243(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate244(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate371(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate372(.a(gate32inter0), .b(s_30), .O(gate32inter1));
  and2  gate373(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate374(.a(s_30), .O(gate32inter3));
  inv1  gate375(.a(s_31), .O(gate32inter4));
  nand2 gate376(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate377(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate378(.a(N34), .O(gate32inter7));
  inv1  gate379(.a(N127), .O(gate32inter8));
  nand2 gate380(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate381(.a(s_31), .b(gate32inter3), .O(gate32inter10));
  nor2  gate382(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate383(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate384(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate441(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate442(.a(gate34inter0), .b(s_40), .O(gate34inter1));
  and2  gate443(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate444(.a(s_40), .O(gate34inter3));
  inv1  gate445(.a(s_41), .O(gate34inter4));
  nand2 gate446(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate447(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate448(.a(N47), .O(gate34inter7));
  inv1  gate449(.a(N131), .O(gate34inter8));
  nand2 gate450(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate451(.a(s_41), .b(gate34inter3), .O(gate34inter10));
  nor2  gate452(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate453(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate454(.a(gate34inter12), .b(gate34inter1), .O(N187));
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate651(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate652(.a(gate37inter0), .b(s_70), .O(gate37inter1));
  and2  gate653(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate654(.a(s_70), .O(gate37inter3));
  inv1  gate655(.a(s_71), .O(gate37inter4));
  nand2 gate656(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate657(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate658(.a(N66), .O(gate37inter7));
  inv1  gate659(.a(N135), .O(gate37inter8));
  nand2 gate660(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate661(.a(s_71), .b(gate37inter3), .O(gate37inter10));
  nor2  gate662(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate663(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate664(.a(gate37inter12), .b(gate37inter1), .O(N190));

  xor2  gate385(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate386(.a(gate38inter0), .b(s_32), .O(gate38inter1));
  and2  gate387(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate388(.a(s_32), .O(gate38inter3));
  inv1  gate389(.a(s_33), .O(gate38inter4));
  nand2 gate390(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate391(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate392(.a(N73), .O(gate38inter7));
  inv1  gate393(.a(N139), .O(gate38inter8));
  nand2 gate394(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate395(.a(s_33), .b(gate38inter3), .O(gate38inter10));
  nor2  gate396(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate397(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate398(.a(gate38inter12), .b(gate38inter1), .O(N191));
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate259(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate260(.a(gate41inter0), .b(s_14), .O(gate41inter1));
  and2  gate261(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate262(.a(s_14), .O(gate41inter3));
  inv1  gate263(.a(s_15), .O(gate41inter4));
  nand2 gate264(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate265(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate266(.a(N92), .O(gate41inter7));
  inv1  gate267(.a(N143), .O(gate41inter8));
  nand2 gate268(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate269(.a(s_15), .b(gate41inter3), .O(gate41inter10));
  nor2  gate270(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate271(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate272(.a(gate41inter12), .b(gate41inter1), .O(N194));

  xor2  gate553(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate554(.a(gate42inter0), .b(s_56), .O(gate42inter1));
  and2  gate555(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate556(.a(s_56), .O(gate42inter3));
  inv1  gate557(.a(s_57), .O(gate42inter4));
  nand2 gate558(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate559(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate560(.a(N99), .O(gate42inter7));
  inv1  gate561(.a(N147), .O(gate42inter8));
  nand2 gate562(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate563(.a(s_57), .b(gate42inter3), .O(gate42inter10));
  nor2  gate564(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate565(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate566(.a(gate42inter12), .b(gate42inter1), .O(N195));

  xor2  gate287(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate288(.a(gate43inter0), .b(s_18), .O(gate43inter1));
  and2  gate289(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate290(.a(s_18), .O(gate43inter3));
  inv1  gate291(.a(s_19), .O(gate43inter4));
  nand2 gate292(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate293(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate294(.a(N105), .O(gate43inter7));
  inv1  gate295(.a(N147), .O(gate43inter8));
  nand2 gate296(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate297(.a(s_19), .b(gate43inter3), .O(gate43inter10));
  nor2  gate298(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate299(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate300(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );

  xor2  gate539(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate540(.a(gate45inter0), .b(s_54), .O(gate45inter1));
  and2  gate541(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate542(.a(s_54), .O(gate45inter3));
  inv1  gate543(.a(s_55), .O(gate45inter4));
  nand2 gate544(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate545(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate546(.a(N115), .O(gate45inter7));
  inv1  gate547(.a(N151), .O(gate45inter8));
  nand2 gate548(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate549(.a(s_55), .b(gate45inter3), .O(gate45inter10));
  nor2  gate550(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate551(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate552(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );

  xor2  gate315(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate316(.a(gate55inter0), .b(s_22), .O(gate55inter1));
  and2  gate317(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate318(.a(s_22), .O(gate55inter3));
  inv1  gate319(.a(s_23), .O(gate55inter4));
  nand2 gate320(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate321(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate322(.a(N203), .O(gate55inter7));
  inv1  gate323(.a(N171), .O(gate55inter8));
  nand2 gate324(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate325(.a(s_23), .b(gate55inter3), .O(gate55inter10));
  nor2  gate326(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate327(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate328(.a(gate55inter12), .b(gate55inter1), .O(N239));
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate189(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate190(.a(gate62inter0), .b(s_4), .O(gate62inter1));
  and2  gate191(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate192(.a(s_4), .O(gate62inter3));
  inv1  gate193(.a(s_5), .O(gate62inter4));
  nand2 gate194(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate195(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate196(.a(N213), .O(gate62inter7));
  inv1  gate197(.a(N37), .O(gate62inter8));
  nand2 gate198(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate199(.a(s_5), .b(gate62inter3), .O(gate62inter10));
  nor2  gate200(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate201(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate202(.a(gate62inter12), .b(gate62inter1), .O(N254));
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );

  xor2  gate301(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate302(.a(gate66inter0), .b(s_20), .O(gate66inter1));
  and2  gate303(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate304(.a(s_20), .O(gate66inter3));
  inv1  gate305(.a(s_21), .O(gate66inter4));
  nand2 gate306(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate307(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate308(.a(N213), .O(gate66inter7));
  inv1  gate309(.a(N89), .O(gate66inter8));
  nand2 gate310(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate311(.a(s_21), .b(gate66inter3), .O(gate66inter10));
  nor2  gate312(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate313(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate314(.a(gate66inter12), .b(gate66inter1), .O(N258));
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );

  xor2  gate595(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate596(.a(gate74inter0), .b(s_62), .O(gate74inter1));
  and2  gate597(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate598(.a(s_62), .O(gate74inter3));
  inv1  gate599(.a(s_63), .O(gate74inter4));
  nand2 gate600(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate601(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate602(.a(N239), .O(gate74inter7));
  inv1  gate603(.a(N191), .O(gate74inter8));
  nand2 gate604(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate605(.a(s_63), .b(gate74inter3), .O(gate74inter10));
  nor2  gate606(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate607(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate608(.a(gate74inter12), .b(gate74inter1), .O(N276));

  xor2  gate693(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate694(.a(gate75inter0), .b(s_76), .O(gate75inter1));
  and2  gate695(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate696(.a(s_76), .O(gate75inter3));
  inv1  gate697(.a(s_77), .O(gate75inter4));
  nand2 gate698(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate699(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate700(.a(N243), .O(gate75inter7));
  inv1  gate701(.a(N193), .O(gate75inter8));
  nand2 gate702(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate703(.a(s_77), .b(gate75inter3), .O(gate75inter10));
  nor2  gate704(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate705(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate706(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate483(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate484(.a(gate77inter0), .b(s_46), .O(gate77inter1));
  and2  gate485(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate486(.a(s_46), .O(gate77inter3));
  inv1  gate487(.a(s_47), .O(gate77inter4));
  nand2 gate488(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate489(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate490(.a(N251), .O(gate77inter7));
  inv1  gate491(.a(N197), .O(gate77inter8));
  nand2 gate492(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate493(.a(s_47), .b(gate77inter3), .O(gate77inter10));
  nor2  gate494(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate495(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate496(.a(gate77inter12), .b(gate77inter1), .O(N285));

  xor2  gate791(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate792(.a(gate78inter0), .b(s_90), .O(gate78inter1));
  and2  gate793(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate794(.a(s_90), .O(gate78inter3));
  inv1  gate795(.a(s_91), .O(gate78inter4));
  nand2 gate796(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate797(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate798(.a(N227), .O(gate78inter7));
  inv1  gate799(.a(N184), .O(gate78inter8));
  nand2 gate800(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate801(.a(s_91), .b(gate78inter3), .O(gate78inter10));
  nor2  gate802(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate803(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate804(.a(gate78inter12), .b(gate78inter1), .O(N288));

  xor2  gate203(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate204(.a(gate79inter0), .b(s_6), .O(gate79inter1));
  and2  gate205(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate206(.a(s_6), .O(gate79inter3));
  inv1  gate207(.a(s_7), .O(gate79inter4));
  nand2 gate208(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate209(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate210(.a(N230), .O(gate79inter7));
  inv1  gate211(.a(N186), .O(gate79inter8));
  nand2 gate212(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate213(.a(s_7), .b(gate79inter3), .O(gate79inter10));
  nor2  gate214(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate215(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate216(.a(gate79inter12), .b(gate79inter1), .O(N289));

  xor2  gate455(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate456(.a(gate80inter0), .b(s_42), .O(gate80inter1));
  and2  gate457(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate458(.a(s_42), .O(gate80inter3));
  inv1  gate459(.a(s_43), .O(gate80inter4));
  nand2 gate460(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate461(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate462(.a(N233), .O(gate80inter7));
  inv1  gate463(.a(N188), .O(gate80inter8));
  nand2 gate464(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate465(.a(s_43), .b(gate80inter3), .O(gate80inter10));
  nor2  gate466(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate467(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate468(.a(gate80inter12), .b(gate80inter1), .O(N290));

  xor2  gate749(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate750(.a(gate81inter0), .b(s_84), .O(gate81inter1));
  and2  gate751(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate752(.a(s_84), .O(gate81inter3));
  inv1  gate753(.a(s_85), .O(gate81inter4));
  nand2 gate754(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate755(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate756(.a(N236), .O(gate81inter7));
  inv1  gate757(.a(N190), .O(gate81inter8));
  nand2 gate758(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate759(.a(s_85), .b(gate81inter3), .O(gate81inter10));
  nor2  gate760(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate761(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate762(.a(gate81inter12), .b(gate81inter1), .O(N291));

  xor2  gate511(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate512(.a(gate82inter0), .b(s_50), .O(gate82inter1));
  and2  gate513(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate514(.a(s_50), .O(gate82inter3));
  inv1  gate515(.a(s_51), .O(gate82inter4));
  nand2 gate516(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate517(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate518(.a(N239), .O(gate82inter7));
  inv1  gate519(.a(N192), .O(gate82inter8));
  nand2 gate520(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate521(.a(s_51), .b(gate82inter3), .O(gate82inter10));
  nor2  gate522(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate523(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate524(.a(gate82inter12), .b(gate82inter1), .O(N292));

  xor2  gate735(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate736(.a(gate83inter0), .b(s_82), .O(gate83inter1));
  and2  gate737(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate738(.a(s_82), .O(gate83inter3));
  inv1  gate739(.a(s_83), .O(gate83inter4));
  nand2 gate740(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate741(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate742(.a(N243), .O(gate83inter7));
  inv1  gate743(.a(N194), .O(gate83inter8));
  nand2 gate744(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate745(.a(s_83), .b(gate83inter3), .O(gate83inter10));
  nor2  gate746(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate747(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate748(.a(gate83inter12), .b(gate83inter1), .O(N293));

  xor2  gate357(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate358(.a(gate84inter0), .b(s_28), .O(gate84inter1));
  and2  gate359(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate360(.a(s_28), .O(gate84inter3));
  inv1  gate361(.a(s_29), .O(gate84inter4));
  nand2 gate362(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate363(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate364(.a(N247), .O(gate84inter7));
  inv1  gate365(.a(N196), .O(gate84inter8));
  nand2 gate366(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate367(.a(s_29), .b(gate84inter3), .O(gate84inter10));
  nor2  gate368(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate369(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate370(.a(gate84inter12), .b(gate84inter1), .O(N294));

  xor2  gate777(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate778(.a(gate85inter0), .b(s_88), .O(gate85inter1));
  and2  gate779(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate780(.a(s_88), .O(gate85inter3));
  inv1  gate781(.a(s_89), .O(gate85inter4));
  nand2 gate782(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate783(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate784(.a(N251), .O(gate85inter7));
  inv1  gate785(.a(N198), .O(gate85inter8));
  nand2 gate786(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate787(.a(s_89), .b(gate85inter3), .O(gate85inter10));
  nor2  gate788(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate789(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate790(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate161(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate162(.a(gate99inter0), .b(s_0), .O(gate99inter1));
  and2  gate163(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate164(.a(s_0), .O(gate99inter3));
  inv1  gate165(.a(s_1), .O(gate99inter4));
  nand2 gate166(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate167(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate168(.a(N309), .O(gate99inter7));
  inv1  gate169(.a(N260), .O(gate99inter8));
  nand2 gate170(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate171(.a(s_1), .b(gate99inter3), .O(gate99inter10));
  nor2  gate172(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate173(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate174(.a(gate99inter12), .b(gate99inter1), .O(N330));

  xor2  gate427(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate428(.a(gate100inter0), .b(s_38), .O(gate100inter1));
  and2  gate429(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate430(.a(s_38), .O(gate100inter3));
  inv1  gate431(.a(s_39), .O(gate100inter4));
  nand2 gate432(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate433(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate434(.a(N309), .O(gate100inter7));
  inv1  gate435(.a(N264), .O(gate100inter8));
  nand2 gate436(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate437(.a(s_39), .b(gate100inter3), .O(gate100inter10));
  nor2  gate438(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate439(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate440(.a(gate100inter12), .b(gate100inter1), .O(N331));

  xor2  gate245(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate246(.a(gate101inter0), .b(s_12), .O(gate101inter1));
  and2  gate247(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate248(.a(s_12), .O(gate101inter3));
  inv1  gate249(.a(s_13), .O(gate101inter4));
  nand2 gate250(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate251(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate252(.a(N309), .O(gate101inter7));
  inv1  gate253(.a(N267), .O(gate101inter8));
  nand2 gate254(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate255(.a(s_13), .b(gate101inter3), .O(gate101inter10));
  nor2  gate256(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate257(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate258(.a(gate101inter12), .b(gate101inter1), .O(N332));
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate665(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate666(.a(gate103inter0), .b(s_72), .O(gate103inter1));
  and2  gate667(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate668(.a(s_72), .O(gate103inter3));
  inv1  gate669(.a(s_73), .O(gate103inter4));
  nand2 gate670(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate671(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate672(.a(N8), .O(gate103inter7));
  inv1  gate673(.a(N319), .O(gate103inter8));
  nand2 gate674(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate675(.a(s_73), .b(gate103inter3), .O(gate103inter10));
  nor2  gate676(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate677(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate678(.a(gate103inter12), .b(gate103inter1), .O(N334));

  xor2  gate679(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate680(.a(gate104inter0), .b(s_74), .O(gate104inter1));
  and2  gate681(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate682(.a(s_74), .O(gate104inter3));
  inv1  gate683(.a(s_75), .O(gate104inter4));
  nand2 gate684(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate685(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate686(.a(N309), .O(gate104inter7));
  inv1  gate687(.a(N273), .O(gate104inter8));
  nand2 gate688(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate689(.a(s_75), .b(gate104inter3), .O(gate104inter10));
  nor2  gate690(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate691(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate692(.a(gate104inter12), .b(gate104inter1), .O(N335));

  xor2  gate399(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate400(.a(gate105inter0), .b(s_34), .O(gate105inter1));
  and2  gate401(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate402(.a(s_34), .O(gate105inter3));
  inv1  gate403(.a(s_35), .O(gate105inter4));
  nand2 gate404(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate405(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate406(.a(N319), .O(gate105inter7));
  inv1  gate407(.a(N21), .O(gate105inter8));
  nand2 gate408(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate409(.a(s_35), .b(gate105inter3), .O(gate105inter10));
  nor2  gate410(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate411(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate412(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );

  xor2  gate609(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate610(.a(gate107inter0), .b(s_64), .O(gate107inter1));
  and2  gate611(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate612(.a(s_64), .O(gate107inter3));
  inv1  gate613(.a(s_65), .O(gate107inter4));
  nand2 gate614(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate615(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate616(.a(N319), .O(gate107inter7));
  inv1  gate617(.a(N34), .O(gate107inter8));
  nand2 gate618(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate619(.a(s_65), .b(gate107inter3), .O(gate107inter10));
  nor2  gate620(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate621(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate622(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate273(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate274(.a(gate110inter0), .b(s_16), .O(gate110inter1));
  and2  gate275(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate276(.a(s_16), .O(gate110inter3));
  inv1  gate277(.a(s_17), .O(gate110inter4));
  nand2 gate278(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate279(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate280(.a(N309), .O(gate110inter7));
  inv1  gate281(.a(N282), .O(gate110inter8));
  nand2 gate282(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate283(.a(s_17), .b(gate110inter3), .O(gate110inter10));
  nor2  gate284(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate285(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate286(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );

  xor2  gate567(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate568(.a(gate112inter0), .b(s_58), .O(gate112inter1));
  and2  gate569(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate570(.a(s_58), .O(gate112inter3));
  inv1  gate571(.a(s_59), .O(gate112inter4));
  nand2 gate572(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate573(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate574(.a(N309), .O(gate112inter7));
  inv1  gate575(.a(N285), .O(gate112inter8));
  nand2 gate576(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate577(.a(s_59), .b(gate112inter3), .O(gate112inter10));
  nor2  gate578(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate579(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate580(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate637(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate638(.a(gate115inter0), .b(s_68), .O(gate115inter1));
  and2  gate639(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate640(.a(s_68), .O(gate115inter3));
  inv1  gate641(.a(s_69), .O(gate115inter4));
  nand2 gate642(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate643(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate644(.a(N319), .O(gate115inter7));
  inv1  gate645(.a(N99), .O(gate115inter8));
  nand2 gate646(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate647(.a(s_69), .b(gate115inter3), .O(gate115inter10));
  nor2  gate648(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate649(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate650(.a(gate115inter12), .b(gate115inter1), .O(N346));

  xor2  gate469(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate470(.a(gate116inter0), .b(s_44), .O(gate116inter1));
  and2  gate471(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate472(.a(s_44), .O(gate116inter3));
  inv1  gate473(.a(s_45), .O(gate116inter4));
  nand2 gate474(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate475(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate476(.a(N319), .O(gate116inter7));
  inv1  gate477(.a(N112), .O(gate116inter8));
  nand2 gate478(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate479(.a(s_45), .b(gate116inter3), .O(gate116inter10));
  nor2  gate480(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate481(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate482(.a(gate116inter12), .b(gate116inter1), .O(N347));
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate175(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate176(.a(gate121inter0), .b(s_2), .O(gate121inter1));
  and2  gate177(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate178(.a(s_2), .O(gate121inter3));
  inv1  gate179(.a(s_3), .O(gate121inter4));
  nand2 gate180(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate181(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate182(.a(N335), .O(gate121inter7));
  inv1  gate183(.a(N304), .O(gate121inter8));
  nand2 gate184(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate185(.a(s_3), .b(gate121inter3), .O(gate121inter10));
  nor2  gate186(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate187(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate188(.a(gate121inter12), .b(gate121inter1), .O(N352));

  xor2  gate707(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate708(.a(gate122inter0), .b(s_78), .O(gate122inter1));
  and2  gate709(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate710(.a(s_78), .O(gate122inter3));
  inv1  gate711(.a(s_79), .O(gate122inter4));
  nand2 gate712(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate713(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate714(.a(N337), .O(gate122inter7));
  inv1  gate715(.a(N305), .O(gate122inter8));
  nand2 gate716(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate717(.a(s_79), .b(gate122inter3), .O(gate122inter10));
  nor2  gate718(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate719(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate720(.a(gate122inter12), .b(gate122inter1), .O(N353));

  xor2  gate721(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate722(.a(gate123inter0), .b(s_80), .O(gate123inter1));
  and2  gate723(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate724(.a(s_80), .O(gate123inter3));
  inv1  gate725(.a(s_81), .O(gate123inter4));
  nand2 gate726(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate727(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate728(.a(N339), .O(gate123inter7));
  inv1  gate729(.a(N306), .O(gate123inter8));
  nand2 gate730(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate731(.a(s_81), .b(gate123inter3), .O(gate123inter10));
  nor2  gate732(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate733(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate734(.a(gate123inter12), .b(gate123inter1), .O(N354));

  xor2  gate763(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate764(.a(gate124inter0), .b(s_86), .O(gate124inter1));
  and2  gate765(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate766(.a(s_86), .O(gate124inter3));
  inv1  gate767(.a(s_87), .O(gate124inter4));
  nand2 gate768(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate769(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate770(.a(N341), .O(gate124inter7));
  inv1  gate771(.a(N307), .O(gate124inter8));
  nand2 gate772(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate773(.a(s_87), .b(gate124inter3), .O(gate124inter10));
  nor2  gate774(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate775(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate776(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate497(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate498(.a(gate131inter0), .b(s_48), .O(gate131inter1));
  and2  gate499(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate500(.a(s_48), .O(gate131inter3));
  inv1  gate501(.a(s_49), .O(gate131inter4));
  nand2 gate502(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate503(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate504(.a(N360), .O(gate131inter7));
  inv1  gate505(.a(N40), .O(gate131inter8));
  nand2 gate506(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate507(.a(s_49), .b(gate131inter3), .O(gate131inter10));
  nor2  gate508(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate509(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate510(.a(gate131inter12), .b(gate131inter1), .O(N373));

  xor2  gate329(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate330(.a(gate132inter0), .b(s_24), .O(gate132inter1));
  and2  gate331(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate332(.a(s_24), .O(gate132inter3));
  inv1  gate333(.a(s_25), .O(gate132inter4));
  nand2 gate334(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate335(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate336(.a(N360), .O(gate132inter7));
  inv1  gate337(.a(N53), .O(gate132inter8));
  nand2 gate338(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate339(.a(s_25), .b(gate132inter3), .O(gate132inter10));
  nor2  gate340(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate341(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate342(.a(gate132inter12), .b(gate132inter1), .O(N374));

  xor2  gate217(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate218(.a(gate133inter0), .b(s_8), .O(gate133inter1));
  and2  gate219(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate220(.a(s_8), .O(gate133inter3));
  inv1  gate221(.a(s_9), .O(gate133inter4));
  nand2 gate222(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate223(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate224(.a(N360), .O(gate133inter7));
  inv1  gate225(.a(N66), .O(gate133inter8));
  nand2 gate226(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate227(.a(s_9), .b(gate133inter3), .O(gate133inter10));
  nor2  gate228(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate229(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate230(.a(gate133inter12), .b(gate133inter1), .O(N375));

  xor2  gate525(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate526(.a(gate134inter0), .b(s_52), .O(gate134inter1));
  and2  gate527(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate528(.a(s_52), .O(gate134inter3));
  inv1  gate529(.a(s_53), .O(gate134inter4));
  nand2 gate530(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate531(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate532(.a(N360), .O(gate134inter7));
  inv1  gate533(.a(N79), .O(gate134inter8));
  nand2 gate534(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate535(.a(s_53), .b(gate134inter3), .O(gate134inter10));
  nor2  gate536(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate537(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate538(.a(gate134inter12), .b(gate134inter1), .O(N376));

  xor2  gate343(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate344(.a(gate135inter0), .b(s_26), .O(gate135inter1));
  and2  gate345(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate346(.a(s_26), .O(gate135inter3));
  inv1  gate347(.a(s_27), .O(gate135inter4));
  nand2 gate348(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate349(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate350(.a(N360), .O(gate135inter7));
  inv1  gate351(.a(N92), .O(gate135inter8));
  nand2 gate352(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate353(.a(s_27), .b(gate135inter3), .O(gate135inter10));
  nor2  gate354(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate355(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate356(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate623(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate624(.a(gate153inter0), .b(s_66), .O(gate153inter1));
  and2  gate625(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate626(.a(s_66), .O(gate153inter3));
  inv1  gate627(.a(s_67), .O(gate153inter4));
  nand2 gate628(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate629(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate630(.a(N415), .O(gate153inter7));
  inv1  gate631(.a(N416), .O(gate153inter8));
  nand2 gate632(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate633(.a(s_67), .b(gate153inter3), .O(gate153inter10));
  nor2  gate634(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate635(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate636(.a(gate153inter12), .b(gate153inter1), .O(N421));
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule