module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1107(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1108(.a(gate9inter0), .b(s_80), .O(gate9inter1));
  and2  gate1109(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1110(.a(s_80), .O(gate9inter3));
  inv1  gate1111(.a(s_81), .O(gate9inter4));
  nand2 gate1112(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1113(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1114(.a(G1), .O(gate9inter7));
  inv1  gate1115(.a(G2), .O(gate9inter8));
  nand2 gate1116(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1117(.a(s_81), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1118(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1119(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1120(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1205(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1206(.a(gate26inter0), .b(s_94), .O(gate26inter1));
  and2  gate1207(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1208(.a(s_94), .O(gate26inter3));
  inv1  gate1209(.a(s_95), .O(gate26inter4));
  nand2 gate1210(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1211(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1212(.a(G9), .O(gate26inter7));
  inv1  gate1213(.a(G13), .O(gate26inter8));
  nand2 gate1214(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1215(.a(s_95), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1216(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1217(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1218(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1093(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1094(.a(gate36inter0), .b(s_78), .O(gate36inter1));
  and2  gate1095(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1096(.a(s_78), .O(gate36inter3));
  inv1  gate1097(.a(s_79), .O(gate36inter4));
  nand2 gate1098(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1099(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1100(.a(G26), .O(gate36inter7));
  inv1  gate1101(.a(G30), .O(gate36inter8));
  nand2 gate1102(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1103(.a(s_79), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1104(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1105(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1106(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate813(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate814(.a(gate38inter0), .b(s_38), .O(gate38inter1));
  and2  gate815(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate816(.a(s_38), .O(gate38inter3));
  inv1  gate817(.a(s_39), .O(gate38inter4));
  nand2 gate818(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate819(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate820(.a(G27), .O(gate38inter7));
  inv1  gate821(.a(G31), .O(gate38inter8));
  nand2 gate822(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate823(.a(s_39), .b(gate38inter3), .O(gate38inter10));
  nor2  gate824(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate825(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate826(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1219(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1220(.a(gate52inter0), .b(s_96), .O(gate52inter1));
  and2  gate1221(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1222(.a(s_96), .O(gate52inter3));
  inv1  gate1223(.a(s_97), .O(gate52inter4));
  nand2 gate1224(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1225(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1226(.a(G12), .O(gate52inter7));
  inv1  gate1227(.a(G281), .O(gate52inter8));
  nand2 gate1228(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1229(.a(s_97), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1230(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1231(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1232(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1163(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1164(.a(gate60inter0), .b(s_88), .O(gate60inter1));
  and2  gate1165(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1166(.a(s_88), .O(gate60inter3));
  inv1  gate1167(.a(s_89), .O(gate60inter4));
  nand2 gate1168(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1169(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1170(.a(G20), .O(gate60inter7));
  inv1  gate1171(.a(G293), .O(gate60inter8));
  nand2 gate1172(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1173(.a(s_89), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1174(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1175(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1176(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate701(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate702(.a(gate62inter0), .b(s_22), .O(gate62inter1));
  and2  gate703(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate704(.a(s_22), .O(gate62inter3));
  inv1  gate705(.a(s_23), .O(gate62inter4));
  nand2 gate706(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate707(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate708(.a(G22), .O(gate62inter7));
  inv1  gate709(.a(G296), .O(gate62inter8));
  nand2 gate710(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate711(.a(s_23), .b(gate62inter3), .O(gate62inter10));
  nor2  gate712(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate713(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate714(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate785(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate786(.a(gate65inter0), .b(s_34), .O(gate65inter1));
  and2  gate787(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate788(.a(s_34), .O(gate65inter3));
  inv1  gate789(.a(s_35), .O(gate65inter4));
  nand2 gate790(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate791(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate792(.a(G25), .O(gate65inter7));
  inv1  gate793(.a(G302), .O(gate65inter8));
  nand2 gate794(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate795(.a(s_35), .b(gate65inter3), .O(gate65inter10));
  nor2  gate796(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate797(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate798(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate729(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate730(.a(gate77inter0), .b(s_26), .O(gate77inter1));
  and2  gate731(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate732(.a(s_26), .O(gate77inter3));
  inv1  gate733(.a(s_27), .O(gate77inter4));
  nand2 gate734(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate735(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate736(.a(G2), .O(gate77inter7));
  inv1  gate737(.a(G320), .O(gate77inter8));
  nand2 gate738(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate739(.a(s_27), .b(gate77inter3), .O(gate77inter10));
  nor2  gate740(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate741(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate742(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1149(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1150(.a(gate79inter0), .b(s_86), .O(gate79inter1));
  and2  gate1151(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1152(.a(s_86), .O(gate79inter3));
  inv1  gate1153(.a(s_87), .O(gate79inter4));
  nand2 gate1154(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1155(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1156(.a(G10), .O(gate79inter7));
  inv1  gate1157(.a(G323), .O(gate79inter8));
  nand2 gate1158(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1159(.a(s_87), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1160(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1161(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1162(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate953(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate954(.a(gate90inter0), .b(s_58), .O(gate90inter1));
  and2  gate955(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate956(.a(s_58), .O(gate90inter3));
  inv1  gate957(.a(s_59), .O(gate90inter4));
  nand2 gate958(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate959(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate960(.a(G21), .O(gate90inter7));
  inv1  gate961(.a(G338), .O(gate90inter8));
  nand2 gate962(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate963(.a(s_59), .b(gate90inter3), .O(gate90inter10));
  nor2  gate964(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate965(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate966(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate757(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate758(.a(gate92inter0), .b(s_30), .O(gate92inter1));
  and2  gate759(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate760(.a(s_30), .O(gate92inter3));
  inv1  gate761(.a(s_31), .O(gate92inter4));
  nand2 gate762(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate763(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate764(.a(G29), .O(gate92inter7));
  inv1  gate765(.a(G341), .O(gate92inter8));
  nand2 gate766(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate767(.a(s_31), .b(gate92inter3), .O(gate92inter10));
  nor2  gate768(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate769(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate770(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate743(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate744(.a(gate96inter0), .b(s_28), .O(gate96inter1));
  and2  gate745(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate746(.a(s_28), .O(gate96inter3));
  inv1  gate747(.a(s_29), .O(gate96inter4));
  nand2 gate748(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate749(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate750(.a(G30), .O(gate96inter7));
  inv1  gate751(.a(G347), .O(gate96inter8));
  nand2 gate752(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate753(.a(s_29), .b(gate96inter3), .O(gate96inter10));
  nor2  gate754(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate755(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate756(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1135(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1136(.a(gate97inter0), .b(s_84), .O(gate97inter1));
  and2  gate1137(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1138(.a(s_84), .O(gate97inter3));
  inv1  gate1139(.a(s_85), .O(gate97inter4));
  nand2 gate1140(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1141(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1142(.a(G19), .O(gate97inter7));
  inv1  gate1143(.a(G350), .O(gate97inter8));
  nand2 gate1144(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1145(.a(s_85), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1146(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1147(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1148(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate603(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate604(.a(gate136inter0), .b(s_8), .O(gate136inter1));
  and2  gate605(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate606(.a(s_8), .O(gate136inter3));
  inv1  gate607(.a(s_9), .O(gate136inter4));
  nand2 gate608(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate609(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate610(.a(G424), .O(gate136inter7));
  inv1  gate611(.a(G425), .O(gate136inter8));
  nand2 gate612(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate613(.a(s_9), .b(gate136inter3), .O(gate136inter10));
  nor2  gate614(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate615(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate616(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1387(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1388(.a(gate138inter0), .b(s_120), .O(gate138inter1));
  and2  gate1389(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1390(.a(s_120), .O(gate138inter3));
  inv1  gate1391(.a(s_121), .O(gate138inter4));
  nand2 gate1392(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1393(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1394(.a(G432), .O(gate138inter7));
  inv1  gate1395(.a(G435), .O(gate138inter8));
  nand2 gate1396(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1397(.a(s_121), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1398(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1399(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1400(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1359(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1360(.a(gate143inter0), .b(s_116), .O(gate143inter1));
  and2  gate1361(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1362(.a(s_116), .O(gate143inter3));
  inv1  gate1363(.a(s_117), .O(gate143inter4));
  nand2 gate1364(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1365(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1366(.a(G462), .O(gate143inter7));
  inv1  gate1367(.a(G465), .O(gate143inter8));
  nand2 gate1368(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1369(.a(s_117), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1370(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1371(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1372(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate897(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate898(.a(gate151inter0), .b(s_50), .O(gate151inter1));
  and2  gate899(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate900(.a(s_50), .O(gate151inter3));
  inv1  gate901(.a(s_51), .O(gate151inter4));
  nand2 gate902(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate903(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate904(.a(G510), .O(gate151inter7));
  inv1  gate905(.a(G513), .O(gate151inter8));
  nand2 gate906(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate907(.a(s_51), .b(gate151inter3), .O(gate151inter10));
  nor2  gate908(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate909(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate910(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate659(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate660(.a(gate161inter0), .b(s_16), .O(gate161inter1));
  and2  gate661(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate662(.a(s_16), .O(gate161inter3));
  inv1  gate663(.a(s_17), .O(gate161inter4));
  nand2 gate664(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate665(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate666(.a(G450), .O(gate161inter7));
  inv1  gate667(.a(G534), .O(gate161inter8));
  nand2 gate668(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate669(.a(s_17), .b(gate161inter3), .O(gate161inter10));
  nor2  gate670(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate671(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate672(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1009(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1010(.a(gate164inter0), .b(s_66), .O(gate164inter1));
  and2  gate1011(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1012(.a(s_66), .O(gate164inter3));
  inv1  gate1013(.a(s_67), .O(gate164inter4));
  nand2 gate1014(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1015(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1016(.a(G459), .O(gate164inter7));
  inv1  gate1017(.a(G537), .O(gate164inter8));
  nand2 gate1018(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1019(.a(s_67), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1020(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1021(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1022(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate617(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate618(.a(gate167inter0), .b(s_10), .O(gate167inter1));
  and2  gate619(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate620(.a(s_10), .O(gate167inter3));
  inv1  gate621(.a(s_11), .O(gate167inter4));
  nand2 gate622(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate623(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate624(.a(G468), .O(gate167inter7));
  inv1  gate625(.a(G543), .O(gate167inter8));
  nand2 gate626(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate627(.a(s_11), .b(gate167inter3), .O(gate167inter10));
  nor2  gate628(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate629(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate630(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1261(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1262(.a(gate170inter0), .b(s_102), .O(gate170inter1));
  and2  gate1263(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1264(.a(s_102), .O(gate170inter3));
  inv1  gate1265(.a(s_103), .O(gate170inter4));
  nand2 gate1266(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1267(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1268(.a(G477), .O(gate170inter7));
  inv1  gate1269(.a(G546), .O(gate170inter8));
  nand2 gate1270(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1271(.a(s_103), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1272(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1273(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1274(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1023(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1024(.a(gate174inter0), .b(s_68), .O(gate174inter1));
  and2  gate1025(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1026(.a(s_68), .O(gate174inter3));
  inv1  gate1027(.a(s_69), .O(gate174inter4));
  nand2 gate1028(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1029(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1030(.a(G489), .O(gate174inter7));
  inv1  gate1031(.a(G552), .O(gate174inter8));
  nand2 gate1032(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1033(.a(s_69), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1034(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1035(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1036(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate715(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate716(.a(gate180inter0), .b(s_24), .O(gate180inter1));
  and2  gate717(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate718(.a(s_24), .O(gate180inter3));
  inv1  gate719(.a(s_25), .O(gate180inter4));
  nand2 gate720(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate721(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate722(.a(G507), .O(gate180inter7));
  inv1  gate723(.a(G561), .O(gate180inter8));
  nand2 gate724(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate725(.a(s_25), .b(gate180inter3), .O(gate180inter10));
  nor2  gate726(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate727(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate728(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1275(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1276(.a(gate184inter0), .b(s_104), .O(gate184inter1));
  and2  gate1277(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1278(.a(s_104), .O(gate184inter3));
  inv1  gate1279(.a(s_105), .O(gate184inter4));
  nand2 gate1280(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1281(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1282(.a(G519), .O(gate184inter7));
  inv1  gate1283(.a(G567), .O(gate184inter8));
  nand2 gate1284(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1285(.a(s_105), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1286(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1287(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1288(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1233(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1234(.a(gate192inter0), .b(s_98), .O(gate192inter1));
  and2  gate1235(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1236(.a(s_98), .O(gate192inter3));
  inv1  gate1237(.a(s_99), .O(gate192inter4));
  nand2 gate1238(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1239(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1240(.a(G584), .O(gate192inter7));
  inv1  gate1241(.a(G585), .O(gate192inter8));
  nand2 gate1242(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1243(.a(s_99), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1244(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1245(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1246(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1065(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1066(.a(gate194inter0), .b(s_74), .O(gate194inter1));
  and2  gate1067(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1068(.a(s_74), .O(gate194inter3));
  inv1  gate1069(.a(s_75), .O(gate194inter4));
  nand2 gate1070(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1071(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1072(.a(G588), .O(gate194inter7));
  inv1  gate1073(.a(G589), .O(gate194inter8));
  nand2 gate1074(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1075(.a(s_75), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1076(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1077(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1078(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1317(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1318(.a(gate196inter0), .b(s_110), .O(gate196inter1));
  and2  gate1319(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1320(.a(s_110), .O(gate196inter3));
  inv1  gate1321(.a(s_111), .O(gate196inter4));
  nand2 gate1322(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1323(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1324(.a(G592), .O(gate196inter7));
  inv1  gate1325(.a(G593), .O(gate196inter8));
  nand2 gate1326(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1327(.a(s_111), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1328(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1329(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1330(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate687(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate688(.a(gate201inter0), .b(s_20), .O(gate201inter1));
  and2  gate689(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate690(.a(s_20), .O(gate201inter3));
  inv1  gate691(.a(s_21), .O(gate201inter4));
  nand2 gate692(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate693(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate694(.a(G602), .O(gate201inter7));
  inv1  gate695(.a(G607), .O(gate201inter8));
  nand2 gate696(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate697(.a(s_21), .b(gate201inter3), .O(gate201inter10));
  nor2  gate698(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate699(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate700(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate981(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate982(.a(gate202inter0), .b(s_62), .O(gate202inter1));
  and2  gate983(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate984(.a(s_62), .O(gate202inter3));
  inv1  gate985(.a(s_63), .O(gate202inter4));
  nand2 gate986(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate987(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate988(.a(G612), .O(gate202inter7));
  inv1  gate989(.a(G617), .O(gate202inter8));
  nand2 gate990(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate991(.a(s_63), .b(gate202inter3), .O(gate202inter10));
  nor2  gate992(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate993(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate994(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate939(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate940(.a(gate208inter0), .b(s_56), .O(gate208inter1));
  and2  gate941(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate942(.a(s_56), .O(gate208inter3));
  inv1  gate943(.a(s_57), .O(gate208inter4));
  nand2 gate944(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate945(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate946(.a(G627), .O(gate208inter7));
  inv1  gate947(.a(G637), .O(gate208inter8));
  nand2 gate948(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate949(.a(s_57), .b(gate208inter3), .O(gate208inter10));
  nor2  gate950(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate951(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate952(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate575(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate576(.a(gate209inter0), .b(s_4), .O(gate209inter1));
  and2  gate577(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate578(.a(s_4), .O(gate209inter3));
  inv1  gate579(.a(s_5), .O(gate209inter4));
  nand2 gate580(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate581(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate582(.a(G602), .O(gate209inter7));
  inv1  gate583(.a(G666), .O(gate209inter8));
  nand2 gate584(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate585(.a(s_5), .b(gate209inter3), .O(gate209inter10));
  nor2  gate586(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate587(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate588(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate967(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate968(.a(gate210inter0), .b(s_60), .O(gate210inter1));
  and2  gate969(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate970(.a(s_60), .O(gate210inter3));
  inv1  gate971(.a(s_61), .O(gate210inter4));
  nand2 gate972(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate973(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate974(.a(G607), .O(gate210inter7));
  inv1  gate975(.a(G666), .O(gate210inter8));
  nand2 gate976(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate977(.a(s_61), .b(gate210inter3), .O(gate210inter10));
  nor2  gate978(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate979(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate980(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1079(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1080(.a(gate232inter0), .b(s_76), .O(gate232inter1));
  and2  gate1081(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1082(.a(s_76), .O(gate232inter3));
  inv1  gate1083(.a(s_77), .O(gate232inter4));
  nand2 gate1084(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1085(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1086(.a(G704), .O(gate232inter7));
  inv1  gate1087(.a(G705), .O(gate232inter8));
  nand2 gate1088(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1089(.a(s_77), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1090(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1091(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1092(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate589(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate590(.a(gate238inter0), .b(s_6), .O(gate238inter1));
  and2  gate591(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate592(.a(s_6), .O(gate238inter3));
  inv1  gate593(.a(s_7), .O(gate238inter4));
  nand2 gate594(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate595(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate596(.a(G257), .O(gate238inter7));
  inv1  gate597(.a(G709), .O(gate238inter8));
  nand2 gate598(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate599(.a(s_7), .b(gate238inter3), .O(gate238inter10));
  nor2  gate600(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate601(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate602(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate827(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate828(.a(gate240inter0), .b(s_40), .O(gate240inter1));
  and2  gate829(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate830(.a(s_40), .O(gate240inter3));
  inv1  gate831(.a(s_41), .O(gate240inter4));
  nand2 gate832(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate833(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate834(.a(G263), .O(gate240inter7));
  inv1  gate835(.a(G715), .O(gate240inter8));
  nand2 gate836(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate837(.a(s_41), .b(gate240inter3), .O(gate240inter10));
  nor2  gate838(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate839(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate840(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate561(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate562(.a(gate264inter0), .b(s_2), .O(gate264inter1));
  and2  gate563(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate564(.a(s_2), .O(gate264inter3));
  inv1  gate565(.a(s_3), .O(gate264inter4));
  nand2 gate566(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate567(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate568(.a(G768), .O(gate264inter7));
  inv1  gate569(.a(G769), .O(gate264inter8));
  nand2 gate570(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate571(.a(s_3), .b(gate264inter3), .O(gate264inter10));
  nor2  gate572(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate573(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate574(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1191(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1192(.a(gate273inter0), .b(s_92), .O(gate273inter1));
  and2  gate1193(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1194(.a(s_92), .O(gate273inter3));
  inv1  gate1195(.a(s_93), .O(gate273inter4));
  nand2 gate1196(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1197(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1198(.a(G642), .O(gate273inter7));
  inv1  gate1199(.a(G794), .O(gate273inter8));
  nand2 gate1200(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1201(.a(s_93), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1202(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1203(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1204(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1373(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1374(.a(gate279inter0), .b(s_118), .O(gate279inter1));
  and2  gate1375(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1376(.a(s_118), .O(gate279inter3));
  inv1  gate1377(.a(s_119), .O(gate279inter4));
  nand2 gate1378(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1379(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1380(.a(G651), .O(gate279inter7));
  inv1  gate1381(.a(G803), .O(gate279inter8));
  nand2 gate1382(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1383(.a(s_119), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1384(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1385(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1386(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1303(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1304(.a(gate280inter0), .b(s_108), .O(gate280inter1));
  and2  gate1305(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1306(.a(s_108), .O(gate280inter3));
  inv1  gate1307(.a(s_109), .O(gate280inter4));
  nand2 gate1308(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1309(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1310(.a(G779), .O(gate280inter7));
  inv1  gate1311(.a(G803), .O(gate280inter8));
  nand2 gate1312(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1313(.a(s_109), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1314(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1315(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1316(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate841(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate842(.a(gate396inter0), .b(s_42), .O(gate396inter1));
  and2  gate843(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate844(.a(s_42), .O(gate396inter3));
  inv1  gate845(.a(s_43), .O(gate396inter4));
  nand2 gate846(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate847(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate848(.a(G10), .O(gate396inter7));
  inv1  gate849(.a(G1063), .O(gate396inter8));
  nand2 gate850(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate851(.a(s_43), .b(gate396inter3), .O(gate396inter10));
  nor2  gate852(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate853(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate854(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate799(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate800(.a(gate398inter0), .b(s_36), .O(gate398inter1));
  and2  gate801(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate802(.a(s_36), .O(gate398inter3));
  inv1  gate803(.a(s_37), .O(gate398inter4));
  nand2 gate804(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate805(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate806(.a(G12), .O(gate398inter7));
  inv1  gate807(.a(G1069), .O(gate398inter8));
  nand2 gate808(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate809(.a(s_37), .b(gate398inter3), .O(gate398inter10));
  nor2  gate810(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate811(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate812(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1247(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1248(.a(gate405inter0), .b(s_100), .O(gate405inter1));
  and2  gate1249(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1250(.a(s_100), .O(gate405inter3));
  inv1  gate1251(.a(s_101), .O(gate405inter4));
  nand2 gate1252(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1253(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1254(.a(G19), .O(gate405inter7));
  inv1  gate1255(.a(G1090), .O(gate405inter8));
  nand2 gate1256(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1257(.a(s_101), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1258(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1259(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1260(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate925(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate926(.a(gate408inter0), .b(s_54), .O(gate408inter1));
  and2  gate927(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate928(.a(s_54), .O(gate408inter3));
  inv1  gate929(.a(s_55), .O(gate408inter4));
  nand2 gate930(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate931(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate932(.a(G22), .O(gate408inter7));
  inv1  gate933(.a(G1099), .O(gate408inter8));
  nand2 gate934(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate935(.a(s_55), .b(gate408inter3), .O(gate408inter10));
  nor2  gate936(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate937(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate938(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1177(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1178(.a(gate421inter0), .b(s_90), .O(gate421inter1));
  and2  gate1179(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1180(.a(s_90), .O(gate421inter3));
  inv1  gate1181(.a(s_91), .O(gate421inter4));
  nand2 gate1182(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1183(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1184(.a(G2), .O(gate421inter7));
  inv1  gate1185(.a(G1135), .O(gate421inter8));
  nand2 gate1186(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1187(.a(s_91), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1188(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1189(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1190(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate855(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate856(.a(gate425inter0), .b(s_44), .O(gate425inter1));
  and2  gate857(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate858(.a(s_44), .O(gate425inter3));
  inv1  gate859(.a(s_45), .O(gate425inter4));
  nand2 gate860(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate861(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate862(.a(G4), .O(gate425inter7));
  inv1  gate863(.a(G1141), .O(gate425inter8));
  nand2 gate864(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate865(.a(s_45), .b(gate425inter3), .O(gate425inter10));
  nor2  gate866(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate867(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate868(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1037(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1038(.a(gate427inter0), .b(s_70), .O(gate427inter1));
  and2  gate1039(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1040(.a(s_70), .O(gate427inter3));
  inv1  gate1041(.a(s_71), .O(gate427inter4));
  nand2 gate1042(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1043(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1044(.a(G5), .O(gate427inter7));
  inv1  gate1045(.a(G1144), .O(gate427inter8));
  nand2 gate1046(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1047(.a(s_71), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1048(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1049(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1050(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1051(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1052(.a(gate431inter0), .b(s_72), .O(gate431inter1));
  and2  gate1053(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1054(.a(s_72), .O(gate431inter3));
  inv1  gate1055(.a(s_73), .O(gate431inter4));
  nand2 gate1056(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1057(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1058(.a(G7), .O(gate431inter7));
  inv1  gate1059(.a(G1150), .O(gate431inter8));
  nand2 gate1060(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1061(.a(s_73), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1062(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1063(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1064(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1345(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1346(.a(gate441inter0), .b(s_114), .O(gate441inter1));
  and2  gate1347(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1348(.a(s_114), .O(gate441inter3));
  inv1  gate1349(.a(s_115), .O(gate441inter4));
  nand2 gate1350(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1351(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1352(.a(G12), .O(gate441inter7));
  inv1  gate1353(.a(G1165), .O(gate441inter8));
  nand2 gate1354(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1355(.a(s_115), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1356(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1357(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1358(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate645(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate646(.a(gate443inter0), .b(s_14), .O(gate443inter1));
  and2  gate647(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate648(.a(s_14), .O(gate443inter3));
  inv1  gate649(.a(s_15), .O(gate443inter4));
  nand2 gate650(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate651(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate652(.a(G13), .O(gate443inter7));
  inv1  gate653(.a(G1168), .O(gate443inter8));
  nand2 gate654(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate655(.a(s_15), .b(gate443inter3), .O(gate443inter10));
  nor2  gate656(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate657(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate658(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1331(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1332(.a(gate446inter0), .b(s_112), .O(gate446inter1));
  and2  gate1333(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1334(.a(s_112), .O(gate446inter3));
  inv1  gate1335(.a(s_113), .O(gate446inter4));
  nand2 gate1336(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1337(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1338(.a(G1075), .O(gate446inter7));
  inv1  gate1339(.a(G1171), .O(gate446inter8));
  nand2 gate1340(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1341(.a(s_113), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1342(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1343(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1344(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate995(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate996(.a(gate455inter0), .b(s_64), .O(gate455inter1));
  and2  gate997(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate998(.a(s_64), .O(gate455inter3));
  inv1  gate999(.a(s_65), .O(gate455inter4));
  nand2 gate1000(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1001(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1002(.a(G19), .O(gate455inter7));
  inv1  gate1003(.a(G1186), .O(gate455inter8));
  nand2 gate1004(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1005(.a(s_65), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1006(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1007(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1008(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate673(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate674(.a(gate465inter0), .b(s_18), .O(gate465inter1));
  and2  gate675(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate676(.a(s_18), .O(gate465inter3));
  inv1  gate677(.a(s_19), .O(gate465inter4));
  nand2 gate678(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate679(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate680(.a(G24), .O(gate465inter7));
  inv1  gate681(.a(G1201), .O(gate465inter8));
  nand2 gate682(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate683(.a(s_19), .b(gate465inter3), .O(gate465inter10));
  nor2  gate684(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate685(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate686(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate547(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate548(.a(gate466inter0), .b(s_0), .O(gate466inter1));
  and2  gate549(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate550(.a(s_0), .O(gate466inter3));
  inv1  gate551(.a(s_1), .O(gate466inter4));
  nand2 gate552(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate553(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate554(.a(G1105), .O(gate466inter7));
  inv1  gate555(.a(G1201), .O(gate466inter8));
  nand2 gate556(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate557(.a(s_1), .b(gate466inter3), .O(gate466inter10));
  nor2  gate558(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate559(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate560(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate631(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate632(.a(gate480inter0), .b(s_12), .O(gate480inter1));
  and2  gate633(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate634(.a(s_12), .O(gate480inter3));
  inv1  gate635(.a(s_13), .O(gate480inter4));
  nand2 gate636(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate637(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate638(.a(G1126), .O(gate480inter7));
  inv1  gate639(.a(G1222), .O(gate480inter8));
  nand2 gate640(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate641(.a(s_13), .b(gate480inter3), .O(gate480inter10));
  nor2  gate642(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate643(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate644(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1289(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1290(.a(gate482inter0), .b(s_106), .O(gate482inter1));
  and2  gate1291(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1292(.a(s_106), .O(gate482inter3));
  inv1  gate1293(.a(s_107), .O(gate482inter4));
  nand2 gate1294(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1295(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1296(.a(G1129), .O(gate482inter7));
  inv1  gate1297(.a(G1225), .O(gate482inter8));
  nand2 gate1298(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1299(.a(s_107), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1300(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1301(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1302(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate883(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate884(.a(gate483inter0), .b(s_48), .O(gate483inter1));
  and2  gate885(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate886(.a(s_48), .O(gate483inter3));
  inv1  gate887(.a(s_49), .O(gate483inter4));
  nand2 gate888(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate889(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate890(.a(G1228), .O(gate483inter7));
  inv1  gate891(.a(G1229), .O(gate483inter8));
  nand2 gate892(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate893(.a(s_49), .b(gate483inter3), .O(gate483inter10));
  nor2  gate894(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate895(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate896(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1121(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1122(.a(gate490inter0), .b(s_82), .O(gate490inter1));
  and2  gate1123(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1124(.a(s_82), .O(gate490inter3));
  inv1  gate1125(.a(s_83), .O(gate490inter4));
  nand2 gate1126(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1127(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1128(.a(G1242), .O(gate490inter7));
  inv1  gate1129(.a(G1243), .O(gate490inter8));
  nand2 gate1130(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1131(.a(s_83), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1132(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1133(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1134(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate911(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate912(.a(gate494inter0), .b(s_52), .O(gate494inter1));
  and2  gate913(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate914(.a(s_52), .O(gate494inter3));
  inv1  gate915(.a(s_53), .O(gate494inter4));
  nand2 gate916(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate917(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate918(.a(G1250), .O(gate494inter7));
  inv1  gate919(.a(G1251), .O(gate494inter8));
  nand2 gate920(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate921(.a(s_53), .b(gate494inter3), .O(gate494inter10));
  nor2  gate922(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate923(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate924(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate771(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate772(.a(gate510inter0), .b(s_32), .O(gate510inter1));
  and2  gate773(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate774(.a(s_32), .O(gate510inter3));
  inv1  gate775(.a(s_33), .O(gate510inter4));
  nand2 gate776(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate777(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate778(.a(G1282), .O(gate510inter7));
  inv1  gate779(.a(G1283), .O(gate510inter8));
  nand2 gate780(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate781(.a(s_33), .b(gate510inter3), .O(gate510inter10));
  nor2  gate782(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate783(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate784(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate869(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate870(.a(gate514inter0), .b(s_46), .O(gate514inter1));
  and2  gate871(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate872(.a(s_46), .O(gate514inter3));
  inv1  gate873(.a(s_47), .O(gate514inter4));
  nand2 gate874(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate875(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate876(.a(G1290), .O(gate514inter7));
  inv1  gate877(.a(G1291), .O(gate514inter8));
  nand2 gate878(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate879(.a(s_47), .b(gate514inter3), .O(gate514inter10));
  nor2  gate880(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate881(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate882(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule