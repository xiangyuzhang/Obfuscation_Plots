module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1387(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1388(.a(gate20inter0), .b(s_120), .O(gate20inter1));
  and2  gate1389(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1390(.a(s_120), .O(gate20inter3));
  inv1  gate1391(.a(s_121), .O(gate20inter4));
  nand2 gate1392(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1393(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1394(.a(G23), .O(gate20inter7));
  inv1  gate1395(.a(G24), .O(gate20inter8));
  nand2 gate1396(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1397(.a(s_121), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1398(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1399(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1400(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1779(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1780(.a(gate27inter0), .b(s_176), .O(gate27inter1));
  and2  gate1781(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1782(.a(s_176), .O(gate27inter3));
  inv1  gate1783(.a(s_177), .O(gate27inter4));
  nand2 gate1784(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1785(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1786(.a(G2), .O(gate27inter7));
  inv1  gate1787(.a(G6), .O(gate27inter8));
  nand2 gate1788(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1789(.a(s_177), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1790(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1791(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1792(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2171(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2172(.a(gate32inter0), .b(s_232), .O(gate32inter1));
  and2  gate2173(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2174(.a(s_232), .O(gate32inter3));
  inv1  gate2175(.a(s_233), .O(gate32inter4));
  nand2 gate2176(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2177(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2178(.a(G12), .O(gate32inter7));
  inv1  gate2179(.a(G16), .O(gate32inter8));
  nand2 gate2180(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2181(.a(s_233), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2182(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2183(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2184(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate925(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate926(.a(gate33inter0), .b(s_54), .O(gate33inter1));
  and2  gate927(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate928(.a(s_54), .O(gate33inter3));
  inv1  gate929(.a(s_55), .O(gate33inter4));
  nand2 gate930(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate931(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate932(.a(G17), .O(gate33inter7));
  inv1  gate933(.a(G21), .O(gate33inter8));
  nand2 gate934(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate935(.a(s_55), .b(gate33inter3), .O(gate33inter10));
  nor2  gate936(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate937(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate938(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1835(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1836(.a(gate35inter0), .b(s_184), .O(gate35inter1));
  and2  gate1837(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1838(.a(s_184), .O(gate35inter3));
  inv1  gate1839(.a(s_185), .O(gate35inter4));
  nand2 gate1840(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1841(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1842(.a(G18), .O(gate35inter7));
  inv1  gate1843(.a(G22), .O(gate35inter8));
  nand2 gate1844(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1845(.a(s_185), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1846(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1847(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1848(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1303(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1304(.a(gate37inter0), .b(s_108), .O(gate37inter1));
  and2  gate1305(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1306(.a(s_108), .O(gate37inter3));
  inv1  gate1307(.a(s_109), .O(gate37inter4));
  nand2 gate1308(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1309(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1310(.a(G19), .O(gate37inter7));
  inv1  gate1311(.a(G23), .O(gate37inter8));
  nand2 gate1312(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1313(.a(s_109), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1314(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1315(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1316(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1583(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1584(.a(gate43inter0), .b(s_148), .O(gate43inter1));
  and2  gate1585(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1586(.a(s_148), .O(gate43inter3));
  inv1  gate1587(.a(s_149), .O(gate43inter4));
  nand2 gate1588(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1589(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1590(.a(G3), .O(gate43inter7));
  inv1  gate1591(.a(G269), .O(gate43inter8));
  nand2 gate1592(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1593(.a(s_149), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1594(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1595(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1596(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1555(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1556(.a(gate50inter0), .b(s_144), .O(gate50inter1));
  and2  gate1557(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1558(.a(s_144), .O(gate50inter3));
  inv1  gate1559(.a(s_145), .O(gate50inter4));
  nand2 gate1560(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1561(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1562(.a(G10), .O(gate50inter7));
  inv1  gate1563(.a(G278), .O(gate50inter8));
  nand2 gate1564(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1565(.a(s_145), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1566(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1567(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1568(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1373(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1374(.a(gate51inter0), .b(s_118), .O(gate51inter1));
  and2  gate1375(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1376(.a(s_118), .O(gate51inter3));
  inv1  gate1377(.a(s_119), .O(gate51inter4));
  nand2 gate1378(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1379(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1380(.a(G11), .O(gate51inter7));
  inv1  gate1381(.a(G281), .O(gate51inter8));
  nand2 gate1382(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1383(.a(s_119), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1384(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1385(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1386(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate939(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate940(.a(gate53inter0), .b(s_56), .O(gate53inter1));
  and2  gate941(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate942(.a(s_56), .O(gate53inter3));
  inv1  gate943(.a(s_57), .O(gate53inter4));
  nand2 gate944(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate945(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate946(.a(G13), .O(gate53inter7));
  inv1  gate947(.a(G284), .O(gate53inter8));
  nand2 gate948(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate949(.a(s_57), .b(gate53inter3), .O(gate53inter10));
  nor2  gate950(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate951(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate952(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate827(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate828(.a(gate59inter0), .b(s_40), .O(gate59inter1));
  and2  gate829(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate830(.a(s_40), .O(gate59inter3));
  inv1  gate831(.a(s_41), .O(gate59inter4));
  nand2 gate832(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate833(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate834(.a(G19), .O(gate59inter7));
  inv1  gate835(.a(G293), .O(gate59inter8));
  nand2 gate836(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate837(.a(s_41), .b(gate59inter3), .O(gate59inter10));
  nor2  gate838(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate839(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate840(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1345(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1346(.a(gate60inter0), .b(s_114), .O(gate60inter1));
  and2  gate1347(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1348(.a(s_114), .O(gate60inter3));
  inv1  gate1349(.a(s_115), .O(gate60inter4));
  nand2 gate1350(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1351(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1352(.a(G20), .O(gate60inter7));
  inv1  gate1353(.a(G293), .O(gate60inter8));
  nand2 gate1354(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1355(.a(s_115), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1356(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1357(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1358(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1961(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1962(.a(gate69inter0), .b(s_202), .O(gate69inter1));
  and2  gate1963(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1964(.a(s_202), .O(gate69inter3));
  inv1  gate1965(.a(s_203), .O(gate69inter4));
  nand2 gate1966(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1967(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1968(.a(G29), .O(gate69inter7));
  inv1  gate1969(.a(G308), .O(gate69inter8));
  nand2 gate1970(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1971(.a(s_203), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1972(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1973(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1974(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1947(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1948(.a(gate70inter0), .b(s_200), .O(gate70inter1));
  and2  gate1949(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1950(.a(s_200), .O(gate70inter3));
  inv1  gate1951(.a(s_201), .O(gate70inter4));
  nand2 gate1952(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1953(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1954(.a(G30), .O(gate70inter7));
  inv1  gate1955(.a(G308), .O(gate70inter8));
  nand2 gate1956(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1957(.a(s_201), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1958(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1959(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1960(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate729(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate730(.a(gate71inter0), .b(s_26), .O(gate71inter1));
  and2  gate731(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate732(.a(s_26), .O(gate71inter3));
  inv1  gate733(.a(s_27), .O(gate71inter4));
  nand2 gate734(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate735(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate736(.a(G31), .O(gate71inter7));
  inv1  gate737(.a(G311), .O(gate71inter8));
  nand2 gate738(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate739(.a(s_27), .b(gate71inter3), .O(gate71inter10));
  nor2  gate740(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate741(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate742(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate841(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate842(.a(gate72inter0), .b(s_42), .O(gate72inter1));
  and2  gate843(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate844(.a(s_42), .O(gate72inter3));
  inv1  gate845(.a(s_43), .O(gate72inter4));
  nand2 gate846(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate847(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate848(.a(G32), .O(gate72inter7));
  inv1  gate849(.a(G311), .O(gate72inter8));
  nand2 gate850(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate851(.a(s_43), .b(gate72inter3), .O(gate72inter10));
  nor2  gate852(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate853(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate854(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1471(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1472(.a(gate73inter0), .b(s_132), .O(gate73inter1));
  and2  gate1473(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1474(.a(s_132), .O(gate73inter3));
  inv1  gate1475(.a(s_133), .O(gate73inter4));
  nand2 gate1476(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1477(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1478(.a(G1), .O(gate73inter7));
  inv1  gate1479(.a(G314), .O(gate73inter8));
  nand2 gate1480(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1481(.a(s_133), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1482(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1483(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1484(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate757(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate758(.a(gate76inter0), .b(s_30), .O(gate76inter1));
  and2  gate759(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate760(.a(s_30), .O(gate76inter3));
  inv1  gate761(.a(s_31), .O(gate76inter4));
  nand2 gate762(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate763(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate764(.a(G13), .O(gate76inter7));
  inv1  gate765(.a(G317), .O(gate76inter8));
  nand2 gate766(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate767(.a(s_31), .b(gate76inter3), .O(gate76inter10));
  nor2  gate768(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate769(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate770(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate2087(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2088(.a(gate77inter0), .b(s_220), .O(gate77inter1));
  and2  gate2089(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2090(.a(s_220), .O(gate77inter3));
  inv1  gate2091(.a(s_221), .O(gate77inter4));
  nand2 gate2092(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2093(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2094(.a(G2), .O(gate77inter7));
  inv1  gate2095(.a(G320), .O(gate77inter8));
  nand2 gate2096(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2097(.a(s_221), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2098(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2099(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2100(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1541(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1542(.a(gate79inter0), .b(s_142), .O(gate79inter1));
  and2  gate1543(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1544(.a(s_142), .O(gate79inter3));
  inv1  gate1545(.a(s_143), .O(gate79inter4));
  nand2 gate1546(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1547(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1548(.a(G10), .O(gate79inter7));
  inv1  gate1549(.a(G323), .O(gate79inter8));
  nand2 gate1550(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1551(.a(s_143), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1552(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1553(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1554(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate547(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate548(.a(gate91inter0), .b(s_0), .O(gate91inter1));
  and2  gate549(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate550(.a(s_0), .O(gate91inter3));
  inv1  gate551(.a(s_1), .O(gate91inter4));
  nand2 gate552(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate553(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate554(.a(G25), .O(gate91inter7));
  inv1  gate555(.a(G341), .O(gate91inter8));
  nand2 gate556(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate557(.a(s_1), .b(gate91inter3), .O(gate91inter10));
  nor2  gate558(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate559(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate560(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1009(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1010(.a(gate95inter0), .b(s_66), .O(gate95inter1));
  and2  gate1011(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1012(.a(s_66), .O(gate95inter3));
  inv1  gate1013(.a(s_67), .O(gate95inter4));
  nand2 gate1014(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1015(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1016(.a(G26), .O(gate95inter7));
  inv1  gate1017(.a(G347), .O(gate95inter8));
  nand2 gate1018(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1019(.a(s_67), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1020(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1021(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1022(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate981(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate982(.a(gate106inter0), .b(s_62), .O(gate106inter1));
  and2  gate983(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate984(.a(s_62), .O(gate106inter3));
  inv1  gate985(.a(s_63), .O(gate106inter4));
  nand2 gate986(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate987(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate988(.a(G364), .O(gate106inter7));
  inv1  gate989(.a(G365), .O(gate106inter8));
  nand2 gate990(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate991(.a(s_63), .b(gate106inter3), .O(gate106inter10));
  nor2  gate992(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate993(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate994(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1513(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1514(.a(gate108inter0), .b(s_138), .O(gate108inter1));
  and2  gate1515(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1516(.a(s_138), .O(gate108inter3));
  inv1  gate1517(.a(s_139), .O(gate108inter4));
  nand2 gate1518(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1519(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1520(.a(G368), .O(gate108inter7));
  inv1  gate1521(.a(G369), .O(gate108inter8));
  nand2 gate1522(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1523(.a(s_139), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1524(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1525(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1526(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1625(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1626(.a(gate109inter0), .b(s_154), .O(gate109inter1));
  and2  gate1627(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1628(.a(s_154), .O(gate109inter3));
  inv1  gate1629(.a(s_155), .O(gate109inter4));
  nand2 gate1630(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1631(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1632(.a(G370), .O(gate109inter7));
  inv1  gate1633(.a(G371), .O(gate109inter8));
  nand2 gate1634(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1635(.a(s_155), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1636(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1637(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1638(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate673(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate674(.a(gate116inter0), .b(s_18), .O(gate116inter1));
  and2  gate675(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate676(.a(s_18), .O(gate116inter3));
  inv1  gate677(.a(s_19), .O(gate116inter4));
  nand2 gate678(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate679(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate680(.a(G384), .O(gate116inter7));
  inv1  gate681(.a(G385), .O(gate116inter8));
  nand2 gate682(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate683(.a(s_19), .b(gate116inter3), .O(gate116inter10));
  nor2  gate684(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate685(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate686(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1751(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1752(.a(gate118inter0), .b(s_172), .O(gate118inter1));
  and2  gate1753(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1754(.a(s_172), .O(gate118inter3));
  inv1  gate1755(.a(s_173), .O(gate118inter4));
  nand2 gate1756(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1757(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1758(.a(G388), .O(gate118inter7));
  inv1  gate1759(.a(G389), .O(gate118inter8));
  nand2 gate1760(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1761(.a(s_173), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1762(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1763(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1764(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2143(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2144(.a(gate120inter0), .b(s_228), .O(gate120inter1));
  and2  gate2145(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2146(.a(s_228), .O(gate120inter3));
  inv1  gate2147(.a(s_229), .O(gate120inter4));
  nand2 gate2148(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2149(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2150(.a(G392), .O(gate120inter7));
  inv1  gate2151(.a(G393), .O(gate120inter8));
  nand2 gate2152(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2153(.a(s_229), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2154(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2155(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2156(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate561(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate562(.a(gate123inter0), .b(s_2), .O(gate123inter1));
  and2  gate563(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate564(.a(s_2), .O(gate123inter3));
  inv1  gate565(.a(s_3), .O(gate123inter4));
  nand2 gate566(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate567(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate568(.a(G398), .O(gate123inter7));
  inv1  gate569(.a(G399), .O(gate123inter8));
  nand2 gate570(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate571(.a(s_3), .b(gate123inter3), .O(gate123inter10));
  nor2  gate572(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate573(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate574(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1863(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1864(.a(gate124inter0), .b(s_188), .O(gate124inter1));
  and2  gate1865(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1866(.a(s_188), .O(gate124inter3));
  inv1  gate1867(.a(s_189), .O(gate124inter4));
  nand2 gate1868(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1869(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1870(.a(G400), .O(gate124inter7));
  inv1  gate1871(.a(G401), .O(gate124inter8));
  nand2 gate1872(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1873(.a(s_189), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1874(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1875(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1876(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2157(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2158(.a(gate126inter0), .b(s_230), .O(gate126inter1));
  and2  gate2159(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2160(.a(s_230), .O(gate126inter3));
  inv1  gate2161(.a(s_231), .O(gate126inter4));
  nand2 gate2162(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2163(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2164(.a(G404), .O(gate126inter7));
  inv1  gate2165(.a(G405), .O(gate126inter8));
  nand2 gate2166(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2167(.a(s_231), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2168(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2169(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2170(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate617(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate618(.a(gate127inter0), .b(s_10), .O(gate127inter1));
  and2  gate619(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate620(.a(s_10), .O(gate127inter3));
  inv1  gate621(.a(s_11), .O(gate127inter4));
  nand2 gate622(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate623(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate624(.a(G406), .O(gate127inter7));
  inv1  gate625(.a(G407), .O(gate127inter8));
  nand2 gate626(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate627(.a(s_11), .b(gate127inter3), .O(gate127inter10));
  nor2  gate628(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate629(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate630(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1653(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1654(.a(gate131inter0), .b(s_158), .O(gate131inter1));
  and2  gate1655(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1656(.a(s_158), .O(gate131inter3));
  inv1  gate1657(.a(s_159), .O(gate131inter4));
  nand2 gate1658(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1659(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1660(.a(G414), .O(gate131inter7));
  inv1  gate1661(.a(G415), .O(gate131inter8));
  nand2 gate1662(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1663(.a(s_159), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1664(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1665(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1666(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1569(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1570(.a(gate132inter0), .b(s_146), .O(gate132inter1));
  and2  gate1571(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1572(.a(s_146), .O(gate132inter3));
  inv1  gate1573(.a(s_147), .O(gate132inter4));
  nand2 gate1574(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1575(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1576(.a(G416), .O(gate132inter7));
  inv1  gate1577(.a(G417), .O(gate132inter8));
  nand2 gate1578(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1579(.a(s_147), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1580(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1581(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1582(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate785(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate786(.a(gate134inter0), .b(s_34), .O(gate134inter1));
  and2  gate787(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate788(.a(s_34), .O(gate134inter3));
  inv1  gate789(.a(s_35), .O(gate134inter4));
  nand2 gate790(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate791(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate792(.a(G420), .O(gate134inter7));
  inv1  gate793(.a(G421), .O(gate134inter8));
  nand2 gate794(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate795(.a(s_35), .b(gate134inter3), .O(gate134inter10));
  nor2  gate796(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate797(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate798(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate743(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate744(.a(gate137inter0), .b(s_28), .O(gate137inter1));
  and2  gate745(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate746(.a(s_28), .O(gate137inter3));
  inv1  gate747(.a(s_29), .O(gate137inter4));
  nand2 gate748(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate749(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate750(.a(G426), .O(gate137inter7));
  inv1  gate751(.a(G429), .O(gate137inter8));
  nand2 gate752(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate753(.a(s_29), .b(gate137inter3), .O(gate137inter10));
  nor2  gate754(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate755(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate756(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1415(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1416(.a(gate138inter0), .b(s_124), .O(gate138inter1));
  and2  gate1417(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1418(.a(s_124), .O(gate138inter3));
  inv1  gate1419(.a(s_125), .O(gate138inter4));
  nand2 gate1420(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1421(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1422(.a(G432), .O(gate138inter7));
  inv1  gate1423(.a(G435), .O(gate138inter8));
  nand2 gate1424(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1425(.a(s_125), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1426(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1427(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1428(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1667(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1668(.a(gate145inter0), .b(s_160), .O(gate145inter1));
  and2  gate1669(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1670(.a(s_160), .O(gate145inter3));
  inv1  gate1671(.a(s_161), .O(gate145inter4));
  nand2 gate1672(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1673(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1674(.a(G474), .O(gate145inter7));
  inv1  gate1675(.a(G477), .O(gate145inter8));
  nand2 gate1676(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1677(.a(s_161), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1678(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1679(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1680(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1037(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1038(.a(gate146inter0), .b(s_70), .O(gate146inter1));
  and2  gate1039(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1040(.a(s_70), .O(gate146inter3));
  inv1  gate1041(.a(s_71), .O(gate146inter4));
  nand2 gate1042(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1043(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1044(.a(G480), .O(gate146inter7));
  inv1  gate1045(.a(G483), .O(gate146inter8));
  nand2 gate1046(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1047(.a(s_71), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1048(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1049(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1050(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1877(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1878(.a(gate148inter0), .b(s_190), .O(gate148inter1));
  and2  gate1879(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1880(.a(s_190), .O(gate148inter3));
  inv1  gate1881(.a(s_191), .O(gate148inter4));
  nand2 gate1882(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1883(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1884(.a(G492), .O(gate148inter7));
  inv1  gate1885(.a(G495), .O(gate148inter8));
  nand2 gate1886(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1887(.a(s_191), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1888(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1889(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1890(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2213(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2214(.a(gate167inter0), .b(s_238), .O(gate167inter1));
  and2  gate2215(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2216(.a(s_238), .O(gate167inter3));
  inv1  gate2217(.a(s_239), .O(gate167inter4));
  nand2 gate2218(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2219(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2220(.a(G468), .O(gate167inter7));
  inv1  gate2221(.a(G543), .O(gate167inter8));
  nand2 gate2222(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2223(.a(s_239), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2224(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2225(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2226(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1989(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1990(.a(gate168inter0), .b(s_206), .O(gate168inter1));
  and2  gate1991(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1992(.a(s_206), .O(gate168inter3));
  inv1  gate1993(.a(s_207), .O(gate168inter4));
  nand2 gate1994(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1995(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1996(.a(G471), .O(gate168inter7));
  inv1  gate1997(.a(G543), .O(gate168inter8));
  nand2 gate1998(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1999(.a(s_207), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2000(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2001(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2002(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1849(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1850(.a(gate172inter0), .b(s_186), .O(gate172inter1));
  and2  gate1851(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1852(.a(s_186), .O(gate172inter3));
  inv1  gate1853(.a(s_187), .O(gate172inter4));
  nand2 gate1854(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1855(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1856(.a(G483), .O(gate172inter7));
  inv1  gate1857(.a(G549), .O(gate172inter8));
  nand2 gate1858(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1859(.a(s_187), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1860(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1861(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1862(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1681(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1682(.a(gate174inter0), .b(s_162), .O(gate174inter1));
  and2  gate1683(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1684(.a(s_162), .O(gate174inter3));
  inv1  gate1685(.a(s_163), .O(gate174inter4));
  nand2 gate1686(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1687(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1688(.a(G489), .O(gate174inter7));
  inv1  gate1689(.a(G552), .O(gate174inter8));
  nand2 gate1690(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1691(.a(s_163), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1692(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1693(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1694(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1765(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1766(.a(gate177inter0), .b(s_174), .O(gate177inter1));
  and2  gate1767(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1768(.a(s_174), .O(gate177inter3));
  inv1  gate1769(.a(s_175), .O(gate177inter4));
  nand2 gate1770(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1771(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1772(.a(G498), .O(gate177inter7));
  inv1  gate1773(.a(G558), .O(gate177inter8));
  nand2 gate1774(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1775(.a(s_175), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1776(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1777(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1778(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1443(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1444(.a(gate178inter0), .b(s_128), .O(gate178inter1));
  and2  gate1445(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1446(.a(s_128), .O(gate178inter3));
  inv1  gate1447(.a(s_129), .O(gate178inter4));
  nand2 gate1448(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1449(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1450(.a(G501), .O(gate178inter7));
  inv1  gate1451(.a(G558), .O(gate178inter8));
  nand2 gate1452(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1453(.a(s_129), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1454(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1455(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1456(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate715(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate716(.a(gate180inter0), .b(s_24), .O(gate180inter1));
  and2  gate717(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate718(.a(s_24), .O(gate180inter3));
  inv1  gate719(.a(s_25), .O(gate180inter4));
  nand2 gate720(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate721(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate722(.a(G507), .O(gate180inter7));
  inv1  gate723(.a(G561), .O(gate180inter8));
  nand2 gate724(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate725(.a(s_25), .b(gate180inter3), .O(gate180inter10));
  nor2  gate726(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate727(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate728(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate645(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate646(.a(gate182inter0), .b(s_14), .O(gate182inter1));
  and2  gate647(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate648(.a(s_14), .O(gate182inter3));
  inv1  gate649(.a(s_15), .O(gate182inter4));
  nand2 gate650(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate651(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate652(.a(G513), .O(gate182inter7));
  inv1  gate653(.a(G564), .O(gate182inter8));
  nand2 gate654(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate655(.a(s_15), .b(gate182inter3), .O(gate182inter10));
  nor2  gate656(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate657(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate658(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1163(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1164(.a(gate186inter0), .b(s_88), .O(gate186inter1));
  and2  gate1165(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1166(.a(s_88), .O(gate186inter3));
  inv1  gate1167(.a(s_89), .O(gate186inter4));
  nand2 gate1168(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1169(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1170(.a(G572), .O(gate186inter7));
  inv1  gate1171(.a(G573), .O(gate186inter8));
  nand2 gate1172(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1173(.a(s_89), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1174(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1175(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1176(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate701(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate702(.a(gate188inter0), .b(s_22), .O(gate188inter1));
  and2  gate703(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate704(.a(s_22), .O(gate188inter3));
  inv1  gate705(.a(s_23), .O(gate188inter4));
  nand2 gate706(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate707(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate708(.a(G576), .O(gate188inter7));
  inv1  gate709(.a(G577), .O(gate188inter8));
  nand2 gate710(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate711(.a(s_23), .b(gate188inter3), .O(gate188inter10));
  nor2  gate712(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate713(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate714(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1219(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1220(.a(gate189inter0), .b(s_96), .O(gate189inter1));
  and2  gate1221(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1222(.a(s_96), .O(gate189inter3));
  inv1  gate1223(.a(s_97), .O(gate189inter4));
  nand2 gate1224(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1225(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1226(.a(G578), .O(gate189inter7));
  inv1  gate1227(.a(G579), .O(gate189inter8));
  nand2 gate1228(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1229(.a(s_97), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1230(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1231(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1232(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate799(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate800(.a(gate193inter0), .b(s_36), .O(gate193inter1));
  and2  gate801(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate802(.a(s_36), .O(gate193inter3));
  inv1  gate803(.a(s_37), .O(gate193inter4));
  nand2 gate804(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate805(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate806(.a(G586), .O(gate193inter7));
  inv1  gate807(.a(G587), .O(gate193inter8));
  nand2 gate808(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate809(.a(s_37), .b(gate193inter3), .O(gate193inter10));
  nor2  gate810(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate811(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate812(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1247(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1248(.a(gate195inter0), .b(s_100), .O(gate195inter1));
  and2  gate1249(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1250(.a(s_100), .O(gate195inter3));
  inv1  gate1251(.a(s_101), .O(gate195inter4));
  nand2 gate1252(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1253(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1254(.a(G590), .O(gate195inter7));
  inv1  gate1255(.a(G591), .O(gate195inter8));
  nand2 gate1256(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1257(.a(s_101), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1258(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1259(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1260(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1499(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1500(.a(gate200inter0), .b(s_136), .O(gate200inter1));
  and2  gate1501(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1502(.a(s_136), .O(gate200inter3));
  inv1  gate1503(.a(s_137), .O(gate200inter4));
  nand2 gate1504(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1505(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1506(.a(G600), .O(gate200inter7));
  inv1  gate1507(.a(G601), .O(gate200inter8));
  nand2 gate1508(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1509(.a(s_137), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1510(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1511(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1512(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate883(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate884(.a(gate201inter0), .b(s_48), .O(gate201inter1));
  and2  gate885(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate886(.a(s_48), .O(gate201inter3));
  inv1  gate887(.a(s_49), .O(gate201inter4));
  nand2 gate888(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate889(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate890(.a(G602), .O(gate201inter7));
  inv1  gate891(.a(G607), .O(gate201inter8));
  nand2 gate892(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate893(.a(s_49), .b(gate201inter3), .O(gate201inter10));
  nor2  gate894(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate895(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate896(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate2199(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2200(.a(gate202inter0), .b(s_236), .O(gate202inter1));
  and2  gate2201(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2202(.a(s_236), .O(gate202inter3));
  inv1  gate2203(.a(s_237), .O(gate202inter4));
  nand2 gate2204(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2205(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2206(.a(G612), .O(gate202inter7));
  inv1  gate2207(.a(G617), .O(gate202inter8));
  nand2 gate2208(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2209(.a(s_237), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2210(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2211(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2212(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1121(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1122(.a(gate203inter0), .b(s_82), .O(gate203inter1));
  and2  gate1123(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1124(.a(s_82), .O(gate203inter3));
  inv1  gate1125(.a(s_83), .O(gate203inter4));
  nand2 gate1126(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1127(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1128(.a(G602), .O(gate203inter7));
  inv1  gate1129(.a(G612), .O(gate203inter8));
  nand2 gate1130(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1131(.a(s_83), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1132(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1133(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1134(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1737(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1738(.a(gate206inter0), .b(s_170), .O(gate206inter1));
  and2  gate1739(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1740(.a(s_170), .O(gate206inter3));
  inv1  gate1741(.a(s_171), .O(gate206inter4));
  nand2 gate1742(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1743(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1744(.a(G632), .O(gate206inter7));
  inv1  gate1745(.a(G637), .O(gate206inter8));
  nand2 gate1746(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1747(.a(s_171), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1748(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1749(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1750(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate813(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate814(.a(gate207inter0), .b(s_38), .O(gate207inter1));
  and2  gate815(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate816(.a(s_38), .O(gate207inter3));
  inv1  gate817(.a(s_39), .O(gate207inter4));
  nand2 gate818(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate819(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate820(.a(G622), .O(gate207inter7));
  inv1  gate821(.a(G632), .O(gate207inter8));
  nand2 gate822(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate823(.a(s_39), .b(gate207inter3), .O(gate207inter10));
  nor2  gate824(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate825(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate826(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1527(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1528(.a(gate208inter0), .b(s_140), .O(gate208inter1));
  and2  gate1529(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1530(.a(s_140), .O(gate208inter3));
  inv1  gate1531(.a(s_141), .O(gate208inter4));
  nand2 gate1532(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1533(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1534(.a(G627), .O(gate208inter7));
  inv1  gate1535(.a(G637), .O(gate208inter8));
  nand2 gate1536(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1537(.a(s_141), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1538(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1539(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1540(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1331(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1332(.a(gate209inter0), .b(s_112), .O(gate209inter1));
  and2  gate1333(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1334(.a(s_112), .O(gate209inter3));
  inv1  gate1335(.a(s_113), .O(gate209inter4));
  nand2 gate1336(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1337(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1338(.a(G602), .O(gate209inter7));
  inv1  gate1339(.a(G666), .O(gate209inter8));
  nand2 gate1340(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1341(.a(s_113), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1342(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1343(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1344(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1975(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1976(.a(gate214inter0), .b(s_204), .O(gate214inter1));
  and2  gate1977(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1978(.a(s_204), .O(gate214inter3));
  inv1  gate1979(.a(s_205), .O(gate214inter4));
  nand2 gate1980(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1981(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1982(.a(G612), .O(gate214inter7));
  inv1  gate1983(.a(G672), .O(gate214inter8));
  nand2 gate1984(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1985(.a(s_205), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1986(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1987(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1988(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1611(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1612(.a(gate221inter0), .b(s_152), .O(gate221inter1));
  and2  gate1613(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1614(.a(s_152), .O(gate221inter3));
  inv1  gate1615(.a(s_153), .O(gate221inter4));
  nand2 gate1616(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1617(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1618(.a(G622), .O(gate221inter7));
  inv1  gate1619(.a(G684), .O(gate221inter8));
  nand2 gate1620(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1621(.a(s_153), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1622(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1623(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1624(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1807(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1808(.a(gate224inter0), .b(s_180), .O(gate224inter1));
  and2  gate1809(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1810(.a(s_180), .O(gate224inter3));
  inv1  gate1811(.a(s_181), .O(gate224inter4));
  nand2 gate1812(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1813(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1814(.a(G637), .O(gate224inter7));
  inv1  gate1815(.a(G687), .O(gate224inter8));
  nand2 gate1816(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1817(.a(s_181), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1818(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1819(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1820(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate869(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate870(.a(gate225inter0), .b(s_46), .O(gate225inter1));
  and2  gate871(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate872(.a(s_46), .O(gate225inter3));
  inv1  gate873(.a(s_47), .O(gate225inter4));
  nand2 gate874(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate875(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate876(.a(G690), .O(gate225inter7));
  inv1  gate877(.a(G691), .O(gate225inter8));
  nand2 gate878(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate879(.a(s_47), .b(gate225inter3), .O(gate225inter10));
  nor2  gate880(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate881(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate882(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1709(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1710(.a(gate241inter0), .b(s_166), .O(gate241inter1));
  and2  gate1711(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1712(.a(s_166), .O(gate241inter3));
  inv1  gate1713(.a(s_167), .O(gate241inter4));
  nand2 gate1714(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1715(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1716(.a(G242), .O(gate241inter7));
  inv1  gate1717(.a(G730), .O(gate241inter8));
  nand2 gate1718(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1719(.a(s_167), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1720(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1721(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1722(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate687(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate688(.a(gate243inter0), .b(s_20), .O(gate243inter1));
  and2  gate689(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate690(.a(s_20), .O(gate243inter3));
  inv1  gate691(.a(s_21), .O(gate243inter4));
  nand2 gate692(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate693(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate694(.a(G245), .O(gate243inter7));
  inv1  gate695(.a(G733), .O(gate243inter8));
  nand2 gate696(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate697(.a(s_21), .b(gate243inter3), .O(gate243inter10));
  nor2  gate698(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate699(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate700(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate2059(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2060(.a(gate244inter0), .b(s_216), .O(gate244inter1));
  and2  gate2061(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2062(.a(s_216), .O(gate244inter3));
  inv1  gate2063(.a(s_217), .O(gate244inter4));
  nand2 gate2064(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2065(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2066(.a(G721), .O(gate244inter7));
  inv1  gate2067(.a(G733), .O(gate244inter8));
  nand2 gate2068(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2069(.a(s_217), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2070(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2071(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2072(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1317(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1318(.a(gate249inter0), .b(s_110), .O(gate249inter1));
  and2  gate1319(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1320(.a(s_110), .O(gate249inter3));
  inv1  gate1321(.a(s_111), .O(gate249inter4));
  nand2 gate1322(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1323(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1324(.a(G254), .O(gate249inter7));
  inv1  gate1325(.a(G742), .O(gate249inter8));
  nand2 gate1326(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1327(.a(s_111), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1328(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1329(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1330(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2031(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2032(.a(gate254inter0), .b(s_212), .O(gate254inter1));
  and2  gate2033(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2034(.a(s_212), .O(gate254inter3));
  inv1  gate2035(.a(s_213), .O(gate254inter4));
  nand2 gate2036(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2037(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2038(.a(G712), .O(gate254inter7));
  inv1  gate2039(.a(G748), .O(gate254inter8));
  nand2 gate2040(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2041(.a(s_213), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2042(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2043(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2044(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1233(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1234(.a(gate255inter0), .b(s_98), .O(gate255inter1));
  and2  gate1235(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1236(.a(s_98), .O(gate255inter3));
  inv1  gate1237(.a(s_99), .O(gate255inter4));
  nand2 gate1238(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1239(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1240(.a(G263), .O(gate255inter7));
  inv1  gate1241(.a(G751), .O(gate255inter8));
  nand2 gate1242(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1243(.a(s_99), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1244(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1245(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1246(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate855(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate856(.a(gate257inter0), .b(s_44), .O(gate257inter1));
  and2  gate857(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate858(.a(s_44), .O(gate257inter3));
  inv1  gate859(.a(s_45), .O(gate257inter4));
  nand2 gate860(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate861(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate862(.a(G754), .O(gate257inter7));
  inv1  gate863(.a(G755), .O(gate257inter8));
  nand2 gate864(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate865(.a(s_45), .b(gate257inter3), .O(gate257inter10));
  nor2  gate866(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate867(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate868(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1107(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1108(.a(gate259inter0), .b(s_80), .O(gate259inter1));
  and2  gate1109(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1110(.a(s_80), .O(gate259inter3));
  inv1  gate1111(.a(s_81), .O(gate259inter4));
  nand2 gate1112(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1113(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1114(.a(G758), .O(gate259inter7));
  inv1  gate1115(.a(G759), .O(gate259inter8));
  nand2 gate1116(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1117(.a(s_81), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1118(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1119(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1120(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1429(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1430(.a(gate261inter0), .b(s_126), .O(gate261inter1));
  and2  gate1431(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1432(.a(s_126), .O(gate261inter3));
  inv1  gate1433(.a(s_127), .O(gate261inter4));
  nand2 gate1434(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1435(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1436(.a(G762), .O(gate261inter7));
  inv1  gate1437(.a(G763), .O(gate261inter8));
  nand2 gate1438(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1439(.a(s_127), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1440(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1441(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1442(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1891(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1892(.a(gate267inter0), .b(s_192), .O(gate267inter1));
  and2  gate1893(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1894(.a(s_192), .O(gate267inter3));
  inv1  gate1895(.a(s_193), .O(gate267inter4));
  nand2 gate1896(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1897(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1898(.a(G648), .O(gate267inter7));
  inv1  gate1899(.a(G776), .O(gate267inter8));
  nand2 gate1900(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1901(.a(s_193), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1902(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1903(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1904(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1191(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1192(.a(gate271inter0), .b(s_92), .O(gate271inter1));
  and2  gate1193(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1194(.a(s_92), .O(gate271inter3));
  inv1  gate1195(.a(s_93), .O(gate271inter4));
  nand2 gate1196(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1197(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1198(.a(G660), .O(gate271inter7));
  inv1  gate1199(.a(G788), .O(gate271inter8));
  nand2 gate1200(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1201(.a(s_93), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1202(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1203(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1204(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1821(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1822(.a(gate276inter0), .b(s_182), .O(gate276inter1));
  and2  gate1823(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1824(.a(s_182), .O(gate276inter3));
  inv1  gate1825(.a(s_183), .O(gate276inter4));
  nand2 gate1826(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1827(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1828(.a(G773), .O(gate276inter7));
  inv1  gate1829(.a(G797), .O(gate276inter8));
  nand2 gate1830(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1831(.a(s_183), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1832(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1833(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1834(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate771(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate772(.a(gate277inter0), .b(s_32), .O(gate277inter1));
  and2  gate773(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate774(.a(s_32), .O(gate277inter3));
  inv1  gate775(.a(s_33), .O(gate277inter4));
  nand2 gate776(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate777(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate778(.a(G648), .O(gate277inter7));
  inv1  gate779(.a(G800), .O(gate277inter8));
  nand2 gate780(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate781(.a(s_33), .b(gate277inter3), .O(gate277inter10));
  nor2  gate782(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate783(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate784(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1205(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1206(.a(gate279inter0), .b(s_94), .O(gate279inter1));
  and2  gate1207(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1208(.a(s_94), .O(gate279inter3));
  inv1  gate1209(.a(s_95), .O(gate279inter4));
  nand2 gate1210(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1211(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1212(.a(G651), .O(gate279inter7));
  inv1  gate1213(.a(G803), .O(gate279inter8));
  nand2 gate1214(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1215(.a(s_95), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1216(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1217(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1218(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2017(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2018(.a(gate283inter0), .b(s_210), .O(gate283inter1));
  and2  gate2019(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2020(.a(s_210), .O(gate283inter3));
  inv1  gate2021(.a(s_211), .O(gate283inter4));
  nand2 gate2022(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2023(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2024(.a(G657), .O(gate283inter7));
  inv1  gate2025(.a(G809), .O(gate283inter8));
  nand2 gate2026(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2027(.a(s_211), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2028(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2029(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2030(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2129(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2130(.a(gate288inter0), .b(s_226), .O(gate288inter1));
  and2  gate2131(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2132(.a(s_226), .O(gate288inter3));
  inv1  gate2133(.a(s_227), .O(gate288inter4));
  nand2 gate2134(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2135(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2136(.a(G791), .O(gate288inter7));
  inv1  gate2137(.a(G815), .O(gate288inter8));
  nand2 gate2138(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2139(.a(s_227), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2140(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2141(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2142(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1359(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1360(.a(gate289inter0), .b(s_116), .O(gate289inter1));
  and2  gate1361(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1362(.a(s_116), .O(gate289inter3));
  inv1  gate1363(.a(s_117), .O(gate289inter4));
  nand2 gate1364(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1365(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1366(.a(G818), .O(gate289inter7));
  inv1  gate1367(.a(G819), .O(gate289inter8));
  nand2 gate1368(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1369(.a(s_117), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1370(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1371(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1372(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate631(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate632(.a(gate291inter0), .b(s_12), .O(gate291inter1));
  and2  gate633(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate634(.a(s_12), .O(gate291inter3));
  inv1  gate635(.a(s_13), .O(gate291inter4));
  nand2 gate636(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate637(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate638(.a(G822), .O(gate291inter7));
  inv1  gate639(.a(G823), .O(gate291inter8));
  nand2 gate640(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate641(.a(s_13), .b(gate291inter3), .O(gate291inter10));
  nor2  gate642(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate643(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate644(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate967(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate968(.a(gate293inter0), .b(s_60), .O(gate293inter1));
  and2  gate969(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate970(.a(s_60), .O(gate293inter3));
  inv1  gate971(.a(s_61), .O(gate293inter4));
  nand2 gate972(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate973(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate974(.a(G828), .O(gate293inter7));
  inv1  gate975(.a(G829), .O(gate293inter8));
  nand2 gate976(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate977(.a(s_61), .b(gate293inter3), .O(gate293inter10));
  nor2  gate978(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate979(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate980(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate589(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate590(.a(gate295inter0), .b(s_6), .O(gate295inter1));
  and2  gate591(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate592(.a(s_6), .O(gate295inter3));
  inv1  gate593(.a(s_7), .O(gate295inter4));
  nand2 gate594(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate595(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate596(.a(G830), .O(gate295inter7));
  inv1  gate597(.a(G831), .O(gate295inter8));
  nand2 gate598(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate599(.a(s_7), .b(gate295inter3), .O(gate295inter10));
  nor2  gate600(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate601(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate602(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1261(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1262(.a(gate391inter0), .b(s_102), .O(gate391inter1));
  and2  gate1263(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1264(.a(s_102), .O(gate391inter3));
  inv1  gate1265(.a(s_103), .O(gate391inter4));
  nand2 gate1266(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1267(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1268(.a(G5), .O(gate391inter7));
  inv1  gate1269(.a(G1048), .O(gate391inter8));
  nand2 gate1270(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1271(.a(s_103), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1272(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1273(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1274(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate575(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate576(.a(gate395inter0), .b(s_4), .O(gate395inter1));
  and2  gate577(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate578(.a(s_4), .O(gate395inter3));
  inv1  gate579(.a(s_5), .O(gate395inter4));
  nand2 gate580(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate581(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate582(.a(G9), .O(gate395inter7));
  inv1  gate583(.a(G1060), .O(gate395inter8));
  nand2 gate584(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate585(.a(s_5), .b(gate395inter3), .O(gate395inter10));
  nor2  gate586(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate587(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate588(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2073(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2074(.a(gate402inter0), .b(s_218), .O(gate402inter1));
  and2  gate2075(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2076(.a(s_218), .O(gate402inter3));
  inv1  gate2077(.a(s_219), .O(gate402inter4));
  nand2 gate2078(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2079(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2080(.a(G16), .O(gate402inter7));
  inv1  gate2081(.a(G1081), .O(gate402inter8));
  nand2 gate2082(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2083(.a(s_219), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2084(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2085(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2086(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1023(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1024(.a(gate405inter0), .b(s_68), .O(gate405inter1));
  and2  gate1025(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1026(.a(s_68), .O(gate405inter3));
  inv1  gate1027(.a(s_69), .O(gate405inter4));
  nand2 gate1028(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1029(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1030(.a(G19), .O(gate405inter7));
  inv1  gate1031(.a(G1090), .O(gate405inter8));
  nand2 gate1032(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1033(.a(s_69), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1034(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1035(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1036(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1933(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1934(.a(gate407inter0), .b(s_198), .O(gate407inter1));
  and2  gate1935(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1936(.a(s_198), .O(gate407inter3));
  inv1  gate1937(.a(s_199), .O(gate407inter4));
  nand2 gate1938(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1939(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1940(.a(G21), .O(gate407inter7));
  inv1  gate1941(.a(G1096), .O(gate407inter8));
  nand2 gate1942(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1943(.a(s_199), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1944(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1945(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1946(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate897(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate898(.a(gate411inter0), .b(s_50), .O(gate411inter1));
  and2  gate899(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate900(.a(s_50), .O(gate411inter3));
  inv1  gate901(.a(s_51), .O(gate411inter4));
  nand2 gate902(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate903(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate904(.a(G25), .O(gate411inter7));
  inv1  gate905(.a(G1108), .O(gate411inter8));
  nand2 gate906(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate907(.a(s_51), .b(gate411inter3), .O(gate411inter10));
  nor2  gate908(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate909(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate910(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1401(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1402(.a(gate414inter0), .b(s_122), .O(gate414inter1));
  and2  gate1403(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1404(.a(s_122), .O(gate414inter3));
  inv1  gate1405(.a(s_123), .O(gate414inter4));
  nand2 gate1406(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1407(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1408(.a(G28), .O(gate414inter7));
  inv1  gate1409(.a(G1117), .O(gate414inter8));
  nand2 gate1410(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1411(.a(s_123), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1412(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1413(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1414(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2045(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2046(.a(gate420inter0), .b(s_214), .O(gate420inter1));
  and2  gate2047(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2048(.a(s_214), .O(gate420inter3));
  inv1  gate2049(.a(s_215), .O(gate420inter4));
  nand2 gate2050(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2051(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2052(.a(G1036), .O(gate420inter7));
  inv1  gate2053(.a(G1132), .O(gate420inter8));
  nand2 gate2054(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2055(.a(s_215), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2056(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2057(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2058(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1793(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1794(.a(gate427inter0), .b(s_178), .O(gate427inter1));
  and2  gate1795(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1796(.a(s_178), .O(gate427inter3));
  inv1  gate1797(.a(s_179), .O(gate427inter4));
  nand2 gate1798(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1799(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1800(.a(G5), .O(gate427inter7));
  inv1  gate1801(.a(G1144), .O(gate427inter8));
  nand2 gate1802(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1803(.a(s_179), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1804(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1805(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1806(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1723(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1724(.a(gate428inter0), .b(s_168), .O(gate428inter1));
  and2  gate1725(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1726(.a(s_168), .O(gate428inter3));
  inv1  gate1727(.a(s_169), .O(gate428inter4));
  nand2 gate1728(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1729(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1730(.a(G1048), .O(gate428inter7));
  inv1  gate1731(.a(G1144), .O(gate428inter8));
  nand2 gate1732(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1733(.a(s_169), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1734(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1735(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1736(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1065(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1066(.a(gate431inter0), .b(s_74), .O(gate431inter1));
  and2  gate1067(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1068(.a(s_74), .O(gate431inter3));
  inv1  gate1069(.a(s_75), .O(gate431inter4));
  nand2 gate1070(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1071(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1072(.a(G7), .O(gate431inter7));
  inv1  gate1073(.a(G1150), .O(gate431inter8));
  nand2 gate1074(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1075(.a(s_75), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1076(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1077(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1078(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1485(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1486(.a(gate440inter0), .b(s_134), .O(gate440inter1));
  and2  gate1487(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1488(.a(s_134), .O(gate440inter3));
  inv1  gate1489(.a(s_135), .O(gate440inter4));
  nand2 gate1490(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1491(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1492(.a(G1066), .O(gate440inter7));
  inv1  gate1493(.a(G1162), .O(gate440inter8));
  nand2 gate1494(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1495(.a(s_135), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1496(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1497(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1498(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate659(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate660(.a(gate441inter0), .b(s_16), .O(gate441inter1));
  and2  gate661(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate662(.a(s_16), .O(gate441inter3));
  inv1  gate663(.a(s_17), .O(gate441inter4));
  nand2 gate664(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate665(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate666(.a(G12), .O(gate441inter7));
  inv1  gate667(.a(G1165), .O(gate441inter8));
  nand2 gate668(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate669(.a(s_17), .b(gate441inter3), .O(gate441inter10));
  nor2  gate670(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate671(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate672(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1177(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1178(.a(gate444inter0), .b(s_90), .O(gate444inter1));
  and2  gate1179(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1180(.a(s_90), .O(gate444inter3));
  inv1  gate1181(.a(s_91), .O(gate444inter4));
  nand2 gate1182(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1183(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1184(.a(G1072), .O(gate444inter7));
  inv1  gate1185(.a(G1168), .O(gate444inter8));
  nand2 gate1186(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1187(.a(s_91), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1188(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1189(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1190(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2115(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2116(.a(gate450inter0), .b(s_224), .O(gate450inter1));
  and2  gate2117(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2118(.a(s_224), .O(gate450inter3));
  inv1  gate2119(.a(s_225), .O(gate450inter4));
  nand2 gate2120(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2121(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2122(.a(G1081), .O(gate450inter7));
  inv1  gate2123(.a(G1177), .O(gate450inter8));
  nand2 gate2124(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2125(.a(s_225), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2126(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2127(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2128(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2101(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2102(.a(gate458inter0), .b(s_222), .O(gate458inter1));
  and2  gate2103(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2104(.a(s_222), .O(gate458inter3));
  inv1  gate2105(.a(s_223), .O(gate458inter4));
  nand2 gate2106(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2107(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2108(.a(G1093), .O(gate458inter7));
  inv1  gate2109(.a(G1189), .O(gate458inter8));
  nand2 gate2110(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2111(.a(s_223), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2112(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2113(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2114(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1905(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1906(.a(gate462inter0), .b(s_194), .O(gate462inter1));
  and2  gate1907(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1908(.a(s_194), .O(gate462inter3));
  inv1  gate1909(.a(s_195), .O(gate462inter4));
  nand2 gate1910(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1911(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1912(.a(G1099), .O(gate462inter7));
  inv1  gate1913(.a(G1195), .O(gate462inter8));
  nand2 gate1914(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1915(.a(s_195), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1916(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1917(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1918(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2227(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2228(.a(gate464inter0), .b(s_240), .O(gate464inter1));
  and2  gate2229(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2230(.a(s_240), .O(gate464inter3));
  inv1  gate2231(.a(s_241), .O(gate464inter4));
  nand2 gate2232(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2233(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2234(.a(G1102), .O(gate464inter7));
  inv1  gate2235(.a(G1198), .O(gate464inter8));
  nand2 gate2236(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2237(.a(s_241), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2238(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2239(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2240(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1597(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1598(.a(gate465inter0), .b(s_150), .O(gate465inter1));
  and2  gate1599(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1600(.a(s_150), .O(gate465inter3));
  inv1  gate1601(.a(s_151), .O(gate465inter4));
  nand2 gate1602(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1603(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1604(.a(G24), .O(gate465inter7));
  inv1  gate1605(.a(G1201), .O(gate465inter8));
  nand2 gate1606(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1607(.a(s_151), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1608(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1609(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1610(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1149(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1150(.a(gate466inter0), .b(s_86), .O(gate466inter1));
  and2  gate1151(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1152(.a(s_86), .O(gate466inter3));
  inv1  gate1153(.a(s_87), .O(gate466inter4));
  nand2 gate1154(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1155(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1156(.a(G1105), .O(gate466inter7));
  inv1  gate1157(.a(G1201), .O(gate466inter8));
  nand2 gate1158(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1159(.a(s_87), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1160(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1161(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1162(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1275(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1276(.a(gate468inter0), .b(s_104), .O(gate468inter1));
  and2  gate1277(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1278(.a(s_104), .O(gate468inter3));
  inv1  gate1279(.a(s_105), .O(gate468inter4));
  nand2 gate1280(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1281(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1282(.a(G1108), .O(gate468inter7));
  inv1  gate1283(.a(G1204), .O(gate468inter8));
  nand2 gate1284(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1285(.a(s_105), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1286(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1287(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1288(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate911(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate912(.a(gate471inter0), .b(s_52), .O(gate471inter1));
  and2  gate913(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate914(.a(s_52), .O(gate471inter3));
  inv1  gate915(.a(s_53), .O(gate471inter4));
  nand2 gate916(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate917(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate918(.a(G27), .O(gate471inter7));
  inv1  gate919(.a(G1210), .O(gate471inter8));
  nand2 gate920(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate921(.a(s_53), .b(gate471inter3), .O(gate471inter10));
  nor2  gate922(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate923(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate924(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1079(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1080(.a(gate479inter0), .b(s_76), .O(gate479inter1));
  and2  gate1081(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1082(.a(s_76), .O(gate479inter3));
  inv1  gate1083(.a(s_77), .O(gate479inter4));
  nand2 gate1084(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1085(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1086(.a(G31), .O(gate479inter7));
  inv1  gate1087(.a(G1222), .O(gate479inter8));
  nand2 gate1088(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1089(.a(s_77), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1090(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1091(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1092(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate995(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate996(.a(gate481inter0), .b(s_64), .O(gate481inter1));
  and2  gate997(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate998(.a(s_64), .O(gate481inter3));
  inv1  gate999(.a(s_65), .O(gate481inter4));
  nand2 gate1000(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1001(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1002(.a(G32), .O(gate481inter7));
  inv1  gate1003(.a(G1225), .O(gate481inter8));
  nand2 gate1004(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1005(.a(s_65), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1006(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1007(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1008(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate953(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate954(.a(gate483inter0), .b(s_58), .O(gate483inter1));
  and2  gate955(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate956(.a(s_58), .O(gate483inter3));
  inv1  gate957(.a(s_59), .O(gate483inter4));
  nand2 gate958(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate959(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate960(.a(G1228), .O(gate483inter7));
  inv1  gate961(.a(G1229), .O(gate483inter8));
  nand2 gate962(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate963(.a(s_59), .b(gate483inter3), .O(gate483inter10));
  nor2  gate964(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate965(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate966(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1695(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1696(.a(gate486inter0), .b(s_164), .O(gate486inter1));
  and2  gate1697(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1698(.a(s_164), .O(gate486inter3));
  inv1  gate1699(.a(s_165), .O(gate486inter4));
  nand2 gate1700(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1701(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1702(.a(G1234), .O(gate486inter7));
  inv1  gate1703(.a(G1235), .O(gate486inter8));
  nand2 gate1704(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1705(.a(s_165), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1706(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1707(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1708(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1639(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1640(.a(gate487inter0), .b(s_156), .O(gate487inter1));
  and2  gate1641(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1642(.a(s_156), .O(gate487inter3));
  inv1  gate1643(.a(s_157), .O(gate487inter4));
  nand2 gate1644(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1645(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1646(.a(G1236), .O(gate487inter7));
  inv1  gate1647(.a(G1237), .O(gate487inter8));
  nand2 gate1648(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1649(.a(s_157), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1650(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1651(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1652(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1919(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1920(.a(gate490inter0), .b(s_196), .O(gate490inter1));
  and2  gate1921(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1922(.a(s_196), .O(gate490inter3));
  inv1  gate1923(.a(s_197), .O(gate490inter4));
  nand2 gate1924(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1925(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1926(.a(G1242), .O(gate490inter7));
  inv1  gate1927(.a(G1243), .O(gate490inter8));
  nand2 gate1928(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1929(.a(s_197), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1930(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1931(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1932(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1093(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1094(.a(gate492inter0), .b(s_78), .O(gate492inter1));
  and2  gate1095(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1096(.a(s_78), .O(gate492inter3));
  inv1  gate1097(.a(s_79), .O(gate492inter4));
  nand2 gate1098(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1099(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1100(.a(G1246), .O(gate492inter7));
  inv1  gate1101(.a(G1247), .O(gate492inter8));
  nand2 gate1102(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1103(.a(s_79), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1104(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1105(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1106(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1289(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1290(.a(gate494inter0), .b(s_106), .O(gate494inter1));
  and2  gate1291(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1292(.a(s_106), .O(gate494inter3));
  inv1  gate1293(.a(s_107), .O(gate494inter4));
  nand2 gate1294(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1295(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1296(.a(G1250), .O(gate494inter7));
  inv1  gate1297(.a(G1251), .O(gate494inter8));
  nand2 gate1298(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1299(.a(s_107), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1300(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1301(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1302(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1457(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1458(.a(gate496inter0), .b(s_130), .O(gate496inter1));
  and2  gate1459(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1460(.a(s_130), .O(gate496inter3));
  inv1  gate1461(.a(s_131), .O(gate496inter4));
  nand2 gate1462(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1463(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1464(.a(G1254), .O(gate496inter7));
  inv1  gate1465(.a(G1255), .O(gate496inter8));
  nand2 gate1466(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1467(.a(s_131), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1468(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1469(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1470(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2185(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2186(.a(gate502inter0), .b(s_234), .O(gate502inter1));
  and2  gate2187(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2188(.a(s_234), .O(gate502inter3));
  inv1  gate2189(.a(s_235), .O(gate502inter4));
  nand2 gate2190(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2191(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2192(.a(G1266), .O(gate502inter7));
  inv1  gate2193(.a(G1267), .O(gate502inter8));
  nand2 gate2194(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2195(.a(s_235), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2196(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2197(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2198(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate603(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate604(.a(gate508inter0), .b(s_8), .O(gate508inter1));
  and2  gate605(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate606(.a(s_8), .O(gate508inter3));
  inv1  gate607(.a(s_9), .O(gate508inter4));
  nand2 gate608(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate609(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate610(.a(G1278), .O(gate508inter7));
  inv1  gate611(.a(G1279), .O(gate508inter8));
  nand2 gate612(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate613(.a(s_9), .b(gate508inter3), .O(gate508inter10));
  nor2  gate614(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate615(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate616(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2003(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2004(.a(gate509inter0), .b(s_208), .O(gate509inter1));
  and2  gate2005(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2006(.a(s_208), .O(gate509inter3));
  inv1  gate2007(.a(s_209), .O(gate509inter4));
  nand2 gate2008(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2009(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2010(.a(G1280), .O(gate509inter7));
  inv1  gate2011(.a(G1281), .O(gate509inter8));
  nand2 gate2012(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2013(.a(s_209), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2014(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2015(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2016(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1135(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1136(.a(gate511inter0), .b(s_84), .O(gate511inter1));
  and2  gate1137(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1138(.a(s_84), .O(gate511inter3));
  inv1  gate1139(.a(s_85), .O(gate511inter4));
  nand2 gate1140(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1141(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1142(.a(G1284), .O(gate511inter7));
  inv1  gate1143(.a(G1285), .O(gate511inter8));
  nand2 gate1144(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1145(.a(s_85), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1146(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1147(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1148(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1051(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1052(.a(gate514inter0), .b(s_72), .O(gate514inter1));
  and2  gate1053(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1054(.a(s_72), .O(gate514inter3));
  inv1  gate1055(.a(s_73), .O(gate514inter4));
  nand2 gate1056(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1057(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1058(.a(G1290), .O(gate514inter7));
  inv1  gate1059(.a(G1291), .O(gate514inter8));
  nand2 gate1060(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1061(.a(s_73), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1062(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1063(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1064(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule