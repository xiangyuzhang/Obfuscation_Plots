module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1891(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1892(.a(gate9inter0), .b(s_192), .O(gate9inter1));
  and2  gate1893(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1894(.a(s_192), .O(gate9inter3));
  inv1  gate1895(.a(s_193), .O(gate9inter4));
  nand2 gate1896(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1897(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1898(.a(G1), .O(gate9inter7));
  inv1  gate1899(.a(G2), .O(gate9inter8));
  nand2 gate1900(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1901(.a(s_193), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1902(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1903(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1904(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2045(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2046(.a(gate11inter0), .b(s_214), .O(gate11inter1));
  and2  gate2047(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2048(.a(s_214), .O(gate11inter3));
  inv1  gate2049(.a(s_215), .O(gate11inter4));
  nand2 gate2050(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2051(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2052(.a(G5), .O(gate11inter7));
  inv1  gate2053(.a(G6), .O(gate11inter8));
  nand2 gate2054(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2055(.a(s_215), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2056(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2057(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2058(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate645(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate646(.a(gate15inter0), .b(s_14), .O(gate15inter1));
  and2  gate647(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate648(.a(s_14), .O(gate15inter3));
  inv1  gate649(.a(s_15), .O(gate15inter4));
  nand2 gate650(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate651(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate652(.a(G13), .O(gate15inter7));
  inv1  gate653(.a(G14), .O(gate15inter8));
  nand2 gate654(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate655(.a(s_15), .b(gate15inter3), .O(gate15inter10));
  nor2  gate656(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate657(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate658(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate631(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate632(.a(gate16inter0), .b(s_12), .O(gate16inter1));
  and2  gate633(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate634(.a(s_12), .O(gate16inter3));
  inv1  gate635(.a(s_13), .O(gate16inter4));
  nand2 gate636(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate637(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate638(.a(G15), .O(gate16inter7));
  inv1  gate639(.a(G16), .O(gate16inter8));
  nand2 gate640(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate641(.a(s_13), .b(gate16inter3), .O(gate16inter10));
  nor2  gate642(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate643(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate644(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2409(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2410(.a(gate17inter0), .b(s_266), .O(gate17inter1));
  and2  gate2411(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2412(.a(s_266), .O(gate17inter3));
  inv1  gate2413(.a(s_267), .O(gate17inter4));
  nand2 gate2414(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2415(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2416(.a(G17), .O(gate17inter7));
  inv1  gate2417(.a(G18), .O(gate17inter8));
  nand2 gate2418(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2419(.a(s_267), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2420(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2421(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2422(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate3123(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate3124(.a(gate18inter0), .b(s_368), .O(gate18inter1));
  and2  gate3125(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate3126(.a(s_368), .O(gate18inter3));
  inv1  gate3127(.a(s_369), .O(gate18inter4));
  nand2 gate3128(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate3129(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate3130(.a(G19), .O(gate18inter7));
  inv1  gate3131(.a(G20), .O(gate18inter8));
  nand2 gate3132(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate3133(.a(s_369), .b(gate18inter3), .O(gate18inter10));
  nor2  gate3134(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate3135(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate3136(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1051(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1052(.a(gate21inter0), .b(s_72), .O(gate21inter1));
  and2  gate1053(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1054(.a(s_72), .O(gate21inter3));
  inv1  gate1055(.a(s_73), .O(gate21inter4));
  nand2 gate1056(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1057(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1058(.a(G25), .O(gate21inter7));
  inv1  gate1059(.a(G26), .O(gate21inter8));
  nand2 gate1060(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1061(.a(s_73), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1062(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1063(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1064(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1443(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1444(.a(gate23inter0), .b(s_128), .O(gate23inter1));
  and2  gate1445(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1446(.a(s_128), .O(gate23inter3));
  inv1  gate1447(.a(s_129), .O(gate23inter4));
  nand2 gate1448(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1449(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1450(.a(G29), .O(gate23inter7));
  inv1  gate1451(.a(G30), .O(gate23inter8));
  nand2 gate1452(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1453(.a(s_129), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1454(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1455(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1456(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1107(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1108(.a(gate24inter0), .b(s_80), .O(gate24inter1));
  and2  gate1109(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1110(.a(s_80), .O(gate24inter3));
  inv1  gate1111(.a(s_81), .O(gate24inter4));
  nand2 gate1112(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1113(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1114(.a(G31), .O(gate24inter7));
  inv1  gate1115(.a(G32), .O(gate24inter8));
  nand2 gate1116(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1117(.a(s_81), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1118(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1119(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1120(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1863(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1864(.a(gate26inter0), .b(s_188), .O(gate26inter1));
  and2  gate1865(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1866(.a(s_188), .O(gate26inter3));
  inv1  gate1867(.a(s_189), .O(gate26inter4));
  nand2 gate1868(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1869(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1870(.a(G9), .O(gate26inter7));
  inv1  gate1871(.a(G13), .O(gate26inter8));
  nand2 gate1872(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1873(.a(s_189), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1874(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1875(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1876(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate673(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate674(.a(gate27inter0), .b(s_18), .O(gate27inter1));
  and2  gate675(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate676(.a(s_18), .O(gate27inter3));
  inv1  gate677(.a(s_19), .O(gate27inter4));
  nand2 gate678(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate679(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate680(.a(G2), .O(gate27inter7));
  inv1  gate681(.a(G6), .O(gate27inter8));
  nand2 gate682(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate683(.a(s_19), .b(gate27inter3), .O(gate27inter10));
  nor2  gate684(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate685(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate686(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate2773(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2774(.a(gate28inter0), .b(s_318), .O(gate28inter1));
  and2  gate2775(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2776(.a(s_318), .O(gate28inter3));
  inv1  gate2777(.a(s_319), .O(gate28inter4));
  nand2 gate2778(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2779(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2780(.a(G10), .O(gate28inter7));
  inv1  gate2781(.a(G14), .O(gate28inter8));
  nand2 gate2782(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2783(.a(s_319), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2784(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2785(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2786(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate2647(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2648(.a(gate30inter0), .b(s_300), .O(gate30inter1));
  and2  gate2649(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2650(.a(s_300), .O(gate30inter3));
  inv1  gate2651(.a(s_301), .O(gate30inter4));
  nand2 gate2652(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2653(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2654(.a(G11), .O(gate30inter7));
  inv1  gate2655(.a(G15), .O(gate30inter8));
  nand2 gate2656(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2657(.a(s_301), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2658(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2659(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2660(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2969(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2970(.a(gate36inter0), .b(s_346), .O(gate36inter1));
  and2  gate2971(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2972(.a(s_346), .O(gate36inter3));
  inv1  gate2973(.a(s_347), .O(gate36inter4));
  nand2 gate2974(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2975(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2976(.a(G26), .O(gate36inter7));
  inv1  gate2977(.a(G30), .O(gate36inter8));
  nand2 gate2978(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2979(.a(s_347), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2980(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2981(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2982(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1695(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1696(.a(gate40inter0), .b(s_164), .O(gate40inter1));
  and2  gate1697(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1698(.a(s_164), .O(gate40inter3));
  inv1  gate1699(.a(s_165), .O(gate40inter4));
  nand2 gate1700(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1701(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1702(.a(G28), .O(gate40inter7));
  inv1  gate1703(.a(G32), .O(gate40inter8));
  nand2 gate1704(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1705(.a(s_165), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1706(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1707(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1708(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1765(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1766(.a(gate41inter0), .b(s_174), .O(gate41inter1));
  and2  gate1767(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1768(.a(s_174), .O(gate41inter3));
  inv1  gate1769(.a(s_175), .O(gate41inter4));
  nand2 gate1770(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1771(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1772(.a(G1), .O(gate41inter7));
  inv1  gate1773(.a(G266), .O(gate41inter8));
  nand2 gate1774(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1775(.a(s_175), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1776(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1777(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1778(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2661(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2662(.a(gate42inter0), .b(s_302), .O(gate42inter1));
  and2  gate2663(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2664(.a(s_302), .O(gate42inter3));
  inv1  gate2665(.a(s_303), .O(gate42inter4));
  nand2 gate2666(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2667(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2668(.a(G2), .O(gate42inter7));
  inv1  gate2669(.a(G266), .O(gate42inter8));
  nand2 gate2670(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2671(.a(s_303), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2672(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2673(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2674(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2731(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2732(.a(gate46inter0), .b(s_312), .O(gate46inter1));
  and2  gate2733(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2734(.a(s_312), .O(gate46inter3));
  inv1  gate2735(.a(s_313), .O(gate46inter4));
  nand2 gate2736(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2737(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2738(.a(G6), .O(gate46inter7));
  inv1  gate2739(.a(G272), .O(gate46inter8));
  nand2 gate2740(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2741(.a(s_313), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2742(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2743(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2744(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate855(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate856(.a(gate48inter0), .b(s_44), .O(gate48inter1));
  and2  gate857(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate858(.a(s_44), .O(gate48inter3));
  inv1  gate859(.a(s_45), .O(gate48inter4));
  nand2 gate860(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate861(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate862(.a(G8), .O(gate48inter7));
  inv1  gate863(.a(G275), .O(gate48inter8));
  nand2 gate864(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate865(.a(s_45), .b(gate48inter3), .O(gate48inter10));
  nor2  gate866(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate867(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate868(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2143(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2144(.a(gate49inter0), .b(s_228), .O(gate49inter1));
  and2  gate2145(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2146(.a(s_228), .O(gate49inter3));
  inv1  gate2147(.a(s_229), .O(gate49inter4));
  nand2 gate2148(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2149(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2150(.a(G9), .O(gate49inter7));
  inv1  gate2151(.a(G278), .O(gate49inter8));
  nand2 gate2152(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2153(.a(s_229), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2154(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2155(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2156(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1359(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1360(.a(gate50inter0), .b(s_116), .O(gate50inter1));
  and2  gate1361(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1362(.a(s_116), .O(gate50inter3));
  inv1  gate1363(.a(s_117), .O(gate50inter4));
  nand2 gate1364(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1365(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1366(.a(G10), .O(gate50inter7));
  inv1  gate1367(.a(G278), .O(gate50inter8));
  nand2 gate1368(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1369(.a(s_117), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1370(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1371(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1372(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2843(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2844(.a(gate51inter0), .b(s_328), .O(gate51inter1));
  and2  gate2845(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2846(.a(s_328), .O(gate51inter3));
  inv1  gate2847(.a(s_329), .O(gate51inter4));
  nand2 gate2848(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2849(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2850(.a(G11), .O(gate51inter7));
  inv1  gate2851(.a(G281), .O(gate51inter8));
  nand2 gate2852(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2853(.a(s_329), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2854(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2855(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2856(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2451(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2452(.a(gate53inter0), .b(s_272), .O(gate53inter1));
  and2  gate2453(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2454(.a(s_272), .O(gate53inter3));
  inv1  gate2455(.a(s_273), .O(gate53inter4));
  nand2 gate2456(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2457(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2458(.a(G13), .O(gate53inter7));
  inv1  gate2459(.a(G284), .O(gate53inter8));
  nand2 gate2460(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2461(.a(s_273), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2462(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2463(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2464(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1415(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1416(.a(gate56inter0), .b(s_124), .O(gate56inter1));
  and2  gate1417(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1418(.a(s_124), .O(gate56inter3));
  inv1  gate1419(.a(s_125), .O(gate56inter4));
  nand2 gate1420(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1421(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1422(.a(G16), .O(gate56inter7));
  inv1  gate1423(.a(G287), .O(gate56inter8));
  nand2 gate1424(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1425(.a(s_125), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1426(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1427(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1428(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate799(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate800(.a(gate57inter0), .b(s_36), .O(gate57inter1));
  and2  gate801(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate802(.a(s_36), .O(gate57inter3));
  inv1  gate803(.a(s_37), .O(gate57inter4));
  nand2 gate804(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate805(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate806(.a(G17), .O(gate57inter7));
  inv1  gate807(.a(G290), .O(gate57inter8));
  nand2 gate808(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate809(.a(s_37), .b(gate57inter3), .O(gate57inter10));
  nor2  gate810(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate811(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate812(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2689(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2690(.a(gate59inter0), .b(s_306), .O(gate59inter1));
  and2  gate2691(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2692(.a(s_306), .O(gate59inter3));
  inv1  gate2693(.a(s_307), .O(gate59inter4));
  nand2 gate2694(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2695(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2696(.a(G19), .O(gate59inter7));
  inv1  gate2697(.a(G293), .O(gate59inter8));
  nand2 gate2698(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2699(.a(s_307), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2700(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2701(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2702(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2297(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2298(.a(gate62inter0), .b(s_250), .O(gate62inter1));
  and2  gate2299(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2300(.a(s_250), .O(gate62inter3));
  inv1  gate2301(.a(s_251), .O(gate62inter4));
  nand2 gate2302(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2303(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2304(.a(G22), .O(gate62inter7));
  inv1  gate2305(.a(G296), .O(gate62inter8));
  nand2 gate2306(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2307(.a(s_251), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2308(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2309(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2310(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1205(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1206(.a(gate69inter0), .b(s_94), .O(gate69inter1));
  and2  gate1207(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1208(.a(s_94), .O(gate69inter3));
  inv1  gate1209(.a(s_95), .O(gate69inter4));
  nand2 gate1210(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1211(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1212(.a(G29), .O(gate69inter7));
  inv1  gate1213(.a(G308), .O(gate69inter8));
  nand2 gate1214(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1215(.a(s_95), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1216(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1217(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1218(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2577(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2578(.a(gate70inter0), .b(s_290), .O(gate70inter1));
  and2  gate2579(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2580(.a(s_290), .O(gate70inter3));
  inv1  gate2581(.a(s_291), .O(gate70inter4));
  nand2 gate2582(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2583(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2584(.a(G30), .O(gate70inter7));
  inv1  gate2585(.a(G308), .O(gate70inter8));
  nand2 gate2586(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2587(.a(s_291), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2588(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2589(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2590(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate2395(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2396(.a(gate71inter0), .b(s_264), .O(gate71inter1));
  and2  gate2397(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2398(.a(s_264), .O(gate71inter3));
  inv1  gate2399(.a(s_265), .O(gate71inter4));
  nand2 gate2400(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2401(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2402(.a(G31), .O(gate71inter7));
  inv1  gate2403(.a(G311), .O(gate71inter8));
  nand2 gate2404(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2405(.a(s_265), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2406(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2407(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2408(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1919(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1920(.a(gate75inter0), .b(s_196), .O(gate75inter1));
  and2  gate1921(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1922(.a(s_196), .O(gate75inter3));
  inv1  gate1923(.a(s_197), .O(gate75inter4));
  nand2 gate1924(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1925(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1926(.a(G9), .O(gate75inter7));
  inv1  gate1927(.a(G317), .O(gate75inter8));
  nand2 gate1928(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1929(.a(s_197), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1930(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1931(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1932(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2871(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2872(.a(gate77inter0), .b(s_332), .O(gate77inter1));
  and2  gate2873(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2874(.a(s_332), .O(gate77inter3));
  inv1  gate2875(.a(s_333), .O(gate77inter4));
  nand2 gate2876(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2877(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2878(.a(G2), .O(gate77inter7));
  inv1  gate2879(.a(G320), .O(gate77inter8));
  nand2 gate2880(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2881(.a(s_333), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2882(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2883(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2884(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate2353(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2354(.a(gate78inter0), .b(s_258), .O(gate78inter1));
  and2  gate2355(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2356(.a(s_258), .O(gate78inter3));
  inv1  gate2357(.a(s_259), .O(gate78inter4));
  nand2 gate2358(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2359(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2360(.a(G6), .O(gate78inter7));
  inv1  gate2361(.a(G320), .O(gate78inter8));
  nand2 gate2362(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2363(.a(s_259), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2364(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2365(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2366(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2927(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2928(.a(gate80inter0), .b(s_340), .O(gate80inter1));
  and2  gate2929(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2930(.a(s_340), .O(gate80inter3));
  inv1  gate2931(.a(s_341), .O(gate80inter4));
  nand2 gate2932(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2933(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2934(.a(G14), .O(gate80inter7));
  inv1  gate2935(.a(G323), .O(gate80inter8));
  nand2 gate2936(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2937(.a(s_341), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2938(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2939(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2940(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2423(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2424(.a(gate81inter0), .b(s_268), .O(gate81inter1));
  and2  gate2425(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2426(.a(s_268), .O(gate81inter3));
  inv1  gate2427(.a(s_269), .O(gate81inter4));
  nand2 gate2428(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2429(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2430(.a(G3), .O(gate81inter7));
  inv1  gate2431(.a(G326), .O(gate81inter8));
  nand2 gate2432(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2433(.a(s_269), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2434(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2435(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2436(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1793(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1794(.a(gate82inter0), .b(s_178), .O(gate82inter1));
  and2  gate1795(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1796(.a(s_178), .O(gate82inter3));
  inv1  gate1797(.a(s_179), .O(gate82inter4));
  nand2 gate1798(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1799(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1800(.a(G7), .O(gate82inter7));
  inv1  gate1801(.a(G326), .O(gate82inter8));
  nand2 gate1802(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1803(.a(s_179), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1804(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1805(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1806(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2367(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2368(.a(gate83inter0), .b(s_260), .O(gate83inter1));
  and2  gate2369(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2370(.a(s_260), .O(gate83inter3));
  inv1  gate2371(.a(s_261), .O(gate83inter4));
  nand2 gate2372(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2373(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2374(.a(G11), .O(gate83inter7));
  inv1  gate2375(.a(G329), .O(gate83inter8));
  nand2 gate2376(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2377(.a(s_261), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2378(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2379(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2380(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate2913(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2914(.a(gate84inter0), .b(s_338), .O(gate84inter1));
  and2  gate2915(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2916(.a(s_338), .O(gate84inter3));
  inv1  gate2917(.a(s_339), .O(gate84inter4));
  nand2 gate2918(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2919(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2920(.a(G15), .O(gate84inter7));
  inv1  gate2921(.a(G329), .O(gate84inter8));
  nand2 gate2922(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2923(.a(s_339), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2924(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2925(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2926(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate771(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate772(.a(gate85inter0), .b(s_32), .O(gate85inter1));
  and2  gate773(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate774(.a(s_32), .O(gate85inter3));
  inv1  gate775(.a(s_33), .O(gate85inter4));
  nand2 gate776(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate777(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate778(.a(G4), .O(gate85inter7));
  inv1  gate779(.a(G332), .O(gate85inter8));
  nand2 gate780(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate781(.a(s_33), .b(gate85inter3), .O(gate85inter10));
  nor2  gate782(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate783(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate784(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate729(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate730(.a(gate95inter0), .b(s_26), .O(gate95inter1));
  and2  gate731(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate732(.a(s_26), .O(gate95inter3));
  inv1  gate733(.a(s_27), .O(gate95inter4));
  nand2 gate734(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate735(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate736(.a(G26), .O(gate95inter7));
  inv1  gate737(.a(G347), .O(gate95inter8));
  nand2 gate738(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate739(.a(s_27), .b(gate95inter3), .O(gate95inter10));
  nor2  gate740(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate741(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate742(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate1471(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1472(.a(gate96inter0), .b(s_132), .O(gate96inter1));
  and2  gate1473(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1474(.a(s_132), .O(gate96inter3));
  inv1  gate1475(.a(s_133), .O(gate96inter4));
  nand2 gate1476(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1477(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1478(.a(G30), .O(gate96inter7));
  inv1  gate1479(.a(G347), .O(gate96inter8));
  nand2 gate1480(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1481(.a(s_133), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1482(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1483(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1484(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate883(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate884(.a(gate100inter0), .b(s_48), .O(gate100inter1));
  and2  gate885(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate886(.a(s_48), .O(gate100inter3));
  inv1  gate887(.a(s_49), .O(gate100inter4));
  nand2 gate888(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate889(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate890(.a(G31), .O(gate100inter7));
  inv1  gate891(.a(G353), .O(gate100inter8));
  nand2 gate892(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate893(.a(s_49), .b(gate100inter3), .O(gate100inter10));
  nor2  gate894(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate895(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate896(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1009(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1010(.a(gate101inter0), .b(s_66), .O(gate101inter1));
  and2  gate1011(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1012(.a(s_66), .O(gate101inter3));
  inv1  gate1013(.a(s_67), .O(gate101inter4));
  nand2 gate1014(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1015(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1016(.a(G20), .O(gate101inter7));
  inv1  gate1017(.a(G356), .O(gate101inter8));
  nand2 gate1018(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1019(.a(s_67), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1020(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1021(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1022(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2241(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2242(.a(gate102inter0), .b(s_242), .O(gate102inter1));
  and2  gate2243(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2244(.a(s_242), .O(gate102inter3));
  inv1  gate2245(.a(s_243), .O(gate102inter4));
  nand2 gate2246(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2247(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2248(.a(G24), .O(gate102inter7));
  inv1  gate2249(.a(G356), .O(gate102inter8));
  nand2 gate2250(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2251(.a(s_243), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2252(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2253(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2254(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate3081(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate3082(.a(gate108inter0), .b(s_362), .O(gate108inter1));
  and2  gate3083(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate3084(.a(s_362), .O(gate108inter3));
  inv1  gate3085(.a(s_363), .O(gate108inter4));
  nand2 gate3086(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate3087(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate3088(.a(G368), .O(gate108inter7));
  inv1  gate3089(.a(G369), .O(gate108inter8));
  nand2 gate3090(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate3091(.a(s_363), .b(gate108inter3), .O(gate108inter10));
  nor2  gate3092(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate3093(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate3094(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2829(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2830(.a(gate111inter0), .b(s_326), .O(gate111inter1));
  and2  gate2831(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2832(.a(s_326), .O(gate111inter3));
  inv1  gate2833(.a(s_327), .O(gate111inter4));
  nand2 gate2834(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2835(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2836(.a(G374), .O(gate111inter7));
  inv1  gate2837(.a(G375), .O(gate111inter8));
  nand2 gate2838(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2839(.a(s_327), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2840(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2841(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2842(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1387(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1388(.a(gate112inter0), .b(s_120), .O(gate112inter1));
  and2  gate1389(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1390(.a(s_120), .O(gate112inter3));
  inv1  gate1391(.a(s_121), .O(gate112inter4));
  nand2 gate1392(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1393(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1394(.a(G376), .O(gate112inter7));
  inv1  gate1395(.a(G377), .O(gate112inter8));
  nand2 gate1396(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1397(.a(s_121), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1398(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1399(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1400(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1877(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1878(.a(gate113inter0), .b(s_190), .O(gate113inter1));
  and2  gate1879(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1880(.a(s_190), .O(gate113inter3));
  inv1  gate1881(.a(s_191), .O(gate113inter4));
  nand2 gate1882(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1883(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1884(.a(G378), .O(gate113inter7));
  inv1  gate1885(.a(G379), .O(gate113inter8));
  nand2 gate1886(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1887(.a(s_191), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1888(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1889(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1890(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate939(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate940(.a(gate115inter0), .b(s_56), .O(gate115inter1));
  and2  gate941(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate942(.a(s_56), .O(gate115inter3));
  inv1  gate943(.a(s_57), .O(gate115inter4));
  nand2 gate944(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate945(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate946(.a(G382), .O(gate115inter7));
  inv1  gate947(.a(G383), .O(gate115inter8));
  nand2 gate948(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate949(.a(s_57), .b(gate115inter3), .O(gate115inter10));
  nor2  gate950(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate951(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate952(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1373(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1374(.a(gate119inter0), .b(s_118), .O(gate119inter1));
  and2  gate1375(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1376(.a(s_118), .O(gate119inter3));
  inv1  gate1377(.a(s_119), .O(gate119inter4));
  nand2 gate1378(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1379(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1380(.a(G390), .O(gate119inter7));
  inv1  gate1381(.a(G391), .O(gate119inter8));
  nand2 gate1382(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1383(.a(s_119), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1384(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1385(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1386(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1555(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1556(.a(gate120inter0), .b(s_144), .O(gate120inter1));
  and2  gate1557(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1558(.a(s_144), .O(gate120inter3));
  inv1  gate1559(.a(s_145), .O(gate120inter4));
  nand2 gate1560(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1561(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1562(.a(G392), .O(gate120inter7));
  inv1  gate1563(.a(G393), .O(gate120inter8));
  nand2 gate1564(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1565(.a(s_145), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1566(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1567(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1568(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate1961(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1962(.a(gate121inter0), .b(s_202), .O(gate121inter1));
  and2  gate1963(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1964(.a(s_202), .O(gate121inter3));
  inv1  gate1965(.a(s_203), .O(gate121inter4));
  nand2 gate1966(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1967(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1968(.a(G394), .O(gate121inter7));
  inv1  gate1969(.a(G395), .O(gate121inter8));
  nand2 gate1970(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1971(.a(s_203), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1972(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1973(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1974(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1779(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1780(.a(gate122inter0), .b(s_176), .O(gate122inter1));
  and2  gate1781(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1782(.a(s_176), .O(gate122inter3));
  inv1  gate1783(.a(s_177), .O(gate122inter4));
  nand2 gate1784(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1785(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1786(.a(G396), .O(gate122inter7));
  inv1  gate1787(.a(G397), .O(gate122inter8));
  nand2 gate1788(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1789(.a(s_177), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1790(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1791(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1792(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate2101(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2102(.a(gate123inter0), .b(s_222), .O(gate123inter1));
  and2  gate2103(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2104(.a(s_222), .O(gate123inter3));
  inv1  gate2105(.a(s_223), .O(gate123inter4));
  nand2 gate2106(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2107(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2108(.a(G398), .O(gate123inter7));
  inv1  gate2109(.a(G399), .O(gate123inter8));
  nand2 gate2110(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2111(.a(s_223), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2112(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2113(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2114(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2521(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2522(.a(gate125inter0), .b(s_282), .O(gate125inter1));
  and2  gate2523(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2524(.a(s_282), .O(gate125inter3));
  inv1  gate2525(.a(s_283), .O(gate125inter4));
  nand2 gate2526(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2527(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2528(.a(G402), .O(gate125inter7));
  inv1  gate2529(.a(G403), .O(gate125inter8));
  nand2 gate2530(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2531(.a(s_283), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2532(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2533(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2534(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate3053(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate3054(.a(gate128inter0), .b(s_358), .O(gate128inter1));
  and2  gate3055(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate3056(.a(s_358), .O(gate128inter3));
  inv1  gate3057(.a(s_359), .O(gate128inter4));
  nand2 gate3058(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate3059(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate3060(.a(G408), .O(gate128inter7));
  inv1  gate3061(.a(G409), .O(gate128inter8));
  nand2 gate3062(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate3063(.a(s_359), .b(gate128inter3), .O(gate128inter10));
  nor2  gate3064(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate3065(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate3066(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate2213(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2214(.a(gate133inter0), .b(s_238), .O(gate133inter1));
  and2  gate2215(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2216(.a(s_238), .O(gate133inter3));
  inv1  gate2217(.a(s_239), .O(gate133inter4));
  nand2 gate2218(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2219(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2220(.a(G418), .O(gate133inter7));
  inv1  gate2221(.a(G419), .O(gate133inter8));
  nand2 gate2222(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2223(.a(s_239), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2224(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2225(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2226(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2703(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2704(.a(gate138inter0), .b(s_308), .O(gate138inter1));
  and2  gate2705(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2706(.a(s_308), .O(gate138inter3));
  inv1  gate2707(.a(s_309), .O(gate138inter4));
  nand2 gate2708(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2709(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2710(.a(G432), .O(gate138inter7));
  inv1  gate2711(.a(G435), .O(gate138inter8));
  nand2 gate2712(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2713(.a(s_309), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2714(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2715(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2716(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2171(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2172(.a(gate143inter0), .b(s_232), .O(gate143inter1));
  and2  gate2173(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2174(.a(s_232), .O(gate143inter3));
  inv1  gate2175(.a(s_233), .O(gate143inter4));
  nand2 gate2176(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2177(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2178(.a(G462), .O(gate143inter7));
  inv1  gate2179(.a(G465), .O(gate143inter8));
  nand2 gate2180(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2181(.a(s_233), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2182(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2183(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2184(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate2339(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2340(.a(gate144inter0), .b(s_256), .O(gate144inter1));
  and2  gate2341(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2342(.a(s_256), .O(gate144inter3));
  inv1  gate2343(.a(s_257), .O(gate144inter4));
  nand2 gate2344(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2345(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2346(.a(G468), .O(gate144inter7));
  inv1  gate2347(.a(G471), .O(gate144inter8));
  nand2 gate2348(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2349(.a(s_257), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2350(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2351(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2352(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2255(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2256(.a(gate149inter0), .b(s_244), .O(gate149inter1));
  and2  gate2257(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2258(.a(s_244), .O(gate149inter3));
  inv1  gate2259(.a(s_245), .O(gate149inter4));
  nand2 gate2260(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2261(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2262(.a(G498), .O(gate149inter7));
  inv1  gate2263(.a(G501), .O(gate149inter8));
  nand2 gate2264(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2265(.a(s_245), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2266(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2267(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2268(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1989(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1990(.a(gate151inter0), .b(s_206), .O(gate151inter1));
  and2  gate1991(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1992(.a(s_206), .O(gate151inter3));
  inv1  gate1993(.a(s_207), .O(gate151inter4));
  nand2 gate1994(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1995(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1996(.a(G510), .O(gate151inter7));
  inv1  gate1997(.a(G513), .O(gate151inter8));
  nand2 gate1998(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1999(.a(s_207), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2000(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2001(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2002(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1261(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1262(.a(gate154inter0), .b(s_102), .O(gate154inter1));
  and2  gate1263(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1264(.a(s_102), .O(gate154inter3));
  inv1  gate1265(.a(s_103), .O(gate154inter4));
  nand2 gate1266(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1267(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1268(.a(G429), .O(gate154inter7));
  inv1  gate1269(.a(G522), .O(gate154inter8));
  nand2 gate1270(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1271(.a(s_103), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1272(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1273(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1274(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1541(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1542(.a(gate161inter0), .b(s_142), .O(gate161inter1));
  and2  gate1543(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1544(.a(s_142), .O(gate161inter3));
  inv1  gate1545(.a(s_143), .O(gate161inter4));
  nand2 gate1546(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1547(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1548(.a(G450), .O(gate161inter7));
  inv1  gate1549(.a(G534), .O(gate161inter8));
  nand2 gate1550(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1551(.a(s_143), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1552(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1553(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1554(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1611(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1612(.a(gate162inter0), .b(s_152), .O(gate162inter1));
  and2  gate1613(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1614(.a(s_152), .O(gate162inter3));
  inv1  gate1615(.a(s_153), .O(gate162inter4));
  nand2 gate1616(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1617(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1618(.a(G453), .O(gate162inter7));
  inv1  gate1619(.a(G534), .O(gate162inter8));
  nand2 gate1620(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1621(.a(s_153), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1622(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1623(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1624(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1345(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1346(.a(gate164inter0), .b(s_114), .O(gate164inter1));
  and2  gate1347(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1348(.a(s_114), .O(gate164inter3));
  inv1  gate1349(.a(s_115), .O(gate164inter4));
  nand2 gate1350(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1351(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1352(.a(G459), .O(gate164inter7));
  inv1  gate1353(.a(G537), .O(gate164inter8));
  nand2 gate1354(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1355(.a(s_115), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1356(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1357(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1358(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate2031(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2032(.a(gate165inter0), .b(s_212), .O(gate165inter1));
  and2  gate2033(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2034(.a(s_212), .O(gate165inter3));
  inv1  gate2035(.a(s_213), .O(gate165inter4));
  nand2 gate2036(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2037(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2038(.a(G462), .O(gate165inter7));
  inv1  gate2039(.a(G540), .O(gate165inter8));
  nand2 gate2040(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2041(.a(s_213), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2042(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2043(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2044(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate2745(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2746(.a(gate166inter0), .b(s_314), .O(gate166inter1));
  and2  gate2747(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2748(.a(s_314), .O(gate166inter3));
  inv1  gate2749(.a(s_315), .O(gate166inter4));
  nand2 gate2750(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2751(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2752(.a(G465), .O(gate166inter7));
  inv1  gate2753(.a(G540), .O(gate166inter8));
  nand2 gate2754(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2755(.a(s_315), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2756(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2757(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2758(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2675(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2676(.a(gate167inter0), .b(s_304), .O(gate167inter1));
  and2  gate2677(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2678(.a(s_304), .O(gate167inter3));
  inv1  gate2679(.a(s_305), .O(gate167inter4));
  nand2 gate2680(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2681(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2682(.a(G468), .O(gate167inter7));
  inv1  gate2683(.a(G543), .O(gate167inter8));
  nand2 gate2684(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2685(.a(s_305), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2686(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2687(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2688(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1905(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1906(.a(gate168inter0), .b(s_194), .O(gate168inter1));
  and2  gate1907(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1908(.a(s_194), .O(gate168inter3));
  inv1  gate1909(.a(s_195), .O(gate168inter4));
  nand2 gate1910(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1911(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1912(.a(G471), .O(gate168inter7));
  inv1  gate1913(.a(G543), .O(gate168inter8));
  nand2 gate1914(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1915(.a(s_195), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1916(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1917(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1918(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate869(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate870(.a(gate169inter0), .b(s_46), .O(gate169inter1));
  and2  gate871(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate872(.a(s_46), .O(gate169inter3));
  inv1  gate873(.a(s_47), .O(gate169inter4));
  nand2 gate874(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate875(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate876(.a(G474), .O(gate169inter7));
  inv1  gate877(.a(G546), .O(gate169inter8));
  nand2 gate878(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate879(.a(s_47), .b(gate169inter3), .O(gate169inter10));
  nor2  gate880(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate881(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate882(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate995(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate996(.a(gate176inter0), .b(s_64), .O(gate176inter1));
  and2  gate997(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate998(.a(s_64), .O(gate176inter3));
  inv1  gate999(.a(s_65), .O(gate176inter4));
  nand2 gate1000(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1001(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1002(.a(G495), .O(gate176inter7));
  inv1  gate1003(.a(G555), .O(gate176inter8));
  nand2 gate1004(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1005(.a(s_65), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1006(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1007(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1008(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate617(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate618(.a(gate178inter0), .b(s_10), .O(gate178inter1));
  and2  gate619(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate620(.a(s_10), .O(gate178inter3));
  inv1  gate621(.a(s_11), .O(gate178inter4));
  nand2 gate622(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate623(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate624(.a(G501), .O(gate178inter7));
  inv1  gate625(.a(G558), .O(gate178inter8));
  nand2 gate626(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate627(.a(s_11), .b(gate178inter3), .O(gate178inter10));
  nor2  gate628(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate629(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate630(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate3095(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate3096(.a(gate183inter0), .b(s_364), .O(gate183inter1));
  and2  gate3097(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate3098(.a(s_364), .O(gate183inter3));
  inv1  gate3099(.a(s_365), .O(gate183inter4));
  nand2 gate3100(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate3101(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate3102(.a(G516), .O(gate183inter7));
  inv1  gate3103(.a(G567), .O(gate183inter8));
  nand2 gate3104(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate3105(.a(s_365), .b(gate183inter3), .O(gate183inter10));
  nor2  gate3106(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate3107(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate3108(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1737(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1738(.a(gate184inter0), .b(s_170), .O(gate184inter1));
  and2  gate1739(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1740(.a(s_170), .O(gate184inter3));
  inv1  gate1741(.a(s_171), .O(gate184inter4));
  nand2 gate1742(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1743(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1744(.a(G519), .O(gate184inter7));
  inv1  gate1745(.a(G567), .O(gate184inter8));
  nand2 gate1746(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1747(.a(s_171), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1748(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1749(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1750(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2157(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2158(.a(gate185inter0), .b(s_230), .O(gate185inter1));
  and2  gate2159(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2160(.a(s_230), .O(gate185inter3));
  inv1  gate2161(.a(s_231), .O(gate185inter4));
  nand2 gate2162(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2163(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2164(.a(G570), .O(gate185inter7));
  inv1  gate2165(.a(G571), .O(gate185inter8));
  nand2 gate2166(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2167(.a(s_231), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2168(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2169(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2170(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2003(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2004(.a(gate186inter0), .b(s_208), .O(gate186inter1));
  and2  gate2005(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2006(.a(s_208), .O(gate186inter3));
  inv1  gate2007(.a(s_209), .O(gate186inter4));
  nand2 gate2008(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2009(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2010(.a(G572), .O(gate186inter7));
  inv1  gate2011(.a(G573), .O(gate186inter8));
  nand2 gate2012(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2013(.a(s_209), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2014(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2015(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2016(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate2381(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2382(.a(gate187inter0), .b(s_262), .O(gate187inter1));
  and2  gate2383(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2384(.a(s_262), .O(gate187inter3));
  inv1  gate2385(.a(s_263), .O(gate187inter4));
  nand2 gate2386(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2387(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2388(.a(G574), .O(gate187inter7));
  inv1  gate2389(.a(G575), .O(gate187inter8));
  nand2 gate2390(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2391(.a(s_263), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2392(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2393(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2394(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate589(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate590(.a(gate190inter0), .b(s_6), .O(gate190inter1));
  and2  gate591(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate592(.a(s_6), .O(gate190inter3));
  inv1  gate593(.a(s_7), .O(gate190inter4));
  nand2 gate594(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate595(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate596(.a(G580), .O(gate190inter7));
  inv1  gate597(.a(G581), .O(gate190inter8));
  nand2 gate598(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate599(.a(s_7), .b(gate190inter3), .O(gate190inter10));
  nor2  gate600(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate601(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate602(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1527(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1528(.a(gate192inter0), .b(s_140), .O(gate192inter1));
  and2  gate1529(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1530(.a(s_140), .O(gate192inter3));
  inv1  gate1531(.a(s_141), .O(gate192inter4));
  nand2 gate1532(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1533(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1534(.a(G584), .O(gate192inter7));
  inv1  gate1535(.a(G585), .O(gate192inter8));
  nand2 gate1536(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1537(.a(s_141), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1538(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1539(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1540(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate701(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate702(.a(gate196inter0), .b(s_22), .O(gate196inter1));
  and2  gate703(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate704(.a(s_22), .O(gate196inter3));
  inv1  gate705(.a(s_23), .O(gate196inter4));
  nand2 gate706(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate707(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate708(.a(G592), .O(gate196inter7));
  inv1  gate709(.a(G593), .O(gate196inter8));
  nand2 gate710(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate711(.a(s_23), .b(gate196inter3), .O(gate196inter10));
  nor2  gate712(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate713(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate714(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2899(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2900(.a(gate198inter0), .b(s_336), .O(gate198inter1));
  and2  gate2901(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2902(.a(s_336), .O(gate198inter3));
  inv1  gate2903(.a(s_337), .O(gate198inter4));
  nand2 gate2904(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2905(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2906(.a(G596), .O(gate198inter7));
  inv1  gate2907(.a(G597), .O(gate198inter8));
  nand2 gate2908(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2909(.a(s_337), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2910(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2911(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2912(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2815(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2816(.a(gate199inter0), .b(s_324), .O(gate199inter1));
  and2  gate2817(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2818(.a(s_324), .O(gate199inter3));
  inv1  gate2819(.a(s_325), .O(gate199inter4));
  nand2 gate2820(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2821(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2822(.a(G598), .O(gate199inter7));
  inv1  gate2823(.a(G599), .O(gate199inter8));
  nand2 gate2824(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2825(.a(s_325), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2826(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2827(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2828(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate687(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate688(.a(gate200inter0), .b(s_20), .O(gate200inter1));
  and2  gate689(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate690(.a(s_20), .O(gate200inter3));
  inv1  gate691(.a(s_21), .O(gate200inter4));
  nand2 gate692(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate693(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate694(.a(G600), .O(gate200inter7));
  inv1  gate695(.a(G601), .O(gate200inter8));
  nand2 gate696(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate697(.a(s_21), .b(gate200inter3), .O(gate200inter10));
  nor2  gate698(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate699(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate700(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate3137(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate3138(.a(gate201inter0), .b(s_370), .O(gate201inter1));
  and2  gate3139(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate3140(.a(s_370), .O(gate201inter3));
  inv1  gate3141(.a(s_371), .O(gate201inter4));
  nand2 gate3142(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate3143(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate3144(.a(G602), .O(gate201inter7));
  inv1  gate3145(.a(G607), .O(gate201inter8));
  nand2 gate3146(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate3147(.a(s_371), .b(gate201inter3), .O(gate201inter10));
  nor2  gate3148(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate3149(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate3150(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2997(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2998(.a(gate205inter0), .b(s_350), .O(gate205inter1));
  and2  gate2999(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate3000(.a(s_350), .O(gate205inter3));
  inv1  gate3001(.a(s_351), .O(gate205inter4));
  nand2 gate3002(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate3003(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate3004(.a(G622), .O(gate205inter7));
  inv1  gate3005(.a(G627), .O(gate205inter8));
  nand2 gate3006(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate3007(.a(s_351), .b(gate205inter3), .O(gate205inter10));
  nor2  gate3008(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate3009(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate3010(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1751(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1752(.a(gate208inter0), .b(s_172), .O(gate208inter1));
  and2  gate1753(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1754(.a(s_172), .O(gate208inter3));
  inv1  gate1755(.a(s_173), .O(gate208inter4));
  nand2 gate1756(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1757(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1758(.a(G627), .O(gate208inter7));
  inv1  gate1759(.a(G637), .O(gate208inter8));
  nand2 gate1760(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1761(.a(s_173), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1762(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1763(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1764(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2115(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2116(.a(gate214inter0), .b(s_224), .O(gate214inter1));
  and2  gate2117(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2118(.a(s_224), .O(gate214inter3));
  inv1  gate2119(.a(s_225), .O(gate214inter4));
  nand2 gate2120(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2121(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2122(.a(G612), .O(gate214inter7));
  inv1  gate2123(.a(G672), .O(gate214inter8));
  nand2 gate2124(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2125(.a(s_225), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2126(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2127(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2128(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate561(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate562(.a(gate215inter0), .b(s_2), .O(gate215inter1));
  and2  gate563(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate564(.a(s_2), .O(gate215inter3));
  inv1  gate565(.a(s_3), .O(gate215inter4));
  nand2 gate566(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate567(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate568(.a(G607), .O(gate215inter7));
  inv1  gate569(.a(G675), .O(gate215inter8));
  nand2 gate570(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate571(.a(s_3), .b(gate215inter3), .O(gate215inter10));
  nor2  gate572(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate573(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate574(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1485(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1486(.a(gate216inter0), .b(s_134), .O(gate216inter1));
  and2  gate1487(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1488(.a(s_134), .O(gate216inter3));
  inv1  gate1489(.a(s_135), .O(gate216inter4));
  nand2 gate1490(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1491(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1492(.a(G617), .O(gate216inter7));
  inv1  gate1493(.a(G675), .O(gate216inter8));
  nand2 gate1494(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1495(.a(s_135), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1496(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1497(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1498(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1093(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1094(.a(gate223inter0), .b(s_78), .O(gate223inter1));
  and2  gate1095(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1096(.a(s_78), .O(gate223inter3));
  inv1  gate1097(.a(s_79), .O(gate223inter4));
  nand2 gate1098(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1099(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1100(.a(G627), .O(gate223inter7));
  inv1  gate1101(.a(G687), .O(gate223inter8));
  nand2 gate1102(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1103(.a(s_79), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1104(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1105(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1106(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate841(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate842(.a(gate231inter0), .b(s_42), .O(gate231inter1));
  and2  gate843(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate844(.a(s_42), .O(gate231inter3));
  inv1  gate845(.a(s_43), .O(gate231inter4));
  nand2 gate846(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate847(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate848(.a(G702), .O(gate231inter7));
  inv1  gate849(.a(G703), .O(gate231inter8));
  nand2 gate850(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate851(.a(s_43), .b(gate231inter3), .O(gate231inter10));
  nor2  gate852(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate853(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate854(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2479(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2480(.a(gate232inter0), .b(s_276), .O(gate232inter1));
  and2  gate2481(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2482(.a(s_276), .O(gate232inter3));
  inv1  gate2483(.a(s_277), .O(gate232inter4));
  nand2 gate2484(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2485(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2486(.a(G704), .O(gate232inter7));
  inv1  gate2487(.a(G705), .O(gate232inter8));
  nand2 gate2488(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2489(.a(s_277), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2490(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2491(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2492(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate813(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate814(.a(gate234inter0), .b(s_38), .O(gate234inter1));
  and2  gate815(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate816(.a(s_38), .O(gate234inter3));
  inv1  gate817(.a(s_39), .O(gate234inter4));
  nand2 gate818(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate819(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate820(.a(G245), .O(gate234inter7));
  inv1  gate821(.a(G721), .O(gate234inter8));
  nand2 gate822(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate823(.a(s_39), .b(gate234inter3), .O(gate234inter10));
  nor2  gate824(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate825(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate826(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1429(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1430(.a(gate236inter0), .b(s_126), .O(gate236inter1));
  and2  gate1431(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1432(.a(s_126), .O(gate236inter3));
  inv1  gate1433(.a(s_127), .O(gate236inter4));
  nand2 gate1434(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1435(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1436(.a(G251), .O(gate236inter7));
  inv1  gate1437(.a(G727), .O(gate236inter8));
  nand2 gate1438(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1439(.a(s_127), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1440(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1441(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1442(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1219(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1220(.a(gate237inter0), .b(s_96), .O(gate237inter1));
  and2  gate1221(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1222(.a(s_96), .O(gate237inter3));
  inv1  gate1223(.a(s_97), .O(gate237inter4));
  nand2 gate1224(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1225(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1226(.a(G254), .O(gate237inter7));
  inv1  gate1227(.a(G706), .O(gate237inter8));
  nand2 gate1228(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1229(.a(s_97), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1230(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1231(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1232(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1513(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1514(.a(gate238inter0), .b(s_138), .O(gate238inter1));
  and2  gate1515(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1516(.a(s_138), .O(gate238inter3));
  inv1  gate1517(.a(s_139), .O(gate238inter4));
  nand2 gate1518(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1519(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1520(.a(G257), .O(gate238inter7));
  inv1  gate1521(.a(G709), .O(gate238inter8));
  nand2 gate1522(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1523(.a(s_139), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1524(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1525(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1526(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate785(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate786(.a(gate240inter0), .b(s_34), .O(gate240inter1));
  and2  gate787(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate788(.a(s_34), .O(gate240inter3));
  inv1  gate789(.a(s_35), .O(gate240inter4));
  nand2 gate790(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate791(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate792(.a(G263), .O(gate240inter7));
  inv1  gate793(.a(G715), .O(gate240inter8));
  nand2 gate794(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate795(.a(s_35), .b(gate240inter3), .O(gate240inter10));
  nor2  gate796(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate797(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate798(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1723(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1724(.a(gate241inter0), .b(s_168), .O(gate241inter1));
  and2  gate1725(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1726(.a(s_168), .O(gate241inter3));
  inv1  gate1727(.a(s_169), .O(gate241inter4));
  nand2 gate1728(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1729(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1730(.a(G242), .O(gate241inter7));
  inv1  gate1731(.a(G730), .O(gate241inter8));
  nand2 gate1732(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1733(.a(s_169), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1734(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1735(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1736(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate911(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate912(.a(gate243inter0), .b(s_52), .O(gate243inter1));
  and2  gate913(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate914(.a(s_52), .O(gate243inter3));
  inv1  gate915(.a(s_53), .O(gate243inter4));
  nand2 gate916(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate917(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate918(.a(G245), .O(gate243inter7));
  inv1  gate919(.a(G733), .O(gate243inter8));
  nand2 gate920(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate921(.a(s_53), .b(gate243inter3), .O(gate243inter10));
  nor2  gate922(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate923(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate924(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1065(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1066(.a(gate244inter0), .b(s_74), .O(gate244inter1));
  and2  gate1067(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1068(.a(s_74), .O(gate244inter3));
  inv1  gate1069(.a(s_75), .O(gate244inter4));
  nand2 gate1070(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1071(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1072(.a(G721), .O(gate244inter7));
  inv1  gate1073(.a(G733), .O(gate244inter8));
  nand2 gate1074(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1075(.a(s_75), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1076(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1077(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1078(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1317(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1318(.a(gate248inter0), .b(s_110), .O(gate248inter1));
  and2  gate1319(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1320(.a(s_110), .O(gate248inter3));
  inv1  gate1321(.a(s_111), .O(gate248inter4));
  nand2 gate1322(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1323(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1324(.a(G727), .O(gate248inter7));
  inv1  gate1325(.a(G739), .O(gate248inter8));
  nand2 gate1326(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1327(.a(s_111), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1328(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1329(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1330(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2087(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2088(.a(gate252inter0), .b(s_220), .O(gate252inter1));
  and2  gate2089(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2090(.a(s_220), .O(gate252inter3));
  inv1  gate2091(.a(s_221), .O(gate252inter4));
  nand2 gate2092(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2093(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2094(.a(G709), .O(gate252inter7));
  inv1  gate2095(.a(G745), .O(gate252inter8));
  nand2 gate2096(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2097(.a(s_221), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2098(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2099(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2100(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate3025(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate3026(.a(gate256inter0), .b(s_354), .O(gate256inter1));
  and2  gate3027(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate3028(.a(s_354), .O(gate256inter3));
  inv1  gate3029(.a(s_355), .O(gate256inter4));
  nand2 gate3030(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate3031(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate3032(.a(G715), .O(gate256inter7));
  inv1  gate3033(.a(G751), .O(gate256inter8));
  nand2 gate3034(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate3035(.a(s_355), .b(gate256inter3), .O(gate256inter10));
  nor2  gate3036(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate3037(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate3038(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1247(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1248(.a(gate257inter0), .b(s_100), .O(gate257inter1));
  and2  gate1249(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1250(.a(s_100), .O(gate257inter3));
  inv1  gate1251(.a(s_101), .O(gate257inter4));
  nand2 gate1252(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1253(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1254(.a(G754), .O(gate257inter7));
  inv1  gate1255(.a(G755), .O(gate257inter8));
  nand2 gate1256(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1257(.a(s_101), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1258(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1259(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1260(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1023(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1024(.a(gate260inter0), .b(s_68), .O(gate260inter1));
  and2  gate1025(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1026(.a(s_68), .O(gate260inter3));
  inv1  gate1027(.a(s_69), .O(gate260inter4));
  nand2 gate1028(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1029(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1030(.a(G760), .O(gate260inter7));
  inv1  gate1031(.a(G761), .O(gate260inter8));
  nand2 gate1032(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1033(.a(s_69), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1034(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1035(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1036(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate3011(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate3012(.a(gate261inter0), .b(s_352), .O(gate261inter1));
  and2  gate3013(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate3014(.a(s_352), .O(gate261inter3));
  inv1  gate3015(.a(s_353), .O(gate261inter4));
  nand2 gate3016(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate3017(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate3018(.a(G762), .O(gate261inter7));
  inv1  gate3019(.a(G763), .O(gate261inter8));
  nand2 gate3020(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate3021(.a(s_353), .b(gate261inter3), .O(gate261inter10));
  nor2  gate3022(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate3023(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate3024(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate2227(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2228(.a(gate262inter0), .b(s_240), .O(gate262inter1));
  and2  gate2229(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2230(.a(s_240), .O(gate262inter3));
  inv1  gate2231(.a(s_241), .O(gate262inter4));
  nand2 gate2232(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2233(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2234(.a(G764), .O(gate262inter7));
  inv1  gate2235(.a(G765), .O(gate262inter8));
  nand2 gate2236(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2237(.a(s_241), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2238(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2239(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2240(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2605(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2606(.a(gate263inter0), .b(s_294), .O(gate263inter1));
  and2  gate2607(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2608(.a(s_294), .O(gate263inter3));
  inv1  gate2609(.a(s_295), .O(gate263inter4));
  nand2 gate2610(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2611(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2612(.a(G766), .O(gate263inter7));
  inv1  gate2613(.a(G767), .O(gate263inter8));
  nand2 gate2614(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2615(.a(s_295), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2616(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2617(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2618(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1401(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1402(.a(gate264inter0), .b(s_122), .O(gate264inter1));
  and2  gate1403(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1404(.a(s_122), .O(gate264inter3));
  inv1  gate1405(.a(s_123), .O(gate264inter4));
  nand2 gate1406(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1407(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1408(.a(G768), .O(gate264inter7));
  inv1  gate1409(.a(G769), .O(gate264inter8));
  nand2 gate1410(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1411(.a(s_123), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1412(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1413(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1414(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate2199(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2200(.a(gate265inter0), .b(s_236), .O(gate265inter1));
  and2  gate2201(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2202(.a(s_236), .O(gate265inter3));
  inv1  gate2203(.a(s_237), .O(gate265inter4));
  nand2 gate2204(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2205(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2206(.a(G642), .O(gate265inter7));
  inv1  gate2207(.a(G770), .O(gate265inter8));
  nand2 gate2208(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2209(.a(s_237), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2210(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2211(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2212(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2787(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2788(.a(gate268inter0), .b(s_320), .O(gate268inter1));
  and2  gate2789(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2790(.a(s_320), .O(gate268inter3));
  inv1  gate2791(.a(s_321), .O(gate268inter4));
  nand2 gate2792(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2793(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2794(.a(G651), .O(gate268inter7));
  inv1  gate2795(.a(G779), .O(gate268inter8));
  nand2 gate2796(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2797(.a(s_321), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2798(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2799(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2800(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1653(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1654(.a(gate269inter0), .b(s_158), .O(gate269inter1));
  and2  gate1655(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1656(.a(s_158), .O(gate269inter3));
  inv1  gate1657(.a(s_159), .O(gate269inter4));
  nand2 gate1658(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1659(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1660(.a(G654), .O(gate269inter7));
  inv1  gate1661(.a(G782), .O(gate269inter8));
  nand2 gate1662(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1663(.a(s_159), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1664(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1665(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1666(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate743(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate744(.a(gate270inter0), .b(s_28), .O(gate270inter1));
  and2  gate745(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate746(.a(s_28), .O(gate270inter3));
  inv1  gate747(.a(s_29), .O(gate270inter4));
  nand2 gate748(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate749(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate750(.a(G657), .O(gate270inter7));
  inv1  gate751(.a(G785), .O(gate270inter8));
  nand2 gate752(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate753(.a(s_29), .b(gate270inter3), .O(gate270inter10));
  nor2  gate754(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate755(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate756(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate603(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate604(.a(gate274inter0), .b(s_8), .O(gate274inter1));
  and2  gate605(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate606(.a(s_8), .O(gate274inter3));
  inv1  gate607(.a(s_9), .O(gate274inter4));
  nand2 gate608(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate609(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate610(.a(G770), .O(gate274inter7));
  inv1  gate611(.a(G794), .O(gate274inter8));
  nand2 gate612(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate613(.a(s_9), .b(gate274inter3), .O(gate274inter10));
  nor2  gate614(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate615(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate616(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2955(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2956(.a(gate275inter0), .b(s_344), .O(gate275inter1));
  and2  gate2957(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2958(.a(s_344), .O(gate275inter3));
  inv1  gate2959(.a(s_345), .O(gate275inter4));
  nand2 gate2960(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2961(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2962(.a(G645), .O(gate275inter7));
  inv1  gate2963(.a(G797), .O(gate275inter8));
  nand2 gate2964(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2965(.a(s_345), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2966(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2967(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2968(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1149(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1150(.a(gate282inter0), .b(s_86), .O(gate282inter1));
  and2  gate1151(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1152(.a(s_86), .O(gate282inter3));
  inv1  gate1153(.a(s_87), .O(gate282inter4));
  nand2 gate1154(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1155(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1156(.a(G782), .O(gate282inter7));
  inv1  gate1157(.a(G806), .O(gate282inter8));
  nand2 gate1158(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1159(.a(s_87), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1160(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1161(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1162(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2325(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2326(.a(gate288inter0), .b(s_254), .O(gate288inter1));
  and2  gate2327(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2328(.a(s_254), .O(gate288inter3));
  inv1  gate2329(.a(s_255), .O(gate288inter4));
  nand2 gate2330(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2331(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2332(.a(G791), .O(gate288inter7));
  inv1  gate2333(.a(G815), .O(gate288inter8));
  nand2 gate2334(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2335(.a(s_255), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2336(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2337(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2338(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1135(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1136(.a(gate289inter0), .b(s_84), .O(gate289inter1));
  and2  gate1137(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1138(.a(s_84), .O(gate289inter3));
  inv1  gate1139(.a(s_85), .O(gate289inter4));
  nand2 gate1140(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1141(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1142(.a(G818), .O(gate289inter7));
  inv1  gate1143(.a(G819), .O(gate289inter8));
  nand2 gate1144(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1145(.a(s_85), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1146(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1147(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1148(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate757(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate758(.a(gate290inter0), .b(s_30), .O(gate290inter1));
  and2  gate759(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate760(.a(s_30), .O(gate290inter3));
  inv1  gate761(.a(s_31), .O(gate290inter4));
  nand2 gate762(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate763(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate764(.a(G820), .O(gate290inter7));
  inv1  gate765(.a(G821), .O(gate290inter8));
  nand2 gate766(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate767(.a(s_31), .b(gate290inter3), .O(gate290inter10));
  nor2  gate768(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate769(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate770(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2983(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2984(.a(gate294inter0), .b(s_348), .O(gate294inter1));
  and2  gate2985(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2986(.a(s_348), .O(gate294inter3));
  inv1  gate2987(.a(s_349), .O(gate294inter4));
  nand2 gate2988(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2989(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2990(.a(G832), .O(gate294inter7));
  inv1  gate2991(.a(G833), .O(gate294inter8));
  nand2 gate2992(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2993(.a(s_349), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2994(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2995(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2996(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2073(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2074(.a(gate295inter0), .b(s_218), .O(gate295inter1));
  and2  gate2075(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2076(.a(s_218), .O(gate295inter3));
  inv1  gate2077(.a(s_219), .O(gate295inter4));
  nand2 gate2078(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2079(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2080(.a(G830), .O(gate295inter7));
  inv1  gate2081(.a(G831), .O(gate295inter8));
  nand2 gate2082(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2083(.a(s_219), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2084(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2085(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2086(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1709(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1710(.a(gate296inter0), .b(s_166), .O(gate296inter1));
  and2  gate1711(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1712(.a(s_166), .O(gate296inter3));
  inv1  gate1713(.a(s_167), .O(gate296inter4));
  nand2 gate1714(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1715(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1716(.a(G826), .O(gate296inter7));
  inv1  gate1717(.a(G827), .O(gate296inter8));
  nand2 gate1718(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1719(.a(s_167), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1720(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1721(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1722(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate659(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate660(.a(gate387inter0), .b(s_16), .O(gate387inter1));
  and2  gate661(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate662(.a(s_16), .O(gate387inter3));
  inv1  gate663(.a(s_17), .O(gate387inter4));
  nand2 gate664(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate665(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate666(.a(G1), .O(gate387inter7));
  inv1  gate667(.a(G1036), .O(gate387inter8));
  nand2 gate668(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate669(.a(s_17), .b(gate387inter3), .O(gate387inter10));
  nor2  gate670(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate671(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate672(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2633(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2634(.a(gate391inter0), .b(s_298), .O(gate391inter1));
  and2  gate2635(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2636(.a(s_298), .O(gate391inter3));
  inv1  gate2637(.a(s_299), .O(gate391inter4));
  nand2 gate2638(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2639(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2640(.a(G5), .O(gate391inter7));
  inv1  gate2641(.a(G1048), .O(gate391inter8));
  nand2 gate2642(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2643(.a(s_299), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2644(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2645(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2646(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate2857(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2858(.a(gate392inter0), .b(s_330), .O(gate392inter1));
  and2  gate2859(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2860(.a(s_330), .O(gate392inter3));
  inv1  gate2861(.a(s_331), .O(gate392inter4));
  nand2 gate2862(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2863(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2864(.a(G6), .O(gate392inter7));
  inv1  gate2865(.a(G1051), .O(gate392inter8));
  nand2 gate2866(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2867(.a(s_331), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2868(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2869(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2870(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1681(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1682(.a(gate394inter0), .b(s_162), .O(gate394inter1));
  and2  gate1683(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1684(.a(s_162), .O(gate394inter3));
  inv1  gate1685(.a(s_163), .O(gate394inter4));
  nand2 gate1686(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1687(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1688(.a(G8), .O(gate394inter7));
  inv1  gate1689(.a(G1057), .O(gate394inter8));
  nand2 gate1690(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1691(.a(s_163), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1692(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1693(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1694(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1331(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1332(.a(gate395inter0), .b(s_112), .O(gate395inter1));
  and2  gate1333(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1334(.a(s_112), .O(gate395inter3));
  inv1  gate1335(.a(s_113), .O(gate395inter4));
  nand2 gate1336(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1337(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1338(.a(G9), .O(gate395inter7));
  inv1  gate1339(.a(G1060), .O(gate395inter8));
  nand2 gate1340(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1341(.a(s_113), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1342(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1343(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1344(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2759(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2760(.a(gate396inter0), .b(s_316), .O(gate396inter1));
  and2  gate2761(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2762(.a(s_316), .O(gate396inter3));
  inv1  gate2763(.a(s_317), .O(gate396inter4));
  nand2 gate2764(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2765(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2766(.a(G10), .O(gate396inter7));
  inv1  gate2767(.a(G1063), .O(gate396inter8));
  nand2 gate2768(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2769(.a(s_317), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2770(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2771(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2772(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate2885(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2886(.a(gate397inter0), .b(s_334), .O(gate397inter1));
  and2  gate2887(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2888(.a(s_334), .O(gate397inter3));
  inv1  gate2889(.a(s_335), .O(gate397inter4));
  nand2 gate2890(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2891(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2892(.a(G11), .O(gate397inter7));
  inv1  gate2893(.a(G1066), .O(gate397inter8));
  nand2 gate2894(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2895(.a(s_335), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2896(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2897(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2898(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate3109(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate3110(.a(gate398inter0), .b(s_366), .O(gate398inter1));
  and2  gate3111(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate3112(.a(s_366), .O(gate398inter3));
  inv1  gate3113(.a(s_367), .O(gate398inter4));
  nand2 gate3114(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate3115(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate3116(.a(G12), .O(gate398inter7));
  inv1  gate3117(.a(G1069), .O(gate398inter8));
  nand2 gate3118(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate3119(.a(s_367), .b(gate398inter3), .O(gate398inter10));
  nor2  gate3120(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate3121(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate3122(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate2619(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2620(.a(gate399inter0), .b(s_296), .O(gate399inter1));
  and2  gate2621(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2622(.a(s_296), .O(gate399inter3));
  inv1  gate2623(.a(s_297), .O(gate399inter4));
  nand2 gate2624(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2625(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2626(.a(G13), .O(gate399inter7));
  inv1  gate2627(.a(G1072), .O(gate399inter8));
  nand2 gate2628(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2629(.a(s_297), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2630(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2631(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2632(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2185(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2186(.a(gate401inter0), .b(s_234), .O(gate401inter1));
  and2  gate2187(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2188(.a(s_234), .O(gate401inter3));
  inv1  gate2189(.a(s_235), .O(gate401inter4));
  nand2 gate2190(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2191(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2192(.a(G15), .O(gate401inter7));
  inv1  gate2193(.a(G1078), .O(gate401inter8));
  nand2 gate2194(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2195(.a(s_235), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2196(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2197(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2198(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate2465(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2466(.a(gate405inter0), .b(s_274), .O(gate405inter1));
  and2  gate2467(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2468(.a(s_274), .O(gate405inter3));
  inv1  gate2469(.a(s_275), .O(gate405inter4));
  nand2 gate2470(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2471(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2472(.a(G19), .O(gate405inter7));
  inv1  gate2473(.a(G1090), .O(gate405inter8));
  nand2 gate2474(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2475(.a(s_275), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2476(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2477(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2478(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2549(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2550(.a(gate407inter0), .b(s_286), .O(gate407inter1));
  and2  gate2551(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2552(.a(s_286), .O(gate407inter3));
  inv1  gate2553(.a(s_287), .O(gate407inter4));
  nand2 gate2554(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2555(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2556(.a(G21), .O(gate407inter7));
  inv1  gate2557(.a(G1096), .O(gate407inter8));
  nand2 gate2558(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2559(.a(s_287), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2560(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2561(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2562(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate575(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate576(.a(gate408inter0), .b(s_4), .O(gate408inter1));
  and2  gate577(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate578(.a(s_4), .O(gate408inter3));
  inv1  gate579(.a(s_5), .O(gate408inter4));
  nand2 gate580(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate581(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate582(.a(G22), .O(gate408inter7));
  inv1  gate583(.a(G1099), .O(gate408inter8));
  nand2 gate584(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate585(.a(s_5), .b(gate408inter3), .O(gate408inter10));
  nor2  gate586(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate587(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate588(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2437(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2438(.a(gate410inter0), .b(s_270), .O(gate410inter1));
  and2  gate2439(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2440(.a(s_270), .O(gate410inter3));
  inv1  gate2441(.a(s_271), .O(gate410inter4));
  nand2 gate2442(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2443(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2444(.a(G24), .O(gate410inter7));
  inv1  gate2445(.a(G1105), .O(gate410inter8));
  nand2 gate2446(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2447(.a(s_271), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2448(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2449(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2450(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2017(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2018(.a(gate413inter0), .b(s_210), .O(gate413inter1));
  and2  gate2019(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2020(.a(s_210), .O(gate413inter3));
  inv1  gate2021(.a(s_211), .O(gate413inter4));
  nand2 gate2022(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2023(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2024(.a(G27), .O(gate413inter7));
  inv1  gate2025(.a(G1114), .O(gate413inter8));
  nand2 gate2026(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2027(.a(s_211), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2028(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2029(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2030(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate981(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate982(.a(gate415inter0), .b(s_62), .O(gate415inter1));
  and2  gate983(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate984(.a(s_62), .O(gate415inter3));
  inv1  gate985(.a(s_63), .O(gate415inter4));
  nand2 gate986(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate987(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate988(.a(G29), .O(gate415inter7));
  inv1  gate989(.a(G1120), .O(gate415inter8));
  nand2 gate990(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate991(.a(s_63), .b(gate415inter3), .O(gate415inter10));
  nor2  gate992(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate993(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate994(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1947(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1948(.a(gate417inter0), .b(s_200), .O(gate417inter1));
  and2  gate1949(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1950(.a(s_200), .O(gate417inter3));
  inv1  gate1951(.a(s_201), .O(gate417inter4));
  nand2 gate1952(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1953(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1954(.a(G31), .O(gate417inter7));
  inv1  gate1955(.a(G1126), .O(gate417inter8));
  nand2 gate1956(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1957(.a(s_201), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1958(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1959(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1960(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2129(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2130(.a(gate420inter0), .b(s_226), .O(gate420inter1));
  and2  gate2131(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2132(.a(s_226), .O(gate420inter3));
  inv1  gate2133(.a(s_227), .O(gate420inter4));
  nand2 gate2134(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2135(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2136(.a(G1036), .O(gate420inter7));
  inv1  gate2137(.a(G1132), .O(gate420inter8));
  nand2 gate2138(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2139(.a(s_227), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2140(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2141(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2142(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2283(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2284(.a(gate423inter0), .b(s_248), .O(gate423inter1));
  and2  gate2285(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2286(.a(s_248), .O(gate423inter3));
  inv1  gate2287(.a(s_249), .O(gate423inter4));
  nand2 gate2288(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2289(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2290(.a(G3), .O(gate423inter7));
  inv1  gate2291(.a(G1138), .O(gate423inter8));
  nand2 gate2292(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2293(.a(s_249), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2294(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2295(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2296(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1975(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1976(.a(gate425inter0), .b(s_204), .O(gate425inter1));
  and2  gate1977(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1978(.a(s_204), .O(gate425inter3));
  inv1  gate1979(.a(s_205), .O(gate425inter4));
  nand2 gate1980(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1981(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1982(.a(G4), .O(gate425inter7));
  inv1  gate1983(.a(G1141), .O(gate425inter8));
  nand2 gate1984(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1985(.a(s_205), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1986(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1987(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1988(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2563(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2564(.a(gate430inter0), .b(s_288), .O(gate430inter1));
  and2  gate2565(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2566(.a(s_288), .O(gate430inter3));
  inv1  gate2567(.a(s_289), .O(gate430inter4));
  nand2 gate2568(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2569(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2570(.a(G1051), .O(gate430inter7));
  inv1  gate2571(.a(G1147), .O(gate430inter8));
  nand2 gate2572(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2573(.a(s_289), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2574(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2575(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2576(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1191(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1192(.a(gate432inter0), .b(s_92), .O(gate432inter1));
  and2  gate1193(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1194(.a(s_92), .O(gate432inter3));
  inv1  gate1195(.a(s_93), .O(gate432inter4));
  nand2 gate1196(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1197(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1198(.a(G1054), .O(gate432inter7));
  inv1  gate1199(.a(G1150), .O(gate432inter8));
  nand2 gate1200(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1201(.a(s_93), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1202(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1203(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1204(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1849(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1850(.a(gate433inter0), .b(s_186), .O(gate433inter1));
  and2  gate1851(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1852(.a(s_186), .O(gate433inter3));
  inv1  gate1853(.a(s_187), .O(gate433inter4));
  nand2 gate1854(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1855(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1856(.a(G8), .O(gate433inter7));
  inv1  gate1857(.a(G1153), .O(gate433inter8));
  nand2 gate1858(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1859(.a(s_187), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1860(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1861(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1862(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1807(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1808(.a(gate434inter0), .b(s_180), .O(gate434inter1));
  and2  gate1809(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1810(.a(s_180), .O(gate434inter3));
  inv1  gate1811(.a(s_181), .O(gate434inter4));
  nand2 gate1812(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1813(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1814(.a(G1057), .O(gate434inter7));
  inv1  gate1815(.a(G1153), .O(gate434inter8));
  nand2 gate1816(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1817(.a(s_181), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1818(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1819(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1820(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2591(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2592(.a(gate435inter0), .b(s_292), .O(gate435inter1));
  and2  gate2593(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2594(.a(s_292), .O(gate435inter3));
  inv1  gate2595(.a(s_293), .O(gate435inter4));
  nand2 gate2596(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2597(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2598(.a(G9), .O(gate435inter7));
  inv1  gate2599(.a(G1156), .O(gate435inter8));
  nand2 gate2600(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2601(.a(s_293), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2602(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2603(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2604(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate967(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate968(.a(gate436inter0), .b(s_60), .O(gate436inter1));
  and2  gate969(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate970(.a(s_60), .O(gate436inter3));
  inv1  gate971(.a(s_61), .O(gate436inter4));
  nand2 gate972(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate973(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate974(.a(G1060), .O(gate436inter7));
  inv1  gate975(.a(G1156), .O(gate436inter8));
  nand2 gate976(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate977(.a(s_61), .b(gate436inter3), .O(gate436inter10));
  nor2  gate978(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate979(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate980(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1583(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1584(.a(gate437inter0), .b(s_148), .O(gate437inter1));
  and2  gate1585(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1586(.a(s_148), .O(gate437inter3));
  inv1  gate1587(.a(s_149), .O(gate437inter4));
  nand2 gate1588(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1589(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1590(.a(G10), .O(gate437inter7));
  inv1  gate1591(.a(G1159), .O(gate437inter8));
  nand2 gate1592(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1593(.a(s_149), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1594(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1595(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1596(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2269(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2270(.a(gate438inter0), .b(s_246), .O(gate438inter1));
  and2  gate2271(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2272(.a(s_246), .O(gate438inter3));
  inv1  gate2273(.a(s_247), .O(gate438inter4));
  nand2 gate2274(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2275(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2276(.a(G1063), .O(gate438inter7));
  inv1  gate2277(.a(G1159), .O(gate438inter8));
  nand2 gate2278(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2279(.a(s_247), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2280(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2281(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2282(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1163(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1164(.a(gate440inter0), .b(s_88), .O(gate440inter1));
  and2  gate1165(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1166(.a(s_88), .O(gate440inter3));
  inv1  gate1167(.a(s_89), .O(gate440inter4));
  nand2 gate1168(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1169(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1170(.a(G1066), .O(gate440inter7));
  inv1  gate1171(.a(G1162), .O(gate440inter8));
  nand2 gate1172(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1173(.a(s_89), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1174(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1175(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1176(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2717(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2718(.a(gate442inter0), .b(s_310), .O(gate442inter1));
  and2  gate2719(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2720(.a(s_310), .O(gate442inter3));
  inv1  gate2721(.a(s_311), .O(gate442inter4));
  nand2 gate2722(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2723(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2724(.a(G1069), .O(gate442inter7));
  inv1  gate2725(.a(G1165), .O(gate442inter8));
  nand2 gate2726(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2727(.a(s_311), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2728(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2729(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2730(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1625(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1626(.a(gate445inter0), .b(s_154), .O(gate445inter1));
  and2  gate1627(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1628(.a(s_154), .O(gate445inter3));
  inv1  gate1629(.a(s_155), .O(gate445inter4));
  nand2 gate1630(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1631(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1632(.a(G14), .O(gate445inter7));
  inv1  gate1633(.a(G1171), .O(gate445inter8));
  nand2 gate1634(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1635(.a(s_155), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1636(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1637(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1638(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1821(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1822(.a(gate446inter0), .b(s_182), .O(gate446inter1));
  and2  gate1823(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1824(.a(s_182), .O(gate446inter3));
  inv1  gate1825(.a(s_183), .O(gate446inter4));
  nand2 gate1826(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1827(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1828(.a(G1075), .O(gate446inter7));
  inv1  gate1829(.a(G1171), .O(gate446inter8));
  nand2 gate1830(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1831(.a(s_183), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1832(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1833(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1834(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2507(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2508(.a(gate448inter0), .b(s_280), .O(gate448inter1));
  and2  gate2509(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2510(.a(s_280), .O(gate448inter3));
  inv1  gate2511(.a(s_281), .O(gate448inter4));
  nand2 gate2512(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2513(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2514(.a(G1078), .O(gate448inter7));
  inv1  gate2515(.a(G1174), .O(gate448inter8));
  nand2 gate2516(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2517(.a(s_281), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2518(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2519(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2520(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1457(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1458(.a(gate449inter0), .b(s_130), .O(gate449inter1));
  and2  gate1459(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1460(.a(s_130), .O(gate449inter3));
  inv1  gate1461(.a(s_131), .O(gate449inter4));
  nand2 gate1462(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1463(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1464(.a(G16), .O(gate449inter7));
  inv1  gate1465(.a(G1177), .O(gate449inter8));
  nand2 gate1466(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1467(.a(s_131), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1468(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1469(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1470(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate715(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate716(.a(gate450inter0), .b(s_24), .O(gate450inter1));
  and2  gate717(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate718(.a(s_24), .O(gate450inter3));
  inv1  gate719(.a(s_25), .O(gate450inter4));
  nand2 gate720(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate721(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate722(.a(G1081), .O(gate450inter7));
  inv1  gate723(.a(G1177), .O(gate450inter8));
  nand2 gate724(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate725(.a(s_25), .b(gate450inter3), .O(gate450inter10));
  nor2  gate726(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate727(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate728(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1933(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1934(.a(gate454inter0), .b(s_198), .O(gate454inter1));
  and2  gate1935(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1936(.a(s_198), .O(gate454inter3));
  inv1  gate1937(.a(s_199), .O(gate454inter4));
  nand2 gate1938(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1939(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1940(.a(G1087), .O(gate454inter7));
  inv1  gate1941(.a(G1183), .O(gate454inter8));
  nand2 gate1942(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1943(.a(s_199), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1944(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1945(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1946(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate2941(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2942(.a(gate455inter0), .b(s_342), .O(gate455inter1));
  and2  gate2943(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2944(.a(s_342), .O(gate455inter3));
  inv1  gate2945(.a(s_343), .O(gate455inter4));
  nand2 gate2946(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2947(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2948(.a(G19), .O(gate455inter7));
  inv1  gate2949(.a(G1186), .O(gate455inter8));
  nand2 gate2950(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2951(.a(s_343), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2952(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2953(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2954(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1275(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1276(.a(gate458inter0), .b(s_104), .O(gate458inter1));
  and2  gate1277(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1278(.a(s_104), .O(gate458inter3));
  inv1  gate1279(.a(s_105), .O(gate458inter4));
  nand2 gate1280(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1281(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1282(.a(G1093), .O(gate458inter7));
  inv1  gate1283(.a(G1189), .O(gate458inter8));
  nand2 gate1284(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1285(.a(s_105), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1286(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1287(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1288(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate2801(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2802(.a(gate459inter0), .b(s_322), .O(gate459inter1));
  and2  gate2803(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2804(.a(s_322), .O(gate459inter3));
  inv1  gate2805(.a(s_323), .O(gate459inter4));
  nand2 gate2806(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2807(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2808(.a(G21), .O(gate459inter7));
  inv1  gate2809(.a(G1192), .O(gate459inter8));
  nand2 gate2810(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2811(.a(s_323), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2812(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2813(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2814(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1233(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1234(.a(gate461inter0), .b(s_98), .O(gate461inter1));
  and2  gate1235(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1236(.a(s_98), .O(gate461inter3));
  inv1  gate1237(.a(s_99), .O(gate461inter4));
  nand2 gate1238(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1239(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1240(.a(G22), .O(gate461inter7));
  inv1  gate1241(.a(G1195), .O(gate461inter8));
  nand2 gate1242(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1243(.a(s_99), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1244(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1245(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1246(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate1667(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1668(.a(gate462inter0), .b(s_160), .O(gate462inter1));
  and2  gate1669(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1670(.a(s_160), .O(gate462inter3));
  inv1  gate1671(.a(s_161), .O(gate462inter4));
  nand2 gate1672(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1673(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1674(.a(G1099), .O(gate462inter7));
  inv1  gate1675(.a(G1195), .O(gate462inter8));
  nand2 gate1676(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1677(.a(s_161), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1678(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1679(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1680(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate897(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate898(.a(gate465inter0), .b(s_50), .O(gate465inter1));
  and2  gate899(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate900(.a(s_50), .O(gate465inter3));
  inv1  gate901(.a(s_51), .O(gate465inter4));
  nand2 gate902(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate903(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate904(.a(G24), .O(gate465inter7));
  inv1  gate905(.a(G1201), .O(gate465inter8));
  nand2 gate906(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate907(.a(s_51), .b(gate465inter3), .O(gate465inter10));
  nor2  gate908(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate909(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate910(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1289(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1290(.a(gate466inter0), .b(s_106), .O(gate466inter1));
  and2  gate1291(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1292(.a(s_106), .O(gate466inter3));
  inv1  gate1293(.a(s_107), .O(gate466inter4));
  nand2 gate1294(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1295(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1296(.a(G1105), .O(gate466inter7));
  inv1  gate1297(.a(G1201), .O(gate466inter8));
  nand2 gate1298(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1299(.a(s_107), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1300(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1301(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1302(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1499(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1500(.a(gate468inter0), .b(s_136), .O(gate468inter1));
  and2  gate1501(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1502(.a(s_136), .O(gate468inter3));
  inv1  gate1503(.a(s_137), .O(gate468inter4));
  nand2 gate1504(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1505(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1506(.a(G1108), .O(gate468inter7));
  inv1  gate1507(.a(G1204), .O(gate468inter8));
  nand2 gate1508(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1509(.a(s_137), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1510(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1511(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1512(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate1079(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1080(.a(gate469inter0), .b(s_76), .O(gate469inter1));
  and2  gate1081(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1082(.a(s_76), .O(gate469inter3));
  inv1  gate1083(.a(s_77), .O(gate469inter4));
  nand2 gate1084(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1085(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1086(.a(G26), .O(gate469inter7));
  inv1  gate1087(.a(G1207), .O(gate469inter8));
  nand2 gate1088(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1089(.a(s_77), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1090(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1091(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1092(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2059(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2060(.a(gate471inter0), .b(s_216), .O(gate471inter1));
  and2  gate2061(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2062(.a(s_216), .O(gate471inter3));
  inv1  gate2063(.a(s_217), .O(gate471inter4));
  nand2 gate2064(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2065(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2066(.a(G27), .O(gate471inter7));
  inv1  gate2067(.a(G1210), .O(gate471inter8));
  nand2 gate2068(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2069(.a(s_217), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2070(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2071(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2072(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1835(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1836(.a(gate476inter0), .b(s_184), .O(gate476inter1));
  and2  gate1837(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1838(.a(s_184), .O(gate476inter3));
  inv1  gate1839(.a(s_185), .O(gate476inter4));
  nand2 gate1840(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1841(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1842(.a(G1120), .O(gate476inter7));
  inv1  gate1843(.a(G1216), .O(gate476inter8));
  nand2 gate1844(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1845(.a(s_185), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1846(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1847(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1848(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1037(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1038(.a(gate479inter0), .b(s_70), .O(gate479inter1));
  and2  gate1039(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1040(.a(s_70), .O(gate479inter3));
  inv1  gate1041(.a(s_71), .O(gate479inter4));
  nand2 gate1042(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1043(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1044(.a(G31), .O(gate479inter7));
  inv1  gate1045(.a(G1222), .O(gate479inter8));
  nand2 gate1046(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1047(.a(s_71), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1048(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1049(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1050(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1177(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1178(.a(gate481inter0), .b(s_90), .O(gate481inter1));
  and2  gate1179(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1180(.a(s_90), .O(gate481inter3));
  inv1  gate1181(.a(s_91), .O(gate481inter4));
  nand2 gate1182(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1183(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1184(.a(G32), .O(gate481inter7));
  inv1  gate1185(.a(G1225), .O(gate481inter8));
  nand2 gate1186(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1187(.a(s_91), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1188(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1189(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1190(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1569(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1570(.a(gate482inter0), .b(s_146), .O(gate482inter1));
  and2  gate1571(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1572(.a(s_146), .O(gate482inter3));
  inv1  gate1573(.a(s_147), .O(gate482inter4));
  nand2 gate1574(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1575(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1576(.a(G1129), .O(gate482inter7));
  inv1  gate1577(.a(G1225), .O(gate482inter8));
  nand2 gate1578(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1579(.a(s_147), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1580(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1581(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1582(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate3039(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate3040(.a(gate486inter0), .b(s_356), .O(gate486inter1));
  and2  gate3041(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate3042(.a(s_356), .O(gate486inter3));
  inv1  gate3043(.a(s_357), .O(gate486inter4));
  nand2 gate3044(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate3045(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate3046(.a(G1234), .O(gate486inter7));
  inv1  gate3047(.a(G1235), .O(gate486inter8));
  nand2 gate3048(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate3049(.a(s_357), .b(gate486inter3), .O(gate486inter10));
  nor2  gate3050(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate3051(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate3052(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1639(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1640(.a(gate487inter0), .b(s_156), .O(gate487inter1));
  and2  gate1641(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1642(.a(s_156), .O(gate487inter3));
  inv1  gate1643(.a(s_157), .O(gate487inter4));
  nand2 gate1644(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1645(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1646(.a(G1236), .O(gate487inter7));
  inv1  gate1647(.a(G1237), .O(gate487inter8));
  nand2 gate1648(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1649(.a(s_157), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1650(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1651(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1652(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1597(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1598(.a(gate488inter0), .b(s_150), .O(gate488inter1));
  and2  gate1599(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1600(.a(s_150), .O(gate488inter3));
  inv1  gate1601(.a(s_151), .O(gate488inter4));
  nand2 gate1602(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1603(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1604(.a(G1238), .O(gate488inter7));
  inv1  gate1605(.a(G1239), .O(gate488inter8));
  nand2 gate1606(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1607(.a(s_151), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1608(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1609(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1610(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2535(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2536(.a(gate492inter0), .b(s_284), .O(gate492inter1));
  and2  gate2537(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2538(.a(s_284), .O(gate492inter3));
  inv1  gate2539(.a(s_285), .O(gate492inter4));
  nand2 gate2540(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2541(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2542(.a(G1246), .O(gate492inter7));
  inv1  gate2543(.a(G1247), .O(gate492inter8));
  nand2 gate2544(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2545(.a(s_285), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2546(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2547(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2548(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1303(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1304(.a(gate493inter0), .b(s_108), .O(gate493inter1));
  and2  gate1305(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1306(.a(s_108), .O(gate493inter3));
  inv1  gate1307(.a(s_109), .O(gate493inter4));
  nand2 gate1308(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1309(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1310(.a(G1248), .O(gate493inter7));
  inv1  gate1311(.a(G1249), .O(gate493inter8));
  nand2 gate1312(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1313(.a(s_109), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1314(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1315(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1316(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate3067(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate3068(.a(gate495inter0), .b(s_360), .O(gate495inter1));
  and2  gate3069(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate3070(.a(s_360), .O(gate495inter3));
  inv1  gate3071(.a(s_361), .O(gate495inter4));
  nand2 gate3072(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate3073(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate3074(.a(G1252), .O(gate495inter7));
  inv1  gate3075(.a(G1253), .O(gate495inter8));
  nand2 gate3076(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate3077(.a(s_361), .b(gate495inter3), .O(gate495inter10));
  nor2  gate3078(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate3079(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate3080(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate953(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate954(.a(gate498inter0), .b(s_58), .O(gate498inter1));
  and2  gate955(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate956(.a(s_58), .O(gate498inter3));
  inv1  gate957(.a(s_59), .O(gate498inter4));
  nand2 gate958(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate959(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate960(.a(G1258), .O(gate498inter7));
  inv1  gate961(.a(G1259), .O(gate498inter8));
  nand2 gate962(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate963(.a(s_59), .b(gate498inter3), .O(gate498inter10));
  nor2  gate964(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate965(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate966(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1121(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1122(.a(gate499inter0), .b(s_82), .O(gate499inter1));
  and2  gate1123(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1124(.a(s_82), .O(gate499inter3));
  inv1  gate1125(.a(s_83), .O(gate499inter4));
  nand2 gate1126(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1127(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1128(.a(G1260), .O(gate499inter7));
  inv1  gate1129(.a(G1261), .O(gate499inter8));
  nand2 gate1130(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1131(.a(s_83), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1132(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1133(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1134(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2311(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2312(.a(gate503inter0), .b(s_252), .O(gate503inter1));
  and2  gate2313(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2314(.a(s_252), .O(gate503inter3));
  inv1  gate2315(.a(s_253), .O(gate503inter4));
  nand2 gate2316(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2317(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2318(.a(G1268), .O(gate503inter7));
  inv1  gate2319(.a(G1269), .O(gate503inter8));
  nand2 gate2320(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2321(.a(s_253), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2322(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2323(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2324(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate547(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate548(.a(gate505inter0), .b(s_0), .O(gate505inter1));
  and2  gate549(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate550(.a(s_0), .O(gate505inter3));
  inv1  gate551(.a(s_1), .O(gate505inter4));
  nand2 gate552(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate553(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate554(.a(G1272), .O(gate505inter7));
  inv1  gate555(.a(G1273), .O(gate505inter8));
  nand2 gate556(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate557(.a(s_1), .b(gate505inter3), .O(gate505inter10));
  nor2  gate558(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate559(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate560(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2493(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2494(.a(gate507inter0), .b(s_278), .O(gate507inter1));
  and2  gate2495(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2496(.a(s_278), .O(gate507inter3));
  inv1  gate2497(.a(s_279), .O(gate507inter4));
  nand2 gate2498(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2499(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2500(.a(G1276), .O(gate507inter7));
  inv1  gate2501(.a(G1277), .O(gate507inter8));
  nand2 gate2502(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2503(.a(s_279), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2504(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2505(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2506(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate827(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate828(.a(gate509inter0), .b(s_40), .O(gate509inter1));
  and2  gate829(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate830(.a(s_40), .O(gate509inter3));
  inv1  gate831(.a(s_41), .O(gate509inter4));
  nand2 gate832(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate833(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate834(.a(G1280), .O(gate509inter7));
  inv1  gate835(.a(G1281), .O(gate509inter8));
  nand2 gate836(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate837(.a(s_41), .b(gate509inter3), .O(gate509inter10));
  nor2  gate838(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate839(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate840(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate925(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate926(.a(gate511inter0), .b(s_54), .O(gate511inter1));
  and2  gate927(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate928(.a(s_54), .O(gate511inter3));
  inv1  gate929(.a(s_55), .O(gate511inter4));
  nand2 gate930(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate931(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate932(.a(G1284), .O(gate511inter7));
  inv1  gate933(.a(G1285), .O(gate511inter8));
  nand2 gate934(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate935(.a(s_55), .b(gate511inter3), .O(gate511inter10));
  nor2  gate936(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate937(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate938(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule