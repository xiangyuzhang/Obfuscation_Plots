module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate3179(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate3180(.a(gate12inter0), .b(s_376), .O(gate12inter1));
  and2  gate3181(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate3182(.a(s_376), .O(gate12inter3));
  inv1  gate3183(.a(s_377), .O(gate12inter4));
  nand2 gate3184(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate3185(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate3186(.a(G7), .O(gate12inter7));
  inv1  gate3187(.a(G8), .O(gate12inter8));
  nand2 gate3188(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate3189(.a(s_377), .b(gate12inter3), .O(gate12inter10));
  nor2  gate3190(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate3191(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate3192(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1051(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1052(.a(gate13inter0), .b(s_72), .O(gate13inter1));
  and2  gate1053(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1054(.a(s_72), .O(gate13inter3));
  inv1  gate1055(.a(s_73), .O(gate13inter4));
  nand2 gate1056(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1057(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1058(.a(G9), .O(gate13inter7));
  inv1  gate1059(.a(G10), .O(gate13inter8));
  nand2 gate1060(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1061(.a(s_73), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1062(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1063(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1064(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1387(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1388(.a(gate14inter0), .b(s_120), .O(gate14inter1));
  and2  gate1389(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1390(.a(s_120), .O(gate14inter3));
  inv1  gate1391(.a(s_121), .O(gate14inter4));
  nand2 gate1392(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1393(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1394(.a(G11), .O(gate14inter7));
  inv1  gate1395(.a(G12), .O(gate14inter8));
  nand2 gate1396(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1397(.a(s_121), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1398(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1399(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1400(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1093(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1094(.a(gate16inter0), .b(s_78), .O(gate16inter1));
  and2  gate1095(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1096(.a(s_78), .O(gate16inter3));
  inv1  gate1097(.a(s_79), .O(gate16inter4));
  nand2 gate1098(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1099(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1100(.a(G15), .O(gate16inter7));
  inv1  gate1101(.a(G16), .O(gate16inter8));
  nand2 gate1102(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1103(.a(s_79), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1104(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1105(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1106(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate771(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate772(.a(gate17inter0), .b(s_32), .O(gate17inter1));
  and2  gate773(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate774(.a(s_32), .O(gate17inter3));
  inv1  gate775(.a(s_33), .O(gate17inter4));
  nand2 gate776(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate777(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate778(.a(G17), .O(gate17inter7));
  inv1  gate779(.a(G18), .O(gate17inter8));
  nand2 gate780(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate781(.a(s_33), .b(gate17inter3), .O(gate17inter10));
  nor2  gate782(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate783(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate784(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2241(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2242(.a(gate19inter0), .b(s_242), .O(gate19inter1));
  and2  gate2243(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2244(.a(s_242), .O(gate19inter3));
  inv1  gate2245(.a(s_243), .O(gate19inter4));
  nand2 gate2246(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2247(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2248(.a(G21), .O(gate19inter7));
  inv1  gate2249(.a(G22), .O(gate19inter8));
  nand2 gate2250(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2251(.a(s_243), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2252(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2253(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2254(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate3207(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate3208(.a(gate21inter0), .b(s_380), .O(gate21inter1));
  and2  gate3209(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate3210(.a(s_380), .O(gate21inter3));
  inv1  gate3211(.a(s_381), .O(gate21inter4));
  nand2 gate3212(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate3213(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate3214(.a(G25), .O(gate21inter7));
  inv1  gate3215(.a(G26), .O(gate21inter8));
  nand2 gate3216(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate3217(.a(s_381), .b(gate21inter3), .O(gate21inter10));
  nor2  gate3218(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate3219(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate3220(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2941(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2942(.a(gate22inter0), .b(s_342), .O(gate22inter1));
  and2  gate2943(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2944(.a(s_342), .O(gate22inter3));
  inv1  gate2945(.a(s_343), .O(gate22inter4));
  nand2 gate2946(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2947(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2948(.a(G27), .O(gate22inter7));
  inv1  gate2949(.a(G28), .O(gate22inter8));
  nand2 gate2950(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2951(.a(s_343), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2952(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2953(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2954(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2913(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2914(.a(gate23inter0), .b(s_338), .O(gate23inter1));
  and2  gate2915(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2916(.a(s_338), .O(gate23inter3));
  inv1  gate2917(.a(s_339), .O(gate23inter4));
  nand2 gate2918(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2919(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2920(.a(G29), .O(gate23inter7));
  inv1  gate2921(.a(G30), .O(gate23inter8));
  nand2 gate2922(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2923(.a(s_339), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2924(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2925(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2926(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate673(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate674(.a(gate24inter0), .b(s_18), .O(gate24inter1));
  and2  gate675(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate676(.a(s_18), .O(gate24inter3));
  inv1  gate677(.a(s_19), .O(gate24inter4));
  nand2 gate678(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate679(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate680(.a(G31), .O(gate24inter7));
  inv1  gate681(.a(G32), .O(gate24inter8));
  nand2 gate682(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate683(.a(s_19), .b(gate24inter3), .O(gate24inter10));
  nor2  gate684(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate685(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate686(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate813(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate814(.a(gate27inter0), .b(s_38), .O(gate27inter1));
  and2  gate815(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate816(.a(s_38), .O(gate27inter3));
  inv1  gate817(.a(s_39), .O(gate27inter4));
  nand2 gate818(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate819(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate820(.a(G2), .O(gate27inter7));
  inv1  gate821(.a(G6), .O(gate27inter8));
  nand2 gate822(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate823(.a(s_39), .b(gate27inter3), .O(gate27inter10));
  nor2  gate824(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate825(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate826(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2535(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2536(.a(gate29inter0), .b(s_284), .O(gate29inter1));
  and2  gate2537(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2538(.a(s_284), .O(gate29inter3));
  inv1  gate2539(.a(s_285), .O(gate29inter4));
  nand2 gate2540(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2541(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2542(.a(G3), .O(gate29inter7));
  inv1  gate2543(.a(G7), .O(gate29inter8));
  nand2 gate2544(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2545(.a(s_285), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2546(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2547(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2548(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2787(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2788(.a(gate30inter0), .b(s_320), .O(gate30inter1));
  and2  gate2789(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2790(.a(s_320), .O(gate30inter3));
  inv1  gate2791(.a(s_321), .O(gate30inter4));
  nand2 gate2792(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2793(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2794(.a(G11), .O(gate30inter7));
  inv1  gate2795(.a(G15), .O(gate30inter8));
  nand2 gate2796(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2797(.a(s_321), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2798(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2799(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2800(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2857(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2858(.a(gate32inter0), .b(s_330), .O(gate32inter1));
  and2  gate2859(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2860(.a(s_330), .O(gate32inter3));
  inv1  gate2861(.a(s_331), .O(gate32inter4));
  nand2 gate2862(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2863(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2864(.a(G12), .O(gate32inter7));
  inv1  gate2865(.a(G16), .O(gate32inter8));
  nand2 gate2866(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2867(.a(s_331), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2868(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2869(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2870(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1037(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1038(.a(gate34inter0), .b(s_70), .O(gate34inter1));
  and2  gate1039(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1040(.a(s_70), .O(gate34inter3));
  inv1  gate1041(.a(s_71), .O(gate34inter4));
  nand2 gate1042(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1043(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1044(.a(G25), .O(gate34inter7));
  inv1  gate1045(.a(G29), .O(gate34inter8));
  nand2 gate1046(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1047(.a(s_71), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1048(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1049(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1050(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2605(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2606(.a(gate38inter0), .b(s_294), .O(gate38inter1));
  and2  gate2607(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2608(.a(s_294), .O(gate38inter3));
  inv1  gate2609(.a(s_295), .O(gate38inter4));
  nand2 gate2610(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2611(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2612(.a(G27), .O(gate38inter7));
  inv1  gate2613(.a(G31), .O(gate38inter8));
  nand2 gate2614(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2615(.a(s_295), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2616(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2617(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2618(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate729(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate730(.a(gate39inter0), .b(s_26), .O(gate39inter1));
  and2  gate731(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate732(.a(s_26), .O(gate39inter3));
  inv1  gate733(.a(s_27), .O(gate39inter4));
  nand2 gate734(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate735(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate736(.a(G20), .O(gate39inter7));
  inv1  gate737(.a(G24), .O(gate39inter8));
  nand2 gate738(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate739(.a(s_27), .b(gate39inter3), .O(gate39inter10));
  nor2  gate740(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate741(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate742(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1331(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1332(.a(gate42inter0), .b(s_112), .O(gate42inter1));
  and2  gate1333(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1334(.a(s_112), .O(gate42inter3));
  inv1  gate1335(.a(s_113), .O(gate42inter4));
  nand2 gate1336(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1337(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1338(.a(G2), .O(gate42inter7));
  inv1  gate1339(.a(G266), .O(gate42inter8));
  nand2 gate1340(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1341(.a(s_113), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1342(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1343(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1344(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1555(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1556(.a(gate44inter0), .b(s_144), .O(gate44inter1));
  and2  gate1557(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1558(.a(s_144), .O(gate44inter3));
  inv1  gate1559(.a(s_145), .O(gate44inter4));
  nand2 gate1560(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1561(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1562(.a(G4), .O(gate44inter7));
  inv1  gate1563(.a(G269), .O(gate44inter8));
  nand2 gate1564(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1565(.a(s_145), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1566(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1567(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1568(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2563(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2564(.a(gate45inter0), .b(s_288), .O(gate45inter1));
  and2  gate2565(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2566(.a(s_288), .O(gate45inter3));
  inv1  gate2567(.a(s_289), .O(gate45inter4));
  nand2 gate2568(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2569(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2570(.a(G5), .O(gate45inter7));
  inv1  gate2571(.a(G272), .O(gate45inter8));
  nand2 gate2572(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2573(.a(s_289), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2574(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2575(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2576(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1891(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1892(.a(gate46inter0), .b(s_192), .O(gate46inter1));
  and2  gate1893(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1894(.a(s_192), .O(gate46inter3));
  inv1  gate1895(.a(s_193), .O(gate46inter4));
  nand2 gate1896(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1897(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1898(.a(G6), .O(gate46inter7));
  inv1  gate1899(.a(G272), .O(gate46inter8));
  nand2 gate1900(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1901(.a(s_193), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1902(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1903(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1904(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1527(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1528(.a(gate50inter0), .b(s_140), .O(gate50inter1));
  and2  gate1529(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1530(.a(s_140), .O(gate50inter3));
  inv1  gate1531(.a(s_141), .O(gate50inter4));
  nand2 gate1532(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1533(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1534(.a(G10), .O(gate50inter7));
  inv1  gate1535(.a(G278), .O(gate50inter8));
  nand2 gate1536(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1537(.a(s_141), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1538(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1539(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1540(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1023(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1024(.a(gate51inter0), .b(s_68), .O(gate51inter1));
  and2  gate1025(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1026(.a(s_68), .O(gate51inter3));
  inv1  gate1027(.a(s_69), .O(gate51inter4));
  nand2 gate1028(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1029(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1030(.a(G11), .O(gate51inter7));
  inv1  gate1031(.a(G281), .O(gate51inter8));
  nand2 gate1032(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1033(.a(s_69), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1034(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1035(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1036(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2129(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2130(.a(gate53inter0), .b(s_226), .O(gate53inter1));
  and2  gate2131(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2132(.a(s_226), .O(gate53inter3));
  inv1  gate2133(.a(s_227), .O(gate53inter4));
  nand2 gate2134(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2135(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2136(.a(G13), .O(gate53inter7));
  inv1  gate2137(.a(G284), .O(gate53inter8));
  nand2 gate2138(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2139(.a(s_227), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2140(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2141(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2142(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate631(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate632(.a(gate54inter0), .b(s_12), .O(gate54inter1));
  and2  gate633(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate634(.a(s_12), .O(gate54inter3));
  inv1  gate635(.a(s_13), .O(gate54inter4));
  nand2 gate636(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate637(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate638(.a(G14), .O(gate54inter7));
  inv1  gate639(.a(G284), .O(gate54inter8));
  nand2 gate640(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate641(.a(s_13), .b(gate54inter3), .O(gate54inter10));
  nor2  gate642(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate643(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate644(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate3095(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate3096(.a(gate57inter0), .b(s_364), .O(gate57inter1));
  and2  gate3097(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate3098(.a(s_364), .O(gate57inter3));
  inv1  gate3099(.a(s_365), .O(gate57inter4));
  nand2 gate3100(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate3101(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate3102(.a(G17), .O(gate57inter7));
  inv1  gate3103(.a(G290), .O(gate57inter8));
  nand2 gate3104(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate3105(.a(s_365), .b(gate57inter3), .O(gate57inter10));
  nor2  gate3106(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate3107(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate3108(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1009(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1010(.a(gate59inter0), .b(s_66), .O(gate59inter1));
  and2  gate1011(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1012(.a(s_66), .O(gate59inter3));
  inv1  gate1013(.a(s_67), .O(gate59inter4));
  nand2 gate1014(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1015(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1016(.a(G19), .O(gate59inter7));
  inv1  gate1017(.a(G293), .O(gate59inter8));
  nand2 gate1018(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1019(.a(s_67), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1020(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1021(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1022(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate2885(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2886(.a(gate60inter0), .b(s_334), .O(gate60inter1));
  and2  gate2887(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2888(.a(s_334), .O(gate60inter3));
  inv1  gate2889(.a(s_335), .O(gate60inter4));
  nand2 gate2890(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2891(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2892(.a(G20), .O(gate60inter7));
  inv1  gate2893(.a(G293), .O(gate60inter8));
  nand2 gate2894(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2895(.a(s_335), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2896(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2897(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2898(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2969(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2970(.a(gate61inter0), .b(s_346), .O(gate61inter1));
  and2  gate2971(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2972(.a(s_346), .O(gate61inter3));
  inv1  gate2973(.a(s_347), .O(gate61inter4));
  nand2 gate2974(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2975(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2976(.a(G21), .O(gate61inter7));
  inv1  gate2977(.a(G296), .O(gate61inter8));
  nand2 gate2978(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2979(.a(s_347), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2980(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2981(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2982(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2815(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2816(.a(gate64inter0), .b(s_324), .O(gate64inter1));
  and2  gate2817(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2818(.a(s_324), .O(gate64inter3));
  inv1  gate2819(.a(s_325), .O(gate64inter4));
  nand2 gate2820(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2821(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2822(.a(G24), .O(gate64inter7));
  inv1  gate2823(.a(G299), .O(gate64inter8));
  nand2 gate2824(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2825(.a(s_325), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2826(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2827(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2828(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1695(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1696(.a(gate67inter0), .b(s_164), .O(gate67inter1));
  and2  gate1697(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1698(.a(s_164), .O(gate67inter3));
  inv1  gate1699(.a(s_165), .O(gate67inter4));
  nand2 gate1700(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1701(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1702(.a(G27), .O(gate67inter7));
  inv1  gate1703(.a(G305), .O(gate67inter8));
  nand2 gate1704(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1705(.a(s_165), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1706(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1707(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1708(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate2647(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2648(.a(gate68inter0), .b(s_300), .O(gate68inter1));
  and2  gate2649(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2650(.a(s_300), .O(gate68inter3));
  inv1  gate2651(.a(s_301), .O(gate68inter4));
  nand2 gate2652(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2653(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2654(.a(G28), .O(gate68inter7));
  inv1  gate2655(.a(G305), .O(gate68inter8));
  nand2 gate2656(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2657(.a(s_301), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2658(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2659(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2660(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate701(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate702(.a(gate69inter0), .b(s_22), .O(gate69inter1));
  and2  gate703(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate704(.a(s_22), .O(gate69inter3));
  inv1  gate705(.a(s_23), .O(gate69inter4));
  nand2 gate706(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate707(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate708(.a(G29), .O(gate69inter7));
  inv1  gate709(.a(G308), .O(gate69inter8));
  nand2 gate710(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate711(.a(s_23), .b(gate69inter3), .O(gate69inter10));
  nor2  gate712(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate713(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate714(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1807(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1808(.a(gate70inter0), .b(s_180), .O(gate70inter1));
  and2  gate1809(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1810(.a(s_180), .O(gate70inter3));
  inv1  gate1811(.a(s_181), .O(gate70inter4));
  nand2 gate1812(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1813(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1814(.a(G30), .O(gate70inter7));
  inv1  gate1815(.a(G308), .O(gate70inter8));
  nand2 gate1816(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1817(.a(s_181), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1818(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1819(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1820(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1541(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1542(.a(gate77inter0), .b(s_142), .O(gate77inter1));
  and2  gate1543(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1544(.a(s_142), .O(gate77inter3));
  inv1  gate1545(.a(s_143), .O(gate77inter4));
  nand2 gate1546(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1547(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1548(.a(G2), .O(gate77inter7));
  inv1  gate1549(.a(G320), .O(gate77inter8));
  nand2 gate1550(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1551(.a(s_143), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1552(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1553(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1554(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1429(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1430(.a(gate79inter0), .b(s_126), .O(gate79inter1));
  and2  gate1431(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1432(.a(s_126), .O(gate79inter3));
  inv1  gate1433(.a(s_127), .O(gate79inter4));
  nand2 gate1434(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1435(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1436(.a(G10), .O(gate79inter7));
  inv1  gate1437(.a(G323), .O(gate79inter8));
  nand2 gate1438(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1439(.a(s_127), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1440(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1441(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1442(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2437(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2438(.a(gate85inter0), .b(s_270), .O(gate85inter1));
  and2  gate2439(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2440(.a(s_270), .O(gate85inter3));
  inv1  gate2441(.a(s_271), .O(gate85inter4));
  nand2 gate2442(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2443(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2444(.a(G4), .O(gate85inter7));
  inv1  gate2445(.a(G332), .O(gate85inter8));
  nand2 gate2446(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2447(.a(s_271), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2448(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2449(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2450(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1653(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1654(.a(gate87inter0), .b(s_158), .O(gate87inter1));
  and2  gate1655(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1656(.a(s_158), .O(gate87inter3));
  inv1  gate1657(.a(s_159), .O(gate87inter4));
  nand2 gate1658(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1659(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1660(.a(G12), .O(gate87inter7));
  inv1  gate1661(.a(G335), .O(gate87inter8));
  nand2 gate1662(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1663(.a(s_159), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1664(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1665(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1666(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1065(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1066(.a(gate88inter0), .b(s_74), .O(gate88inter1));
  and2  gate1067(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1068(.a(s_74), .O(gate88inter3));
  inv1  gate1069(.a(s_75), .O(gate88inter4));
  nand2 gate1070(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1071(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1072(.a(G16), .O(gate88inter7));
  inv1  gate1073(.a(G335), .O(gate88inter8));
  nand2 gate1074(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1075(.a(s_75), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1076(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1077(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1078(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1177(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1178(.a(gate94inter0), .b(s_90), .O(gate94inter1));
  and2  gate1179(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1180(.a(s_90), .O(gate94inter3));
  inv1  gate1181(.a(s_91), .O(gate94inter4));
  nand2 gate1182(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1183(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1184(.a(G22), .O(gate94inter7));
  inv1  gate1185(.a(G344), .O(gate94inter8));
  nand2 gate1186(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1187(.a(s_91), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1188(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1189(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1190(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1947(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1948(.a(gate97inter0), .b(s_200), .O(gate97inter1));
  and2  gate1949(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1950(.a(s_200), .O(gate97inter3));
  inv1  gate1951(.a(s_201), .O(gate97inter4));
  nand2 gate1952(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1953(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1954(.a(G19), .O(gate97inter7));
  inv1  gate1955(.a(G350), .O(gate97inter8));
  nand2 gate1956(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1957(.a(s_201), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1958(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1959(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1960(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate3081(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate3082(.a(gate98inter0), .b(s_362), .O(gate98inter1));
  and2  gate3083(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate3084(.a(s_362), .O(gate98inter3));
  inv1  gate3085(.a(s_363), .O(gate98inter4));
  nand2 gate3086(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate3087(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate3088(.a(G23), .O(gate98inter7));
  inv1  gate3089(.a(G350), .O(gate98inter8));
  nand2 gate3090(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate3091(.a(s_363), .b(gate98inter3), .O(gate98inter10));
  nor2  gate3092(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate3093(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate3094(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2367(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2368(.a(gate100inter0), .b(s_260), .O(gate100inter1));
  and2  gate2369(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2370(.a(s_260), .O(gate100inter3));
  inv1  gate2371(.a(s_261), .O(gate100inter4));
  nand2 gate2372(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2373(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2374(.a(G31), .O(gate100inter7));
  inv1  gate2375(.a(G353), .O(gate100inter8));
  nand2 gate2376(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2377(.a(s_261), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2378(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2379(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2380(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1289(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1290(.a(gate101inter0), .b(s_106), .O(gate101inter1));
  and2  gate1291(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1292(.a(s_106), .O(gate101inter3));
  inv1  gate1293(.a(s_107), .O(gate101inter4));
  nand2 gate1294(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1295(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1296(.a(G20), .O(gate101inter7));
  inv1  gate1297(.a(G356), .O(gate101inter8));
  nand2 gate1298(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1299(.a(s_107), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1300(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1301(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1302(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1149(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1150(.a(gate102inter0), .b(s_86), .O(gate102inter1));
  and2  gate1151(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1152(.a(s_86), .O(gate102inter3));
  inv1  gate1153(.a(s_87), .O(gate102inter4));
  nand2 gate1154(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1155(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1156(.a(G24), .O(gate102inter7));
  inv1  gate1157(.a(G356), .O(gate102inter8));
  nand2 gate1158(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1159(.a(s_87), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1160(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1161(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1162(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate953(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate954(.a(gate104inter0), .b(s_58), .O(gate104inter1));
  and2  gate955(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate956(.a(s_58), .O(gate104inter3));
  inv1  gate957(.a(s_59), .O(gate104inter4));
  nand2 gate958(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate959(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate960(.a(G32), .O(gate104inter7));
  inv1  gate961(.a(G359), .O(gate104inter8));
  nand2 gate962(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate963(.a(s_59), .b(gate104inter3), .O(gate104inter10));
  nor2  gate964(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate965(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate966(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate2549(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2550(.a(gate105inter0), .b(s_286), .O(gate105inter1));
  and2  gate2551(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2552(.a(s_286), .O(gate105inter3));
  inv1  gate2553(.a(s_287), .O(gate105inter4));
  nand2 gate2554(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2555(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2556(.a(G362), .O(gate105inter7));
  inv1  gate2557(.a(G363), .O(gate105inter8));
  nand2 gate2558(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2559(.a(s_287), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2560(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2561(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2562(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate3151(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate3152(.a(gate107inter0), .b(s_372), .O(gate107inter1));
  and2  gate3153(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate3154(.a(s_372), .O(gate107inter3));
  inv1  gate3155(.a(s_373), .O(gate107inter4));
  nand2 gate3156(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate3157(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate3158(.a(G366), .O(gate107inter7));
  inv1  gate3159(.a(G367), .O(gate107inter8));
  nand2 gate3160(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate3161(.a(s_373), .b(gate107inter3), .O(gate107inter10));
  nor2  gate3162(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate3163(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate3164(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate981(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate982(.a(gate109inter0), .b(s_62), .O(gate109inter1));
  and2  gate983(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate984(.a(s_62), .O(gate109inter3));
  inv1  gate985(.a(s_63), .O(gate109inter4));
  nand2 gate986(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate987(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate988(.a(G370), .O(gate109inter7));
  inv1  gate989(.a(G371), .O(gate109inter8));
  nand2 gate990(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate991(.a(s_63), .b(gate109inter3), .O(gate109inter10));
  nor2  gate992(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate993(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate994(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1779(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1780(.a(gate110inter0), .b(s_176), .O(gate110inter1));
  and2  gate1781(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1782(.a(s_176), .O(gate110inter3));
  inv1  gate1783(.a(s_177), .O(gate110inter4));
  nand2 gate1784(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1785(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1786(.a(G372), .O(gate110inter7));
  inv1  gate1787(.a(G373), .O(gate110inter8));
  nand2 gate1788(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1789(.a(s_177), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1790(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1791(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1792(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2801(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2802(.a(gate111inter0), .b(s_322), .O(gate111inter1));
  and2  gate2803(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2804(.a(s_322), .O(gate111inter3));
  inv1  gate2805(.a(s_323), .O(gate111inter4));
  nand2 gate2806(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2807(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2808(.a(G374), .O(gate111inter7));
  inv1  gate2809(.a(G375), .O(gate111inter8));
  nand2 gate2810(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2811(.a(s_323), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2812(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2813(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2814(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2675(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2676(.a(gate119inter0), .b(s_304), .O(gate119inter1));
  and2  gate2677(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2678(.a(s_304), .O(gate119inter3));
  inv1  gate2679(.a(s_305), .O(gate119inter4));
  nand2 gate2680(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2681(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2682(.a(G390), .O(gate119inter7));
  inv1  gate2683(.a(G391), .O(gate119inter8));
  nand2 gate2684(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2685(.a(s_305), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2686(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2687(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2688(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1765(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1766(.a(gate124inter0), .b(s_174), .O(gate124inter1));
  and2  gate1767(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1768(.a(s_174), .O(gate124inter3));
  inv1  gate1769(.a(s_175), .O(gate124inter4));
  nand2 gate1770(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1771(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1772(.a(G400), .O(gate124inter7));
  inv1  gate1773(.a(G401), .O(gate124inter8));
  nand2 gate1774(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1775(.a(s_175), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1776(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1777(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1778(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate967(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate968(.a(gate125inter0), .b(s_60), .O(gate125inter1));
  and2  gate969(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate970(.a(s_60), .O(gate125inter3));
  inv1  gate971(.a(s_61), .O(gate125inter4));
  nand2 gate972(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate973(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate974(.a(G402), .O(gate125inter7));
  inv1  gate975(.a(G403), .O(gate125inter8));
  nand2 gate976(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate977(.a(s_61), .b(gate125inter3), .O(gate125inter10));
  nor2  gate978(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate979(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate980(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1121(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1122(.a(gate126inter0), .b(s_82), .O(gate126inter1));
  and2  gate1123(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1124(.a(s_82), .O(gate126inter3));
  inv1  gate1125(.a(s_83), .O(gate126inter4));
  nand2 gate1126(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1127(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1128(.a(G404), .O(gate126inter7));
  inv1  gate1129(.a(G405), .O(gate126inter8));
  nand2 gate1130(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1131(.a(s_83), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1132(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1133(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1134(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1219(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1220(.a(gate128inter0), .b(s_96), .O(gate128inter1));
  and2  gate1221(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1222(.a(s_96), .O(gate128inter3));
  inv1  gate1223(.a(s_97), .O(gate128inter4));
  nand2 gate1224(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1225(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1226(.a(G408), .O(gate128inter7));
  inv1  gate1227(.a(G409), .O(gate128inter8));
  nand2 gate1228(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1229(.a(s_97), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1230(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1231(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1232(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate575(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate576(.a(gate129inter0), .b(s_4), .O(gate129inter1));
  and2  gate577(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate578(.a(s_4), .O(gate129inter3));
  inv1  gate579(.a(s_5), .O(gate129inter4));
  nand2 gate580(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate581(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate582(.a(G410), .O(gate129inter7));
  inv1  gate583(.a(G411), .O(gate129inter8));
  nand2 gate584(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate585(.a(s_5), .b(gate129inter3), .O(gate129inter10));
  nor2  gate586(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate587(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate588(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate1597(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1598(.a(gate130inter0), .b(s_150), .O(gate130inter1));
  and2  gate1599(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1600(.a(s_150), .O(gate130inter3));
  inv1  gate1601(.a(s_151), .O(gate130inter4));
  nand2 gate1602(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1603(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1604(.a(G412), .O(gate130inter7));
  inv1  gate1605(.a(G413), .O(gate130inter8));
  nand2 gate1606(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1607(.a(s_151), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1608(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1609(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1610(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate3109(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate3110(.a(gate131inter0), .b(s_366), .O(gate131inter1));
  and2  gate3111(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate3112(.a(s_366), .O(gate131inter3));
  inv1  gate3113(.a(s_367), .O(gate131inter4));
  nand2 gate3114(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate3115(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate3116(.a(G414), .O(gate131inter7));
  inv1  gate3117(.a(G415), .O(gate131inter8));
  nand2 gate3118(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate3119(.a(s_367), .b(gate131inter3), .O(gate131inter10));
  nor2  gate3120(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate3121(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate3122(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1233(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1234(.a(gate132inter0), .b(s_98), .O(gate132inter1));
  and2  gate1235(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1236(.a(s_98), .O(gate132inter3));
  inv1  gate1237(.a(s_99), .O(gate132inter4));
  nand2 gate1238(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1239(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1240(.a(G416), .O(gate132inter7));
  inv1  gate1241(.a(G417), .O(gate132inter8));
  nand2 gate1242(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1243(.a(s_99), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1244(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1245(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1246(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2199(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2200(.a(gate135inter0), .b(s_236), .O(gate135inter1));
  and2  gate2201(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2202(.a(s_236), .O(gate135inter3));
  inv1  gate2203(.a(s_237), .O(gate135inter4));
  nand2 gate2204(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2205(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2206(.a(G422), .O(gate135inter7));
  inv1  gate2207(.a(G423), .O(gate135inter8));
  nand2 gate2208(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2209(.a(s_237), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2210(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2211(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2212(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate2311(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2312(.a(gate136inter0), .b(s_252), .O(gate136inter1));
  and2  gate2313(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2314(.a(s_252), .O(gate136inter3));
  inv1  gate2315(.a(s_253), .O(gate136inter4));
  nand2 gate2316(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2317(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2318(.a(G424), .O(gate136inter7));
  inv1  gate2319(.a(G425), .O(gate136inter8));
  nand2 gate2320(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2321(.a(s_253), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2322(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2323(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2324(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate785(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate786(.a(gate137inter0), .b(s_34), .O(gate137inter1));
  and2  gate787(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate788(.a(s_34), .O(gate137inter3));
  inv1  gate789(.a(s_35), .O(gate137inter4));
  nand2 gate790(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate791(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate792(.a(G426), .O(gate137inter7));
  inv1  gate793(.a(G429), .O(gate137inter8));
  nand2 gate794(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate795(.a(s_35), .b(gate137inter3), .O(gate137inter10));
  nor2  gate796(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate797(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate798(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1681(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1682(.a(gate139inter0), .b(s_162), .O(gate139inter1));
  and2  gate1683(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1684(.a(s_162), .O(gate139inter3));
  inv1  gate1685(.a(s_163), .O(gate139inter4));
  nand2 gate1686(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1687(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1688(.a(G438), .O(gate139inter7));
  inv1  gate1689(.a(G441), .O(gate139inter8));
  nand2 gate1690(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1691(.a(s_163), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1692(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1693(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1694(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1471(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1472(.a(gate143inter0), .b(s_132), .O(gate143inter1));
  and2  gate1473(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1474(.a(s_132), .O(gate143inter3));
  inv1  gate1475(.a(s_133), .O(gate143inter4));
  nand2 gate1476(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1477(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1478(.a(G462), .O(gate143inter7));
  inv1  gate1479(.a(G465), .O(gate143inter8));
  nand2 gate1480(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1481(.a(s_133), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1482(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1483(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1484(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1261(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1262(.a(gate145inter0), .b(s_102), .O(gate145inter1));
  and2  gate1263(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1264(.a(s_102), .O(gate145inter3));
  inv1  gate1265(.a(s_103), .O(gate145inter4));
  nand2 gate1266(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1267(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1268(.a(G474), .O(gate145inter7));
  inv1  gate1269(.a(G477), .O(gate145inter8));
  nand2 gate1270(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1271(.a(s_103), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1272(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1273(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1274(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2339(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2340(.a(gate149inter0), .b(s_256), .O(gate149inter1));
  and2  gate2341(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2342(.a(s_256), .O(gate149inter3));
  inv1  gate2343(.a(s_257), .O(gate149inter4));
  nand2 gate2344(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2345(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2346(.a(G498), .O(gate149inter7));
  inv1  gate2347(.a(G501), .O(gate149inter8));
  nand2 gate2348(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2349(.a(s_257), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2350(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2351(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2352(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2325(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2326(.a(gate150inter0), .b(s_254), .O(gate150inter1));
  and2  gate2327(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2328(.a(s_254), .O(gate150inter3));
  inv1  gate2329(.a(s_255), .O(gate150inter4));
  nand2 gate2330(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2331(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2332(.a(G504), .O(gate150inter7));
  inv1  gate2333(.a(G507), .O(gate150inter8));
  nand2 gate2334(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2335(.a(s_255), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2336(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2337(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2338(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate603(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate604(.a(gate152inter0), .b(s_8), .O(gate152inter1));
  and2  gate605(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate606(.a(s_8), .O(gate152inter3));
  inv1  gate607(.a(s_9), .O(gate152inter4));
  nand2 gate608(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate609(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate610(.a(G516), .O(gate152inter7));
  inv1  gate611(.a(G519), .O(gate152inter8));
  nand2 gate612(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate613(.a(s_9), .b(gate152inter3), .O(gate152inter10));
  nor2  gate614(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate615(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate616(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate799(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate800(.a(gate153inter0), .b(s_36), .O(gate153inter1));
  and2  gate801(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate802(.a(s_36), .O(gate153inter3));
  inv1  gate803(.a(s_37), .O(gate153inter4));
  nand2 gate804(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate805(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate806(.a(G426), .O(gate153inter7));
  inv1  gate807(.a(G522), .O(gate153inter8));
  nand2 gate808(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate809(.a(s_37), .b(gate153inter3), .O(gate153inter10));
  nor2  gate810(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate811(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate812(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2171(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2172(.a(gate157inter0), .b(s_232), .O(gate157inter1));
  and2  gate2173(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2174(.a(s_232), .O(gate157inter3));
  inv1  gate2175(.a(s_233), .O(gate157inter4));
  nand2 gate2176(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2177(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2178(.a(G438), .O(gate157inter7));
  inv1  gate2179(.a(G528), .O(gate157inter8));
  nand2 gate2180(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2181(.a(s_233), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2182(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2183(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2184(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1513(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1514(.a(gate159inter0), .b(s_138), .O(gate159inter1));
  and2  gate1515(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1516(.a(s_138), .O(gate159inter3));
  inv1  gate1517(.a(s_139), .O(gate159inter4));
  nand2 gate1518(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1519(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1520(.a(G444), .O(gate159inter7));
  inv1  gate1521(.a(G531), .O(gate159inter8));
  nand2 gate1522(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1523(.a(s_139), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1524(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1525(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1526(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1863(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1864(.a(gate160inter0), .b(s_188), .O(gate160inter1));
  and2  gate1865(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1866(.a(s_188), .O(gate160inter3));
  inv1  gate1867(.a(s_189), .O(gate160inter4));
  nand2 gate1868(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1869(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1870(.a(G447), .O(gate160inter7));
  inv1  gate1871(.a(G531), .O(gate160inter8));
  nand2 gate1872(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1873(.a(s_189), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1874(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1875(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1876(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1163(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1164(.a(gate161inter0), .b(s_88), .O(gate161inter1));
  and2  gate1165(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1166(.a(s_88), .O(gate161inter3));
  inv1  gate1167(.a(s_89), .O(gate161inter4));
  nand2 gate1168(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1169(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1170(.a(G450), .O(gate161inter7));
  inv1  gate1171(.a(G534), .O(gate161inter8));
  nand2 gate1172(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1173(.a(s_89), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1174(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1175(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1176(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1905(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1906(.a(gate162inter0), .b(s_194), .O(gate162inter1));
  and2  gate1907(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1908(.a(s_194), .O(gate162inter3));
  inv1  gate1909(.a(s_195), .O(gate162inter4));
  nand2 gate1910(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1911(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1912(.a(G453), .O(gate162inter7));
  inv1  gate1913(.a(G534), .O(gate162inter8));
  nand2 gate1914(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1915(.a(s_195), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1916(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1917(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1918(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2521(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2522(.a(gate170inter0), .b(s_282), .O(gate170inter1));
  and2  gate2523(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2524(.a(s_282), .O(gate170inter3));
  inv1  gate2525(.a(s_283), .O(gate170inter4));
  nand2 gate2526(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2527(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2528(.a(G477), .O(gate170inter7));
  inv1  gate2529(.a(G546), .O(gate170inter8));
  nand2 gate2530(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2531(.a(s_283), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2532(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2533(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2534(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate3193(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate3194(.a(gate171inter0), .b(s_378), .O(gate171inter1));
  and2  gate3195(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate3196(.a(s_378), .O(gate171inter3));
  inv1  gate3197(.a(s_379), .O(gate171inter4));
  nand2 gate3198(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate3199(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate3200(.a(G480), .O(gate171inter7));
  inv1  gate3201(.a(G549), .O(gate171inter8));
  nand2 gate3202(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate3203(.a(s_379), .b(gate171inter3), .O(gate171inter10));
  nor2  gate3204(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate3205(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate3206(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate3165(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate3166(.a(gate172inter0), .b(s_374), .O(gate172inter1));
  and2  gate3167(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate3168(.a(s_374), .O(gate172inter3));
  inv1  gate3169(.a(s_375), .O(gate172inter4));
  nand2 gate3170(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate3171(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate3172(.a(G483), .O(gate172inter7));
  inv1  gate3173(.a(G549), .O(gate172inter8));
  nand2 gate3174(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate3175(.a(s_375), .b(gate172inter3), .O(gate172inter10));
  nor2  gate3176(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate3177(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate3178(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2115(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2116(.a(gate173inter0), .b(s_224), .O(gate173inter1));
  and2  gate2117(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2118(.a(s_224), .O(gate173inter3));
  inv1  gate2119(.a(s_225), .O(gate173inter4));
  nand2 gate2120(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2121(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2122(.a(G486), .O(gate173inter7));
  inv1  gate2123(.a(G552), .O(gate173inter8));
  nand2 gate2124(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2125(.a(s_225), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2126(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2127(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2128(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2143(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2144(.a(gate176inter0), .b(s_228), .O(gate176inter1));
  and2  gate2145(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2146(.a(s_228), .O(gate176inter3));
  inv1  gate2147(.a(s_229), .O(gate176inter4));
  nand2 gate2148(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2149(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2150(.a(G495), .O(gate176inter7));
  inv1  gate2151(.a(G555), .O(gate176inter8));
  nand2 gate2152(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2153(.a(s_229), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2154(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2155(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2156(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1107(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1108(.a(gate178inter0), .b(s_80), .O(gate178inter1));
  and2  gate1109(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1110(.a(s_80), .O(gate178inter3));
  inv1  gate1111(.a(s_81), .O(gate178inter4));
  nand2 gate1112(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1113(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1114(.a(G501), .O(gate178inter7));
  inv1  gate1115(.a(G558), .O(gate178inter8));
  nand2 gate1116(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1117(.a(s_81), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1118(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1119(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1120(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2759(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2760(.a(gate181inter0), .b(s_316), .O(gate181inter1));
  and2  gate2761(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2762(.a(s_316), .O(gate181inter3));
  inv1  gate2763(.a(s_317), .O(gate181inter4));
  nand2 gate2764(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2765(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2766(.a(G510), .O(gate181inter7));
  inv1  gate2767(.a(G564), .O(gate181inter8));
  nand2 gate2768(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2769(.a(s_317), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2770(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2771(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2772(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate3123(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate3124(.a(gate182inter0), .b(s_368), .O(gate182inter1));
  and2  gate3125(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate3126(.a(s_368), .O(gate182inter3));
  inv1  gate3127(.a(s_369), .O(gate182inter4));
  nand2 gate3128(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate3129(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate3130(.a(G513), .O(gate182inter7));
  inv1  gate3131(.a(G564), .O(gate182inter8));
  nand2 gate3132(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate3133(.a(s_369), .b(gate182inter3), .O(gate182inter10));
  nor2  gate3134(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate3135(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate3136(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1485(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1486(.a(gate183inter0), .b(s_134), .O(gate183inter1));
  and2  gate1487(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1488(.a(s_134), .O(gate183inter3));
  inv1  gate1489(.a(s_135), .O(gate183inter4));
  nand2 gate1490(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1491(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1492(.a(G516), .O(gate183inter7));
  inv1  gate1493(.a(G567), .O(gate183inter8));
  nand2 gate1494(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1495(.a(s_135), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1496(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1497(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1498(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate2017(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2018(.a(gate184inter0), .b(s_210), .O(gate184inter1));
  and2  gate2019(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2020(.a(s_210), .O(gate184inter3));
  inv1  gate2021(.a(s_211), .O(gate184inter4));
  nand2 gate2022(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2023(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2024(.a(G519), .O(gate184inter7));
  inv1  gate2025(.a(G567), .O(gate184inter8));
  nand2 gate2026(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2027(.a(s_211), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2028(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2029(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2030(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2899(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2900(.a(gate185inter0), .b(s_336), .O(gate185inter1));
  and2  gate2901(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2902(.a(s_336), .O(gate185inter3));
  inv1  gate2903(.a(s_337), .O(gate185inter4));
  nand2 gate2904(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2905(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2906(.a(G570), .O(gate185inter7));
  inv1  gate2907(.a(G571), .O(gate185inter8));
  nand2 gate2908(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2909(.a(s_337), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2910(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2911(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2912(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1975(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1976(.a(gate186inter0), .b(s_204), .O(gate186inter1));
  and2  gate1977(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1978(.a(s_204), .O(gate186inter3));
  inv1  gate1979(.a(s_205), .O(gate186inter4));
  nand2 gate1980(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1981(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1982(.a(G572), .O(gate186inter7));
  inv1  gate1983(.a(G573), .O(gate186inter8));
  nand2 gate1984(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1985(.a(s_205), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1986(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1987(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1988(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2185(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2186(.a(gate189inter0), .b(s_234), .O(gate189inter1));
  and2  gate2187(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2188(.a(s_234), .O(gate189inter3));
  inv1  gate2189(.a(s_235), .O(gate189inter4));
  nand2 gate2190(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2191(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2192(.a(G578), .O(gate189inter7));
  inv1  gate2193(.a(G579), .O(gate189inter8));
  nand2 gate2194(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2195(.a(s_235), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2196(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2197(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2198(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1961(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1962(.a(gate192inter0), .b(s_202), .O(gate192inter1));
  and2  gate1963(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1964(.a(s_202), .O(gate192inter3));
  inv1  gate1965(.a(s_203), .O(gate192inter4));
  nand2 gate1966(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1967(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1968(.a(G584), .O(gate192inter7));
  inv1  gate1969(.a(G585), .O(gate192inter8));
  nand2 gate1970(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1971(.a(s_203), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1972(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1973(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1974(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate547(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate548(.a(gate194inter0), .b(s_0), .O(gate194inter1));
  and2  gate549(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate550(.a(s_0), .O(gate194inter3));
  inv1  gate551(.a(s_1), .O(gate194inter4));
  nand2 gate552(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate553(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate554(.a(G588), .O(gate194inter7));
  inv1  gate555(.a(G589), .O(gate194inter8));
  nand2 gate556(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate557(.a(s_1), .b(gate194inter3), .O(gate194inter10));
  nor2  gate558(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate559(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate560(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2871(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2872(.a(gate197inter0), .b(s_332), .O(gate197inter1));
  and2  gate2873(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2874(.a(s_332), .O(gate197inter3));
  inv1  gate2875(.a(s_333), .O(gate197inter4));
  nand2 gate2876(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2877(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2878(.a(G594), .O(gate197inter7));
  inv1  gate2879(.a(G595), .O(gate197inter8));
  nand2 gate2880(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2881(.a(s_333), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2882(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2883(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2884(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate2353(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2354(.a(gate198inter0), .b(s_258), .O(gate198inter1));
  and2  gate2355(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2356(.a(s_258), .O(gate198inter3));
  inv1  gate2357(.a(s_259), .O(gate198inter4));
  nand2 gate2358(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2359(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2360(.a(G596), .O(gate198inter7));
  inv1  gate2361(.a(G597), .O(gate198inter8));
  nand2 gate2362(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2363(.a(s_259), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2364(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2365(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2366(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2689(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2690(.a(gate200inter0), .b(s_306), .O(gate200inter1));
  and2  gate2691(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2692(.a(s_306), .O(gate200inter3));
  inv1  gate2693(.a(s_307), .O(gate200inter4));
  nand2 gate2694(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2695(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2696(.a(G600), .O(gate200inter7));
  inv1  gate2697(.a(G601), .O(gate200inter8));
  nand2 gate2698(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2699(.a(s_307), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2700(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2701(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2702(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate2059(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2060(.a(gate201inter0), .b(s_216), .O(gate201inter1));
  and2  gate2061(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2062(.a(s_216), .O(gate201inter3));
  inv1  gate2063(.a(s_217), .O(gate201inter4));
  nand2 gate2064(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2065(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2066(.a(G602), .O(gate201inter7));
  inv1  gate2067(.a(G607), .O(gate201inter8));
  nand2 gate2068(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2069(.a(s_217), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2070(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2071(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2072(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2255(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2256(.a(gate204inter0), .b(s_244), .O(gate204inter1));
  and2  gate2257(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2258(.a(s_244), .O(gate204inter3));
  inv1  gate2259(.a(s_245), .O(gate204inter4));
  nand2 gate2260(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2261(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2262(.a(G607), .O(gate204inter7));
  inv1  gate2263(.a(G617), .O(gate204inter8));
  nand2 gate2264(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2265(.a(s_245), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2266(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2267(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2268(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1583(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1584(.a(gate209inter0), .b(s_148), .O(gate209inter1));
  and2  gate1585(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1586(.a(s_148), .O(gate209inter3));
  inv1  gate1587(.a(s_149), .O(gate209inter4));
  nand2 gate1588(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1589(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1590(.a(G602), .O(gate209inter7));
  inv1  gate1591(.a(G666), .O(gate209inter8));
  nand2 gate1592(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1593(.a(s_149), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1594(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1595(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1596(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2297(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2298(.a(gate213inter0), .b(s_250), .O(gate213inter1));
  and2  gate2299(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2300(.a(s_250), .O(gate213inter3));
  inv1  gate2301(.a(s_251), .O(gate213inter4));
  nand2 gate2302(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2303(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2304(.a(G602), .O(gate213inter7));
  inv1  gate2305(.a(G672), .O(gate213inter8));
  nand2 gate2306(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2307(.a(s_251), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2308(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2309(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2310(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1359(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1360(.a(gate219inter0), .b(s_116), .O(gate219inter1));
  and2  gate1361(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1362(.a(s_116), .O(gate219inter3));
  inv1  gate1363(.a(s_117), .O(gate219inter4));
  nand2 gate1364(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1365(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1366(.a(G632), .O(gate219inter7));
  inv1  gate1367(.a(G681), .O(gate219inter8));
  nand2 gate1368(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1369(.a(s_117), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1370(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1371(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1372(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate883(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate884(.a(gate221inter0), .b(s_48), .O(gate221inter1));
  and2  gate885(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate886(.a(s_48), .O(gate221inter3));
  inv1  gate887(.a(s_49), .O(gate221inter4));
  nand2 gate888(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate889(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate890(.a(G622), .O(gate221inter7));
  inv1  gate891(.a(G684), .O(gate221inter8));
  nand2 gate892(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate893(.a(s_49), .b(gate221inter3), .O(gate221inter10));
  nor2  gate894(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate895(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate896(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2003(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2004(.a(gate224inter0), .b(s_208), .O(gate224inter1));
  and2  gate2005(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2006(.a(s_208), .O(gate224inter3));
  inv1  gate2007(.a(s_209), .O(gate224inter4));
  nand2 gate2008(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2009(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2010(.a(G637), .O(gate224inter7));
  inv1  gate2011(.a(G687), .O(gate224inter8));
  nand2 gate2012(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2013(.a(s_209), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2014(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2015(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2016(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1415(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1416(.a(gate225inter0), .b(s_124), .O(gate225inter1));
  and2  gate1417(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1418(.a(s_124), .O(gate225inter3));
  inv1  gate1419(.a(s_125), .O(gate225inter4));
  nand2 gate1420(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1421(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1422(.a(G690), .O(gate225inter7));
  inv1  gate1423(.a(G691), .O(gate225inter8));
  nand2 gate1424(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1425(.a(s_125), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1426(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1427(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1428(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2493(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2494(.a(gate231inter0), .b(s_278), .O(gate231inter1));
  and2  gate2495(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2496(.a(s_278), .O(gate231inter3));
  inv1  gate2497(.a(s_279), .O(gate231inter4));
  nand2 gate2498(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2499(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2500(.a(G702), .O(gate231inter7));
  inv1  gate2501(.a(G703), .O(gate231inter8));
  nand2 gate2502(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2503(.a(s_279), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2504(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2505(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2506(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2717(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2718(.a(gate232inter0), .b(s_310), .O(gate232inter1));
  and2  gate2719(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2720(.a(s_310), .O(gate232inter3));
  inv1  gate2721(.a(s_311), .O(gate232inter4));
  nand2 gate2722(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2723(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2724(.a(G704), .O(gate232inter7));
  inv1  gate2725(.a(G705), .O(gate232inter8));
  nand2 gate2726(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2727(.a(s_311), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2728(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2729(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2730(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate897(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate898(.a(gate233inter0), .b(s_50), .O(gate233inter1));
  and2  gate899(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate900(.a(s_50), .O(gate233inter3));
  inv1  gate901(.a(s_51), .O(gate233inter4));
  nand2 gate902(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate903(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate904(.a(G242), .O(gate233inter7));
  inv1  gate905(.a(G718), .O(gate233inter8));
  nand2 gate906(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate907(.a(s_51), .b(gate233inter3), .O(gate233inter10));
  nor2  gate908(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate909(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate910(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1849(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1850(.a(gate234inter0), .b(s_186), .O(gate234inter1));
  and2  gate1851(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1852(.a(s_186), .O(gate234inter3));
  inv1  gate1853(.a(s_187), .O(gate234inter4));
  nand2 gate1854(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1855(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1856(.a(G245), .O(gate234inter7));
  inv1  gate1857(.a(G721), .O(gate234inter8));
  nand2 gate1858(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1859(.a(s_187), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1860(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1861(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1862(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1667(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1668(.a(gate236inter0), .b(s_160), .O(gate236inter1));
  and2  gate1669(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1670(.a(s_160), .O(gate236inter3));
  inv1  gate1671(.a(s_161), .O(gate236inter4));
  nand2 gate1672(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1673(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1674(.a(G251), .O(gate236inter7));
  inv1  gate1675(.a(G727), .O(gate236inter8));
  nand2 gate1676(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1677(.a(s_161), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1678(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1679(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1680(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate2843(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2844(.a(gate238inter0), .b(s_328), .O(gate238inter1));
  and2  gate2845(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2846(.a(s_328), .O(gate238inter3));
  inv1  gate2847(.a(s_329), .O(gate238inter4));
  nand2 gate2848(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2849(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2850(.a(G257), .O(gate238inter7));
  inv1  gate2851(.a(G709), .O(gate238inter8));
  nand2 gate2852(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2853(.a(s_329), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2854(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2855(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2856(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate3011(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate3012(.a(gate239inter0), .b(s_352), .O(gate239inter1));
  and2  gate3013(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate3014(.a(s_352), .O(gate239inter3));
  inv1  gate3015(.a(s_353), .O(gate239inter4));
  nand2 gate3016(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate3017(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate3018(.a(G260), .O(gate239inter7));
  inv1  gate3019(.a(G712), .O(gate239inter8));
  nand2 gate3020(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate3021(.a(s_353), .b(gate239inter3), .O(gate239inter10));
  nor2  gate3022(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate3023(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate3024(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2927(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2928(.a(gate241inter0), .b(s_340), .O(gate241inter1));
  and2  gate2929(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2930(.a(s_340), .O(gate241inter3));
  inv1  gate2931(.a(s_341), .O(gate241inter4));
  nand2 gate2932(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2933(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2934(.a(G242), .O(gate241inter7));
  inv1  gate2935(.a(G730), .O(gate241inter8));
  nand2 gate2936(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2937(.a(s_341), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2938(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2939(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2940(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate2731(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2732(.a(gate242inter0), .b(s_312), .O(gate242inter1));
  and2  gate2733(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2734(.a(s_312), .O(gate242inter3));
  inv1  gate2735(.a(s_313), .O(gate242inter4));
  nand2 gate2736(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2737(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2738(.a(G718), .O(gate242inter7));
  inv1  gate2739(.a(G730), .O(gate242inter8));
  nand2 gate2740(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2741(.a(s_313), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2742(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2743(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2744(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate2983(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2984(.a(gate243inter0), .b(s_348), .O(gate243inter1));
  and2  gate2985(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2986(.a(s_348), .O(gate243inter3));
  inv1  gate2987(.a(s_349), .O(gate243inter4));
  nand2 gate2988(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2989(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2990(.a(G245), .O(gate243inter7));
  inv1  gate2991(.a(G733), .O(gate243inter8));
  nand2 gate2992(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2993(.a(s_349), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2994(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2995(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2996(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2773(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2774(.a(gate246inter0), .b(s_318), .O(gate246inter1));
  and2  gate2775(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2776(.a(s_318), .O(gate246inter3));
  inv1  gate2777(.a(s_319), .O(gate246inter4));
  nand2 gate2778(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2779(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2780(.a(G724), .O(gate246inter7));
  inv1  gate2781(.a(G736), .O(gate246inter8));
  nand2 gate2782(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2783(.a(s_319), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2784(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2785(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2786(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1443(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1444(.a(gate248inter0), .b(s_128), .O(gate248inter1));
  and2  gate1445(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1446(.a(s_128), .O(gate248inter3));
  inv1  gate1447(.a(s_129), .O(gate248inter4));
  nand2 gate1448(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1449(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1450(.a(G727), .O(gate248inter7));
  inv1  gate1451(.a(G739), .O(gate248inter8));
  nand2 gate1452(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1453(.a(s_129), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1454(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1455(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1456(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate925(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate926(.a(gate250inter0), .b(s_54), .O(gate250inter1));
  and2  gate927(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate928(.a(s_54), .O(gate250inter3));
  inv1  gate929(.a(s_55), .O(gate250inter4));
  nand2 gate930(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate931(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate932(.a(G706), .O(gate250inter7));
  inv1  gate933(.a(G742), .O(gate250inter8));
  nand2 gate934(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate935(.a(s_55), .b(gate250inter3), .O(gate250inter10));
  nor2  gate936(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate937(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate938(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2703(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2704(.a(gate251inter0), .b(s_308), .O(gate251inter1));
  and2  gate2705(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2706(.a(s_308), .O(gate251inter3));
  inv1  gate2707(.a(s_309), .O(gate251inter4));
  nand2 gate2708(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2709(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2710(.a(G257), .O(gate251inter7));
  inv1  gate2711(.a(G745), .O(gate251inter8));
  nand2 gate2712(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2713(.a(s_309), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2714(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2715(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2716(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate589(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate590(.a(gate252inter0), .b(s_6), .O(gate252inter1));
  and2  gate591(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate592(.a(s_6), .O(gate252inter3));
  inv1  gate593(.a(s_7), .O(gate252inter4));
  nand2 gate594(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate595(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate596(.a(G709), .O(gate252inter7));
  inv1  gate597(.a(G745), .O(gate252inter8));
  nand2 gate598(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate599(.a(s_7), .b(gate252inter3), .O(gate252inter10));
  nor2  gate600(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate601(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate602(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate3137(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate3138(.a(gate253inter0), .b(s_370), .O(gate253inter1));
  and2  gate3139(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate3140(.a(s_370), .O(gate253inter3));
  inv1  gate3141(.a(s_371), .O(gate253inter4));
  nand2 gate3142(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate3143(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate3144(.a(G260), .O(gate253inter7));
  inv1  gate3145(.a(G748), .O(gate253inter8));
  nand2 gate3146(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate3147(.a(s_371), .b(gate253inter3), .O(gate253inter10));
  nor2  gate3148(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate3149(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate3150(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2479(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2480(.a(gate255inter0), .b(s_276), .O(gate255inter1));
  and2  gate2481(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2482(.a(s_276), .O(gate255inter3));
  inv1  gate2483(.a(s_277), .O(gate255inter4));
  nand2 gate2484(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2485(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2486(.a(G263), .O(gate255inter7));
  inv1  gate2487(.a(G751), .O(gate255inter8));
  nand2 gate2488(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2489(.a(s_277), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2490(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2491(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2492(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2283(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2284(.a(gate257inter0), .b(s_248), .O(gate257inter1));
  and2  gate2285(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2286(.a(s_248), .O(gate257inter3));
  inv1  gate2287(.a(s_249), .O(gate257inter4));
  nand2 gate2288(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2289(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2290(.a(G754), .O(gate257inter7));
  inv1  gate2291(.a(G755), .O(gate257inter8));
  nand2 gate2292(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2293(.a(s_249), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2294(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2295(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2296(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate2619(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2620(.a(gate259inter0), .b(s_296), .O(gate259inter1));
  and2  gate2621(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2622(.a(s_296), .O(gate259inter3));
  inv1  gate2623(.a(s_297), .O(gate259inter4));
  nand2 gate2624(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2625(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2626(.a(G758), .O(gate259inter7));
  inv1  gate2627(.a(G759), .O(gate259inter8));
  nand2 gate2628(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2629(.a(s_297), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2630(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2631(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2632(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1723(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1724(.a(gate260inter0), .b(s_168), .O(gate260inter1));
  and2  gate1725(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1726(.a(s_168), .O(gate260inter3));
  inv1  gate1727(.a(s_169), .O(gate260inter4));
  nand2 gate1728(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1729(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1730(.a(G760), .O(gate260inter7));
  inv1  gate1731(.a(G761), .O(gate260inter8));
  nand2 gate1732(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1733(.a(s_169), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1734(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1735(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1736(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate2395(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2396(.a(gate266inter0), .b(s_264), .O(gate266inter1));
  and2  gate2397(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2398(.a(s_264), .O(gate266inter3));
  inv1  gate2399(.a(s_265), .O(gate266inter4));
  nand2 gate2400(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2401(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2402(.a(G645), .O(gate266inter7));
  inv1  gate2403(.a(G773), .O(gate266inter8));
  nand2 gate2404(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2405(.a(s_265), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2406(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2407(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2408(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1317(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1318(.a(gate269inter0), .b(s_110), .O(gate269inter1));
  and2  gate1319(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1320(.a(s_110), .O(gate269inter3));
  inv1  gate1321(.a(s_111), .O(gate269inter4));
  nand2 gate1322(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1323(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1324(.a(G654), .O(gate269inter7));
  inv1  gate1325(.a(G782), .O(gate269inter8));
  nand2 gate1326(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1327(.a(s_111), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1328(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1329(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1330(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate3067(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate3068(.a(gate270inter0), .b(s_360), .O(gate270inter1));
  and2  gate3069(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate3070(.a(s_360), .O(gate270inter3));
  inv1  gate3071(.a(s_361), .O(gate270inter4));
  nand2 gate3072(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate3073(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate3074(.a(G657), .O(gate270inter7));
  inv1  gate3075(.a(G785), .O(gate270inter8));
  nand2 gate3076(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate3077(.a(s_361), .b(gate270inter3), .O(gate270inter10));
  nor2  gate3078(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate3079(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate3080(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate715(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate716(.a(gate272inter0), .b(s_24), .O(gate272inter1));
  and2  gate717(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate718(.a(s_24), .O(gate272inter3));
  inv1  gate719(.a(s_25), .O(gate272inter4));
  nand2 gate720(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate721(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate722(.a(G663), .O(gate272inter7));
  inv1  gate723(.a(G791), .O(gate272inter8));
  nand2 gate724(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate725(.a(s_25), .b(gate272inter3), .O(gate272inter10));
  nor2  gate726(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate727(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate728(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate2087(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2088(.a(gate273inter0), .b(s_220), .O(gate273inter1));
  and2  gate2089(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2090(.a(s_220), .O(gate273inter3));
  inv1  gate2091(.a(s_221), .O(gate273inter4));
  nand2 gate2092(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2093(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2094(.a(G642), .O(gate273inter7));
  inv1  gate2095(.a(G794), .O(gate273inter8));
  nand2 gate2096(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2097(.a(s_221), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2098(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2099(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2100(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate855(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate856(.a(gate277inter0), .b(s_44), .O(gate277inter1));
  and2  gate857(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate858(.a(s_44), .O(gate277inter3));
  inv1  gate859(.a(s_45), .O(gate277inter4));
  nand2 gate860(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate861(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate862(.a(G648), .O(gate277inter7));
  inv1  gate863(.a(G800), .O(gate277inter8));
  nand2 gate864(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate865(.a(s_45), .b(gate277inter3), .O(gate277inter10));
  nor2  gate866(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate867(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate868(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate2507(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2508(.a(gate278inter0), .b(s_280), .O(gate278inter1));
  and2  gate2509(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2510(.a(s_280), .O(gate278inter3));
  inv1  gate2511(.a(s_281), .O(gate278inter4));
  nand2 gate2512(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2513(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2514(.a(G776), .O(gate278inter7));
  inv1  gate2515(.a(G800), .O(gate278inter8));
  nand2 gate2516(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2517(.a(s_281), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2518(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2519(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2520(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1373(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1374(.a(gate281inter0), .b(s_118), .O(gate281inter1));
  and2  gate1375(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1376(.a(s_118), .O(gate281inter3));
  inv1  gate1377(.a(s_119), .O(gate281inter4));
  nand2 gate1378(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1379(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1380(.a(G654), .O(gate281inter7));
  inv1  gate1381(.a(G806), .O(gate281inter8));
  nand2 gate1382(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1383(.a(s_119), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1384(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1385(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1386(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2829(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2830(.a(gate282inter0), .b(s_326), .O(gate282inter1));
  and2  gate2831(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2832(.a(s_326), .O(gate282inter3));
  inv1  gate2833(.a(s_327), .O(gate282inter4));
  nand2 gate2834(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2835(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2836(.a(G782), .O(gate282inter7));
  inv1  gate2837(.a(G806), .O(gate282inter8));
  nand2 gate2838(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2839(.a(s_327), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2840(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2841(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2842(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1611(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1612(.a(gate283inter0), .b(s_152), .O(gate283inter1));
  and2  gate1613(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1614(.a(s_152), .O(gate283inter3));
  inv1  gate1615(.a(s_153), .O(gate283inter4));
  nand2 gate1616(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1617(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1618(.a(G657), .O(gate283inter7));
  inv1  gate1619(.a(G809), .O(gate283inter8));
  nand2 gate1620(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1621(.a(s_153), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1622(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1623(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1624(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1877(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1878(.a(gate284inter0), .b(s_190), .O(gate284inter1));
  and2  gate1879(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1880(.a(s_190), .O(gate284inter3));
  inv1  gate1881(.a(s_191), .O(gate284inter4));
  nand2 gate1882(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1883(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1884(.a(G785), .O(gate284inter7));
  inv1  gate1885(.a(G809), .O(gate284inter8));
  nand2 gate1886(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1887(.a(s_191), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1888(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1889(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1890(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2031(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2032(.a(gate286inter0), .b(s_212), .O(gate286inter1));
  and2  gate2033(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2034(.a(s_212), .O(gate286inter3));
  inv1  gate2035(.a(s_213), .O(gate286inter4));
  nand2 gate2036(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2037(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2038(.a(G788), .O(gate286inter7));
  inv1  gate2039(.a(G812), .O(gate286inter8));
  nand2 gate2040(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2041(.a(s_213), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2042(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2043(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2044(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1821(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1822(.a(gate287inter0), .b(s_182), .O(gate287inter1));
  and2  gate1823(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1824(.a(s_182), .O(gate287inter3));
  inv1  gate1825(.a(s_183), .O(gate287inter4));
  nand2 gate1826(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1827(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1828(.a(G663), .O(gate287inter7));
  inv1  gate1829(.a(G815), .O(gate287inter8));
  nand2 gate1830(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1831(.a(s_183), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1832(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1833(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1834(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate3053(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate3054(.a(gate288inter0), .b(s_358), .O(gate288inter1));
  and2  gate3055(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate3056(.a(s_358), .O(gate288inter3));
  inv1  gate3057(.a(s_359), .O(gate288inter4));
  nand2 gate3058(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate3059(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate3060(.a(G791), .O(gate288inter7));
  inv1  gate3061(.a(G815), .O(gate288inter8));
  nand2 gate3062(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate3063(.a(s_359), .b(gate288inter3), .O(gate288inter10));
  nor2  gate3064(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate3065(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate3066(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1793(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1794(.a(gate293inter0), .b(s_178), .O(gate293inter1));
  and2  gate1795(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1796(.a(s_178), .O(gate293inter3));
  inv1  gate1797(.a(s_179), .O(gate293inter4));
  nand2 gate1798(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1799(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1800(.a(G828), .O(gate293inter7));
  inv1  gate1801(.a(G829), .O(gate293inter8));
  nand2 gate1802(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1803(.a(s_179), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1804(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1805(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1806(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate3039(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate3040(.a(gate294inter0), .b(s_356), .O(gate294inter1));
  and2  gate3041(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate3042(.a(s_356), .O(gate294inter3));
  inv1  gate3043(.a(s_357), .O(gate294inter4));
  nand2 gate3044(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate3045(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate3046(.a(G832), .O(gate294inter7));
  inv1  gate3047(.a(G833), .O(gate294inter8));
  nand2 gate3048(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate3049(.a(s_357), .b(gate294inter3), .O(gate294inter10));
  nor2  gate3050(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate3051(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate3052(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate757(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate758(.a(gate388inter0), .b(s_30), .O(gate388inter1));
  and2  gate759(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate760(.a(s_30), .O(gate388inter3));
  inv1  gate761(.a(s_31), .O(gate388inter4));
  nand2 gate762(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate763(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate764(.a(G2), .O(gate388inter7));
  inv1  gate765(.a(G1039), .O(gate388inter8));
  nand2 gate766(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate767(.a(s_31), .b(gate388inter3), .O(gate388inter10));
  nor2  gate768(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate769(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate770(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2423(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2424(.a(gate389inter0), .b(s_268), .O(gate389inter1));
  and2  gate2425(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2426(.a(s_268), .O(gate389inter3));
  inv1  gate2427(.a(s_269), .O(gate389inter4));
  nand2 gate2428(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2429(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2430(.a(G3), .O(gate389inter7));
  inv1  gate2431(.a(G1042), .O(gate389inter8));
  nand2 gate2432(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2433(.a(s_269), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2434(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2435(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2436(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1989(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1990(.a(gate392inter0), .b(s_206), .O(gate392inter1));
  and2  gate1991(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1992(.a(s_206), .O(gate392inter3));
  inv1  gate1993(.a(s_207), .O(gate392inter4));
  nand2 gate1994(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1995(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1996(.a(G6), .O(gate392inter7));
  inv1  gate1997(.a(G1051), .O(gate392inter8));
  nand2 gate1998(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1999(.a(s_207), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2000(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2001(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2002(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1135(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1136(.a(gate395inter0), .b(s_84), .O(gate395inter1));
  and2  gate1137(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1138(.a(s_84), .O(gate395inter3));
  inv1  gate1139(.a(s_85), .O(gate395inter4));
  nand2 gate1140(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1141(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1142(.a(G9), .O(gate395inter7));
  inv1  gate1143(.a(G1060), .O(gate395inter8));
  nand2 gate1144(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1145(.a(s_85), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1146(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1147(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1148(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1499(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1500(.a(gate396inter0), .b(s_136), .O(gate396inter1));
  and2  gate1501(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1502(.a(s_136), .O(gate396inter3));
  inv1  gate1503(.a(s_137), .O(gate396inter4));
  nand2 gate1504(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1505(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1506(.a(G10), .O(gate396inter7));
  inv1  gate1507(.a(G1063), .O(gate396inter8));
  nand2 gate1508(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1509(.a(s_137), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1510(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1511(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1512(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1275(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1276(.a(gate397inter0), .b(s_104), .O(gate397inter1));
  and2  gate1277(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1278(.a(s_104), .O(gate397inter3));
  inv1  gate1279(.a(s_105), .O(gate397inter4));
  nand2 gate1280(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1281(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1282(.a(G11), .O(gate397inter7));
  inv1  gate1283(.a(G1066), .O(gate397inter8));
  nand2 gate1284(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1285(.a(s_105), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1286(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1287(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1288(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1457(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1458(.a(gate402inter0), .b(s_130), .O(gate402inter1));
  and2  gate1459(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1460(.a(s_130), .O(gate402inter3));
  inv1  gate1461(.a(s_131), .O(gate402inter4));
  nand2 gate1462(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1463(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1464(.a(G16), .O(gate402inter7));
  inv1  gate1465(.a(G1081), .O(gate402inter8));
  nand2 gate1466(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1467(.a(s_131), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1468(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1469(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1470(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1205(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1206(.a(gate403inter0), .b(s_94), .O(gate403inter1));
  and2  gate1207(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1208(.a(s_94), .O(gate403inter3));
  inv1  gate1209(.a(s_95), .O(gate403inter4));
  nand2 gate1210(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1211(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1212(.a(G17), .O(gate403inter7));
  inv1  gate1213(.a(G1084), .O(gate403inter8));
  nand2 gate1214(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1215(.a(s_95), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1216(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1217(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1218(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2227(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2228(.a(gate407inter0), .b(s_240), .O(gate407inter1));
  and2  gate2229(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2230(.a(s_240), .O(gate407inter3));
  inv1  gate2231(.a(s_241), .O(gate407inter4));
  nand2 gate2232(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2233(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2234(.a(G21), .O(gate407inter7));
  inv1  gate2235(.a(G1096), .O(gate407inter8));
  nand2 gate2236(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2237(.a(s_241), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2238(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2239(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2240(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate911(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate912(.a(gate408inter0), .b(s_52), .O(gate408inter1));
  and2  gate913(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate914(.a(s_52), .O(gate408inter3));
  inv1  gate915(.a(s_53), .O(gate408inter4));
  nand2 gate916(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate917(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate918(.a(G22), .O(gate408inter7));
  inv1  gate919(.a(G1099), .O(gate408inter8));
  nand2 gate920(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate921(.a(s_53), .b(gate408inter3), .O(gate408inter10));
  nor2  gate922(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate923(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate924(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1247(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1248(.a(gate412inter0), .b(s_100), .O(gate412inter1));
  and2  gate1249(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1250(.a(s_100), .O(gate412inter3));
  inv1  gate1251(.a(s_101), .O(gate412inter4));
  nand2 gate1252(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1253(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1254(.a(G26), .O(gate412inter7));
  inv1  gate1255(.a(G1111), .O(gate412inter8));
  nand2 gate1256(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1257(.a(s_101), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1258(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1259(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1260(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1933(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1934(.a(gate417inter0), .b(s_198), .O(gate417inter1));
  and2  gate1935(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1936(.a(s_198), .O(gate417inter3));
  inv1  gate1937(.a(s_199), .O(gate417inter4));
  nand2 gate1938(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1939(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1940(.a(G31), .O(gate417inter7));
  inv1  gate1941(.a(G1126), .O(gate417inter8));
  nand2 gate1942(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1943(.a(s_199), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1944(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1945(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1946(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2591(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2592(.a(gate423inter0), .b(s_292), .O(gate423inter1));
  and2  gate2593(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2594(.a(s_292), .O(gate423inter3));
  inv1  gate2595(.a(s_293), .O(gate423inter4));
  nand2 gate2596(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2597(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2598(.a(G3), .O(gate423inter7));
  inv1  gate2599(.a(G1138), .O(gate423inter8));
  nand2 gate2600(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2601(.a(s_293), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2602(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2603(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2604(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate687(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate688(.a(gate431inter0), .b(s_20), .O(gate431inter1));
  and2  gate689(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate690(.a(s_20), .O(gate431inter3));
  inv1  gate691(.a(s_21), .O(gate431inter4));
  nand2 gate692(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate693(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate694(.a(G7), .O(gate431inter7));
  inv1  gate695(.a(G1150), .O(gate431inter8));
  nand2 gate696(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate697(.a(s_21), .b(gate431inter3), .O(gate431inter10));
  nor2  gate698(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate699(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate700(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2045(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2046(.a(gate432inter0), .b(s_214), .O(gate432inter1));
  and2  gate2047(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2048(.a(s_214), .O(gate432inter3));
  inv1  gate2049(.a(s_215), .O(gate432inter4));
  nand2 gate2050(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2051(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2052(.a(G1054), .O(gate432inter7));
  inv1  gate2053(.a(G1150), .O(gate432inter8));
  nand2 gate2054(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2055(.a(s_215), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2056(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2057(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2058(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2633(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2634(.a(gate434inter0), .b(s_298), .O(gate434inter1));
  and2  gate2635(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2636(.a(s_298), .O(gate434inter3));
  inv1  gate2637(.a(s_299), .O(gate434inter4));
  nand2 gate2638(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2639(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2640(.a(G1057), .O(gate434inter7));
  inv1  gate2641(.a(G1153), .O(gate434inter8));
  nand2 gate2642(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2643(.a(s_299), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2644(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2645(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2646(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1751(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1752(.a(gate437inter0), .b(s_172), .O(gate437inter1));
  and2  gate1753(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1754(.a(s_172), .O(gate437inter3));
  inv1  gate1755(.a(s_173), .O(gate437inter4));
  nand2 gate1756(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1757(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1758(.a(G10), .O(gate437inter7));
  inv1  gate1759(.a(G1159), .O(gate437inter8));
  nand2 gate1760(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1761(.a(s_173), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1762(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1763(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1764(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1569(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1570(.a(gate438inter0), .b(s_146), .O(gate438inter1));
  and2  gate1571(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1572(.a(s_146), .O(gate438inter3));
  inv1  gate1573(.a(s_147), .O(gate438inter4));
  nand2 gate1574(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1575(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1576(.a(G1063), .O(gate438inter7));
  inv1  gate1577(.a(G1159), .O(gate438inter8));
  nand2 gate1578(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1579(.a(s_147), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1580(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1581(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1582(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2997(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2998(.a(gate440inter0), .b(s_350), .O(gate440inter1));
  and2  gate2999(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate3000(.a(s_350), .O(gate440inter3));
  inv1  gate3001(.a(s_351), .O(gate440inter4));
  nand2 gate3002(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate3003(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate3004(.a(G1066), .O(gate440inter7));
  inv1  gate3005(.a(G1162), .O(gate440inter8));
  nand2 gate3006(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate3007(.a(s_351), .b(gate440inter3), .O(gate440inter10));
  nor2  gate3008(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate3009(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate3010(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2073(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2074(.a(gate445inter0), .b(s_218), .O(gate445inter1));
  and2  gate2075(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2076(.a(s_218), .O(gate445inter3));
  inv1  gate2077(.a(s_219), .O(gate445inter4));
  nand2 gate2078(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2079(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2080(.a(G14), .O(gate445inter7));
  inv1  gate2081(.a(G1171), .O(gate445inter8));
  nand2 gate2082(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2083(.a(s_219), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2084(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2085(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2086(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate659(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate660(.a(gate446inter0), .b(s_16), .O(gate446inter1));
  and2  gate661(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate662(.a(s_16), .O(gate446inter3));
  inv1  gate663(.a(s_17), .O(gate446inter4));
  nand2 gate664(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate665(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate666(.a(G1075), .O(gate446inter7));
  inv1  gate667(.a(G1171), .O(gate446inter8));
  nand2 gate668(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate669(.a(s_17), .b(gate446inter3), .O(gate446inter10));
  nor2  gate670(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate671(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate672(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2465(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2466(.a(gate451inter0), .b(s_274), .O(gate451inter1));
  and2  gate2467(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2468(.a(s_274), .O(gate451inter3));
  inv1  gate2469(.a(s_275), .O(gate451inter4));
  nand2 gate2470(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2471(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2472(.a(G17), .O(gate451inter7));
  inv1  gate2473(.a(G1180), .O(gate451inter8));
  nand2 gate2474(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2475(.a(s_275), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2476(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2477(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2478(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate869(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate870(.a(gate454inter0), .b(s_46), .O(gate454inter1));
  and2  gate871(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate872(.a(s_46), .O(gate454inter3));
  inv1  gate873(.a(s_47), .O(gate454inter4));
  nand2 gate874(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate875(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate876(.a(G1087), .O(gate454inter7));
  inv1  gate877(.a(G1183), .O(gate454inter8));
  nand2 gate878(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate879(.a(s_47), .b(gate454inter3), .O(gate454inter10));
  nor2  gate880(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate881(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate882(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate995(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate996(.a(gate455inter0), .b(s_64), .O(gate455inter1));
  and2  gate997(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate998(.a(s_64), .O(gate455inter3));
  inv1  gate999(.a(s_65), .O(gate455inter4));
  nand2 gate1000(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1001(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1002(.a(G19), .O(gate455inter7));
  inv1  gate1003(.a(G1186), .O(gate455inter8));
  nand2 gate1004(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1005(.a(s_65), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1006(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1007(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1008(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1303(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1304(.a(gate456inter0), .b(s_108), .O(gate456inter1));
  and2  gate1305(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1306(.a(s_108), .O(gate456inter3));
  inv1  gate1307(.a(s_109), .O(gate456inter4));
  nand2 gate1308(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1309(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1310(.a(G1090), .O(gate456inter7));
  inv1  gate1311(.a(G1186), .O(gate456inter8));
  nand2 gate1312(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1313(.a(s_109), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1314(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1315(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1316(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1625(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1626(.a(gate460inter0), .b(s_154), .O(gate460inter1));
  and2  gate1627(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1628(.a(s_154), .O(gate460inter3));
  inv1  gate1629(.a(s_155), .O(gate460inter4));
  nand2 gate1630(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1631(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1632(.a(G1096), .O(gate460inter7));
  inv1  gate1633(.a(G1192), .O(gate460inter8));
  nand2 gate1634(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1635(.a(s_155), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1636(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1637(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1638(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate1639(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1640(.a(gate461inter0), .b(s_156), .O(gate461inter1));
  and2  gate1641(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1642(.a(s_156), .O(gate461inter3));
  inv1  gate1643(.a(s_157), .O(gate461inter4));
  nand2 gate1644(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1645(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1646(.a(G22), .O(gate461inter7));
  inv1  gate1647(.a(G1195), .O(gate461inter8));
  nand2 gate1648(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1649(.a(s_157), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1650(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1651(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1652(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate939(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate940(.a(gate462inter0), .b(s_56), .O(gate462inter1));
  and2  gate941(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate942(.a(s_56), .O(gate462inter3));
  inv1  gate943(.a(s_57), .O(gate462inter4));
  nand2 gate944(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate945(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate946(.a(G1099), .O(gate462inter7));
  inv1  gate947(.a(G1195), .O(gate462inter8));
  nand2 gate948(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate949(.a(s_57), .b(gate462inter3), .O(gate462inter10));
  nor2  gate950(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate951(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate952(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2157(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2158(.a(gate463inter0), .b(s_230), .O(gate463inter1));
  and2  gate2159(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2160(.a(s_230), .O(gate463inter3));
  inv1  gate2161(.a(s_231), .O(gate463inter4));
  nand2 gate2162(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2163(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2164(.a(G23), .O(gate463inter7));
  inv1  gate2165(.a(G1198), .O(gate463inter8));
  nand2 gate2166(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2167(.a(s_231), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2168(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2169(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2170(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1079(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1080(.a(gate465inter0), .b(s_76), .O(gate465inter1));
  and2  gate1081(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1082(.a(s_76), .O(gate465inter3));
  inv1  gate1083(.a(s_77), .O(gate465inter4));
  nand2 gate1084(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1085(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1086(.a(G24), .O(gate465inter7));
  inv1  gate1087(.a(G1201), .O(gate465inter8));
  nand2 gate1088(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1089(.a(s_77), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1090(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1091(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1092(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2955(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2956(.a(gate466inter0), .b(s_344), .O(gate466inter1));
  and2  gate2957(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2958(.a(s_344), .O(gate466inter3));
  inv1  gate2959(.a(s_345), .O(gate466inter4));
  nand2 gate2960(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2961(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2962(.a(G1105), .O(gate466inter7));
  inv1  gate2963(.a(G1201), .O(gate466inter8));
  nand2 gate2964(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2965(.a(s_345), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2966(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2967(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2968(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate645(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate646(.a(gate468inter0), .b(s_14), .O(gate468inter1));
  and2  gate647(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate648(.a(s_14), .O(gate468inter3));
  inv1  gate649(.a(s_15), .O(gate468inter4));
  nand2 gate650(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate651(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate652(.a(G1108), .O(gate468inter7));
  inv1  gate653(.a(G1204), .O(gate468inter8));
  nand2 gate654(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate655(.a(s_15), .b(gate468inter3), .O(gate468inter10));
  nor2  gate656(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate657(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate658(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2269(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2270(.a(gate470inter0), .b(s_246), .O(gate470inter1));
  and2  gate2271(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2272(.a(s_246), .O(gate470inter3));
  inv1  gate2273(.a(s_247), .O(gate470inter4));
  nand2 gate2274(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2275(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2276(.a(G1111), .O(gate470inter7));
  inv1  gate2277(.a(G1207), .O(gate470inter8));
  nand2 gate2278(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2279(.a(s_247), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2280(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2281(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2282(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2213(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2214(.a(gate472inter0), .b(s_238), .O(gate472inter1));
  and2  gate2215(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2216(.a(s_238), .O(gate472inter3));
  inv1  gate2217(.a(s_239), .O(gate472inter4));
  nand2 gate2218(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2219(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2220(.a(G1114), .O(gate472inter7));
  inv1  gate2221(.a(G1210), .O(gate472inter8));
  nand2 gate2222(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2223(.a(s_239), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2224(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2225(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2226(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1709(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1710(.a(gate475inter0), .b(s_166), .O(gate475inter1));
  and2  gate1711(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1712(.a(s_166), .O(gate475inter3));
  inv1  gate1713(.a(s_167), .O(gate475inter4));
  nand2 gate1714(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1715(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1716(.a(G29), .O(gate475inter7));
  inv1  gate1717(.a(G1216), .O(gate475inter8));
  nand2 gate1718(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1719(.a(s_167), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1720(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1721(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1722(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate3025(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate3026(.a(gate476inter0), .b(s_354), .O(gate476inter1));
  and2  gate3027(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate3028(.a(s_354), .O(gate476inter3));
  inv1  gate3029(.a(s_355), .O(gate476inter4));
  nand2 gate3030(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate3031(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate3032(.a(G1120), .O(gate476inter7));
  inv1  gate3033(.a(G1216), .O(gate476inter8));
  nand2 gate3034(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate3035(.a(s_355), .b(gate476inter3), .O(gate476inter10));
  nor2  gate3036(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate3037(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate3038(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate743(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate744(.a(gate477inter0), .b(s_28), .O(gate477inter1));
  and2  gate745(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate746(.a(s_28), .O(gate477inter3));
  inv1  gate747(.a(s_29), .O(gate477inter4));
  nand2 gate748(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate749(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate750(.a(G30), .O(gate477inter7));
  inv1  gate751(.a(G1219), .O(gate477inter8));
  nand2 gate752(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate753(.a(s_29), .b(gate477inter3), .O(gate477inter10));
  nor2  gate754(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate755(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate756(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1191(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1192(.a(gate478inter0), .b(s_92), .O(gate478inter1));
  and2  gate1193(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1194(.a(s_92), .O(gate478inter3));
  inv1  gate1195(.a(s_93), .O(gate478inter4));
  nand2 gate1196(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1197(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1198(.a(G1123), .O(gate478inter7));
  inv1  gate1199(.a(G1219), .O(gate478inter8));
  nand2 gate1200(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1201(.a(s_93), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1202(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1203(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1204(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate617(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate618(.a(gate479inter0), .b(s_10), .O(gate479inter1));
  and2  gate619(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate620(.a(s_10), .O(gate479inter3));
  inv1  gate621(.a(s_11), .O(gate479inter4));
  nand2 gate622(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate623(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate624(.a(G31), .O(gate479inter7));
  inv1  gate625(.a(G1222), .O(gate479inter8));
  nand2 gate626(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate627(.a(s_11), .b(gate479inter3), .O(gate479inter10));
  nor2  gate628(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate629(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate630(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate841(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate842(.a(gate482inter0), .b(s_42), .O(gate482inter1));
  and2  gate843(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate844(.a(s_42), .O(gate482inter3));
  inv1  gate845(.a(s_43), .O(gate482inter4));
  nand2 gate846(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate847(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate848(.a(G1129), .O(gate482inter7));
  inv1  gate849(.a(G1225), .O(gate482inter8));
  nand2 gate850(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate851(.a(s_43), .b(gate482inter3), .O(gate482inter10));
  nor2  gate852(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate853(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate854(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1345(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1346(.a(gate483inter0), .b(s_114), .O(gate483inter1));
  and2  gate1347(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1348(.a(s_114), .O(gate483inter3));
  inv1  gate1349(.a(s_115), .O(gate483inter4));
  nand2 gate1350(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1351(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1352(.a(G1228), .O(gate483inter7));
  inv1  gate1353(.a(G1229), .O(gate483inter8));
  nand2 gate1354(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1355(.a(s_115), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1356(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1357(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1358(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1401(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1402(.a(gate484inter0), .b(s_122), .O(gate484inter1));
  and2  gate1403(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1404(.a(s_122), .O(gate484inter3));
  inv1  gate1405(.a(s_123), .O(gate484inter4));
  nand2 gate1406(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1407(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1408(.a(G1230), .O(gate484inter7));
  inv1  gate1409(.a(G1231), .O(gate484inter8));
  nand2 gate1410(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1411(.a(s_123), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1412(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1413(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1414(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate827(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate828(.a(gate487inter0), .b(s_40), .O(gate487inter1));
  and2  gate829(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate830(.a(s_40), .O(gate487inter3));
  inv1  gate831(.a(s_41), .O(gate487inter4));
  nand2 gate832(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate833(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate834(.a(G1236), .O(gate487inter7));
  inv1  gate835(.a(G1237), .O(gate487inter8));
  nand2 gate836(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate837(.a(s_41), .b(gate487inter3), .O(gate487inter10));
  nor2  gate838(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate839(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate840(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2381(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2382(.a(gate489inter0), .b(s_262), .O(gate489inter1));
  and2  gate2383(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2384(.a(s_262), .O(gate489inter3));
  inv1  gate2385(.a(s_263), .O(gate489inter4));
  nand2 gate2386(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2387(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2388(.a(G1240), .O(gate489inter7));
  inv1  gate2389(.a(G1241), .O(gate489inter8));
  nand2 gate2390(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2391(.a(s_263), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2392(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2393(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2394(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate2451(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2452(.a(gate490inter0), .b(s_272), .O(gate490inter1));
  and2  gate2453(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2454(.a(s_272), .O(gate490inter3));
  inv1  gate2455(.a(s_273), .O(gate490inter4));
  nand2 gate2456(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2457(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2458(.a(G1242), .O(gate490inter7));
  inv1  gate2459(.a(G1243), .O(gate490inter8));
  nand2 gate2460(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2461(.a(s_273), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2462(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2463(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2464(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate2101(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2102(.a(gate491inter0), .b(s_222), .O(gate491inter1));
  and2  gate2103(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2104(.a(s_222), .O(gate491inter3));
  inv1  gate2105(.a(s_223), .O(gate491inter4));
  nand2 gate2106(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2107(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2108(.a(G1244), .O(gate491inter7));
  inv1  gate2109(.a(G1245), .O(gate491inter8));
  nand2 gate2110(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2111(.a(s_223), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2112(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2113(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2114(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2577(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2578(.a(gate493inter0), .b(s_290), .O(gate493inter1));
  and2  gate2579(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2580(.a(s_290), .O(gate493inter3));
  inv1  gate2581(.a(s_291), .O(gate493inter4));
  nand2 gate2582(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2583(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2584(.a(G1248), .O(gate493inter7));
  inv1  gate2585(.a(G1249), .O(gate493inter8));
  nand2 gate2586(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2587(.a(s_291), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2588(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2589(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2590(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate2661(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2662(.a(gate495inter0), .b(s_302), .O(gate495inter1));
  and2  gate2663(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2664(.a(s_302), .O(gate495inter3));
  inv1  gate2665(.a(s_303), .O(gate495inter4));
  nand2 gate2666(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2667(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2668(.a(G1252), .O(gate495inter7));
  inv1  gate2669(.a(G1253), .O(gate495inter8));
  nand2 gate2670(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2671(.a(s_303), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2672(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2673(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2674(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1835(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1836(.a(gate499inter0), .b(s_184), .O(gate499inter1));
  and2  gate1837(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1838(.a(s_184), .O(gate499inter3));
  inv1  gate1839(.a(s_185), .O(gate499inter4));
  nand2 gate1840(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1841(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1842(.a(G1260), .O(gate499inter7));
  inv1  gate1843(.a(G1261), .O(gate499inter8));
  nand2 gate1844(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1845(.a(s_185), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1846(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1847(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1848(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1919(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1920(.a(gate505inter0), .b(s_196), .O(gate505inter1));
  and2  gate1921(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1922(.a(s_196), .O(gate505inter3));
  inv1  gate1923(.a(s_197), .O(gate505inter4));
  nand2 gate1924(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1925(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1926(.a(G1272), .O(gate505inter7));
  inv1  gate1927(.a(G1273), .O(gate505inter8));
  nand2 gate1928(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1929(.a(s_197), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1930(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1931(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1932(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate2409(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2410(.a(gate506inter0), .b(s_266), .O(gate506inter1));
  and2  gate2411(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2412(.a(s_266), .O(gate506inter3));
  inv1  gate2413(.a(s_267), .O(gate506inter4));
  nand2 gate2414(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2415(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2416(.a(G1274), .O(gate506inter7));
  inv1  gate2417(.a(G1275), .O(gate506inter8));
  nand2 gate2418(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2419(.a(s_267), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2420(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2421(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2422(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1737(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1738(.a(gate507inter0), .b(s_170), .O(gate507inter1));
  and2  gate1739(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1740(.a(s_170), .O(gate507inter3));
  inv1  gate1741(.a(s_171), .O(gate507inter4));
  nand2 gate1742(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1743(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1744(.a(G1276), .O(gate507inter7));
  inv1  gate1745(.a(G1277), .O(gate507inter8));
  nand2 gate1746(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1747(.a(s_171), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1748(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1749(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1750(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2745(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2746(.a(gate508inter0), .b(s_314), .O(gate508inter1));
  and2  gate2747(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2748(.a(s_314), .O(gate508inter3));
  inv1  gate2749(.a(s_315), .O(gate508inter4));
  nand2 gate2750(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2751(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2752(.a(G1278), .O(gate508inter7));
  inv1  gate2753(.a(G1279), .O(gate508inter8));
  nand2 gate2754(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2755(.a(s_315), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2756(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2757(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2758(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate561(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate562(.a(gate509inter0), .b(s_2), .O(gate509inter1));
  and2  gate563(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate564(.a(s_2), .O(gate509inter3));
  inv1  gate565(.a(s_3), .O(gate509inter4));
  nand2 gate566(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate567(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate568(.a(G1280), .O(gate509inter7));
  inv1  gate569(.a(G1281), .O(gate509inter8));
  nand2 gate570(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate571(.a(s_3), .b(gate509inter3), .O(gate509inter10));
  nor2  gate572(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate573(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate574(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule